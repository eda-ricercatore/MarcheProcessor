
module RegFileWW ( rd1data, rd2data, wrdata, rd1addr, rd2addr, wraddr, rd1en, 
        rd2en, wren, wrbyteen, clk );
  output [127:0] rd1data;
  output [127:0] rd2data;
  input [0:127] wrdata;
  input [4:0] rd1addr;
  input [4:0] rd2addr;
  input [4:0] wraddr;
  input [15:0] wrbyteen;
  input rd1en, rd2en, wren, clk;
  wire   rd1data1033_127_, rd1data1033_126_, rd1data1033_125_,
         rd1data1033_124_, rd1data1033_123_, rd1data1033_122_,
         rd1data1033_121_, rd1data1033_120_, rd1data1033_119_,
         rd1data1033_118_, rd1data1033_117_, rd1data1033_116_,
         rd1data1033_115_, rd1data1033_114_, rd1data1033_113_,
         rd1data1033_112_, rd1data1033_111_, rd1data1033_110_,
         rd1data1033_109_, rd1data1033_108_, rd1data1033_107_,
         rd1data1033_106_, rd1data1033_105_, rd1data1033_104_,
         rd1data1033_103_, rd1data1033_102_, rd1data1033_101_,
         rd1data1033_100_, rd1data1033_99_, rd1data1033_98_, rd1data1033_97_,
         rd1data1033_96_, rd1data1033_95_, rd1data1033_94_, rd1data1033_93_,
         rd1data1033_92_, rd1data1033_91_, rd1data1033_90_, rd1data1033_89_,
         rd1data1033_88_, rd1data1033_87_, rd1data1033_86_, rd1data1033_85_,
         rd1data1033_84_, rd1data1033_83_, rd1data1033_82_, rd1data1033_81_,
         rd1data1033_80_, rd1data1033_79_, rd1data1033_78_, rd1data1033_77_,
         rd1data1033_76_, rd1data1033_75_, rd1data1033_74_, rd1data1033_73_,
         rd1data1033_72_, rd1data1033_71_, rd1data1033_70_, rd1data1033_69_,
         rd1data1033_68_, rd1data1033_67_, rd1data1033_66_, rd1data1033_65_,
         rd1data1033_64_, rd1data1033_63_, rd1data1033_62_, rd1data1033_61_,
         rd1data1033_60_, rd1data1033_59_, rd1data1033_58_, rd1data1033_57_,
         rd1data1033_56_, rd1data1033_55_, rd1data1033_54_, rd1data1033_53_,
         rd1data1033_52_, rd1data1033_51_, rd1data1033_50_, rd1data1033_49_,
         rd1data1033_48_, rd1data1033_47_, rd1data1033_46_, rd1data1033_45_,
         rd1data1033_44_, rd1data1033_43_, rd1data1033_42_, rd1data1033_41_,
         rd1data1033_40_, rd1data1033_39_, rd1data1033_38_, rd1data1033_37_,
         rd1data1033_36_, rd1data1033_35_, rd1data1033_34_, rd1data1033_33_,
         rd1data1033_32_, rd1data1033_31_, rd1data1033_30_, rd1data1033_29_,
         rd1data1033_28_, rd1data1033_27_, rd1data1033_26_, rd1data1033_25_,
         rd1data1033_24_, rd1data1033_23_, rd1data1033_22_, rd1data1033_21_,
         rd1data1033_20_, rd1data1033_19_, rd1data1033_18_, rd1data1033_17_,
         rd1data1033_16_, rd1data1033_15_, rd1data1033_14_, rd1data1033_13_,
         rd1data1033_12_, rd1data1033_11_, rd1data1033_10_, rd1data1033_9_,
         rd1data1033_8_, rd1data1033_7_, rd1data1033_6_, rd1data1033_5_,
         rd1data1033_4_, rd1data1033_3_, rd1data1033_2_, rd1data1033_1_,
         rd1data1033_0_, rd2data1040_127_, rd2data1040_126_, rd2data1040_125_,
         rd2data1040_124_, rd2data1040_123_, rd2data1040_122_,
         rd2data1040_121_, rd2data1040_120_, rd2data1040_119_,
         rd2data1040_118_, rd2data1040_117_, rd2data1040_116_,
         rd2data1040_115_, rd2data1040_114_, rd2data1040_113_,
         rd2data1040_112_, rd2data1040_111_, rd2data1040_110_,
         rd2data1040_109_, rd2data1040_108_, rd2data1040_107_,
         rd2data1040_106_, rd2data1040_105_, rd2data1040_104_,
         rd2data1040_103_, rd2data1040_102_, rd2data1040_101_,
         rd2data1040_100_, rd2data1040_99_, rd2data1040_98_, rd2data1040_97_,
         rd2data1040_96_, rd2data1040_95_, rd2data1040_94_, rd2data1040_93_,
         rd2data1040_92_, rd2data1040_91_, rd2data1040_90_, rd2data1040_89_,
         rd2data1040_88_, rd2data1040_87_, rd2data1040_86_, rd2data1040_85_,
         rd2data1040_84_, rd2data1040_83_, rd2data1040_82_, rd2data1040_81_,
         rd2data1040_80_, rd2data1040_79_, rd2data1040_78_, rd2data1040_77_,
         rd2data1040_76_, rd2data1040_75_, rd2data1040_74_, rd2data1040_73_,
         rd2data1040_72_, rd2data1040_71_, rd2data1040_70_, rd2data1040_69_,
         rd2data1040_68_, rd2data1040_67_, rd2data1040_66_, rd2data1040_65_,
         rd2data1040_64_, rd2data1040_63_, rd2data1040_62_, rd2data1040_61_,
         rd2data1040_60_, rd2data1040_59_, rd2data1040_58_, rd2data1040_57_,
         rd2data1040_56_, rd2data1040_55_, rd2data1040_54_, rd2data1040_53_,
         rd2data1040_52_, rd2data1040_51_, rd2data1040_50_, rd2data1040_49_,
         rd2data1040_48_, rd2data1040_47_, rd2data1040_46_, rd2data1040_45_,
         rd2data1040_44_, rd2data1040_43_, rd2data1040_42_, rd2data1040_41_,
         rd2data1040_40_, rd2data1040_39_, rd2data1040_38_, rd2data1040_37_,
         rd2data1040_36_, rd2data1040_35_, rd2data1040_34_, rd2data1040_33_,
         rd2data1040_32_, rd2data1040_31_, rd2data1040_30_, rd2data1040_29_,
         rd2data1040_28_, rd2data1040_27_, rd2data1040_26_, rd2data1040_25_,
         rd2data1040_24_, rd2data1040_23_, rd2data1040_22_, rd2data1040_21_,
         rd2data1040_20_, rd2data1040_19_, rd2data1040_18_, rd2data1040_17_,
         rd2data1040_16_, rd2data1040_15_, rd2data1040_14_, rd2data1040_13_,
         rd2data1040_12_, rd2data1040_11_, rd2data1040_10_, rd2data1040_9_,
         rd2data1040_8_, rd2data1040_7_, rd2data1040_6_, rd2data1040_5_,
         rd2data1040_4_, rd2data1040_3_, rd2data1040_2_, rd2data1040_1_,
         rd2data1040_0_, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
         n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
         n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
         n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750,
         n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
         n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
         n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782,
         n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
         n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798,
         n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
         n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
         n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822,
         n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
         n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
         n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
         n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
         n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
         n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
         n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
         n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942,
         n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
         n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958,
         n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966,
         n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
         n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
         n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990,
         n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
         n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
         n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014,
         n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
         n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
         n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
         n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
         n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
         n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
         n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
         n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
         n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086,
         n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
         n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302,
         n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
         n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
         n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
         n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334,
         n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
         n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350,
         n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358,
         n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366,
         n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374,
         n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
         n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
         n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
         n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406,
         n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
         n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422,
         n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430,
         n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438,
         n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446,
         n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
         n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
         n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470,
         n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478,
         n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486,
         n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494,
         n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502,
         n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510,
         n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518,
         n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526,
         n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
         n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542,
         n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550,
         n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558,
         n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566,
         n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574,
         n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582,
         n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590,
         n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598,
         n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606,
         n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614,
         n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
         n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630,
         n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638,
         n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
         n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654,
         n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662,
         n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
         n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
         n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686,
         n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694,
         n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
         n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710,
         n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718,
         n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726,
         n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734,
         n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742,
         n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750,
         n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758,
         n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766,
         n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774,
         n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782,
         n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790,
         n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798,
         n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806,
         n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814,
         n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822,
         n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830,
         n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838,
         n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846,
         n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854,
         n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862,
         n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870,
         n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878,
         n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886,
         n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894,
         n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902,
         n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910,
         n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918,
         n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926,
         n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934,
         n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942,
         n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950,
         n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958,
         n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966,
         n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974,
         n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982,
         n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990,
         n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998,
         n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006,
         n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014,
         n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022,
         n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030,
         n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038,
         n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046,
         n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054,
         n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
         n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070,
         n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078,
         n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086,
         n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094,
         n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102,
         n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110,
         n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118,
         n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
         n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134,
         n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142,
         n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150,
         n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158,
         n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166,
         n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174,
         n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182,
         n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
         n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
         n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
         n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214,
         n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222,
         n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230,
         n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238,
         n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
         n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254,
         n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262,
         n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270,
         n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278,
         n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286,
         n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294,
         n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
         n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310,
         n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318,
         n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326,
         n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334,
         n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342,
         n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350,
         n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358,
         n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366,
         n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
         n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382,
         n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390,
         n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398,
         n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406,
         n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414,
         n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422,
         n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430,
         n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438,
         n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446,
         n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454,
         n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462,
         n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470,
         n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478,
         n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486,
         n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
         n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502,
         n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510,
         n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
         n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526,
         n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534,
         n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542,
         n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550,
         n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558,
         n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
         n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
         n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582,
         n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
         n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598,
         n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
         n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
         n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
         n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630,
         n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
         n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646,
         n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654,
         n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
         n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670,
         n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678,
         n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686,
         n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
         n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
         n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
         n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
         n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
         n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
         n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742,
         n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750,
         n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
         n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
         n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774,
         n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782,
         n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790,
         n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
         n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
         n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814,
         n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822,
         n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
         n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838,
         n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846,
         n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854,
         n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862,
         n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870,
         n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878,
         n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886,
         n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894,
         n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
         n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910,
         n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918,
         n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926,
         n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934,
         n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942,
         n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950,
         n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958,
         n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966,
         n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
         n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982,
         n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990,
         n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
         n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006,
         n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014,
         n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022,
         n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030,
         n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038,
         n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
         n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054,
         n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062,
         n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
         n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078,
         n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086,
         n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094,
         n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102,
         n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110,
         n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
         n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126,
         n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134,
         n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
         n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150,
         n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158,
         n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166,
         n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174,
         n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
         n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
         n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198,
         n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206,
         n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
         n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222,
         n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230,
         n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238,
         n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246,
         n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
         n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262,
         n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270,
         n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
         n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
         n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294,
         n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302,
         n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310,
         n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318,
         n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
         n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
         n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
         n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350,
         n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
         n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366,
         n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374,
         n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382,
         n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390,
         n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
         n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
         n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414,
         n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422,
         n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430,
         n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438,
         n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446,
         n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454,
         n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462,
         n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
         n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478,
         n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486,
         n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
         n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
         n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510,
         n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518,
         n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
         n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534,
         n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
         n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550,
         n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558,
         n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566,
         n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
         n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582,
         n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590,
         n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598,
         n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606,
         n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
         n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622,
         n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630,
         n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638,
         n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
         n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654,
         n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662,
         n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670,
         n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678,
         n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686,
         n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694,
         n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702,
         n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710,
         n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
         n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726,
         n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734,
         n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
         n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
         n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758,
         n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766,
         n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774,
         n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782,
         n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
         n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798,
         n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806,
         n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
         n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
         n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
         n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
         n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846,
         n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
         n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
         n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870,
         n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878,
         n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
         n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
         n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902,
         n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
         n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918,
         n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
         n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934,
         n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942,
         n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950,
         n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958,
         n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966,
         n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974,
         n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982,
         n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990,
         n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998,
         n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006,
         n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014,
         n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022,
         n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
         n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038,
         n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046,
         n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054,
         n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062,
         n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070,
         n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
         n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086,
         n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094,
         n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102,
         n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
         n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118,
         n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126,
         n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134,
         n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142,
         n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150,
         n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158,
         n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166,
         n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
         n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182,
         n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190,
         n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
         n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206,
         n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214,
         n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222,
         n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230,
         n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238,
         n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
         n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254,
         n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262,
         n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270,
         n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278,
         n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286,
         n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294,
         n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302,
         n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310,
         n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
         n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326,
         n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334,
         n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342,
         n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350,
         n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358,
         n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366,
         n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374,
         n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382,
         n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
         n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398,
         n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
         n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414,
         n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422,
         n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430,
         n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
         n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446,
         n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454,
         n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
         n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470,
         n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
         n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486,
         n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494,
         n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502,
         n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
         n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
         n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526,
         n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
         n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542,
         n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
         n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558,
         n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566,
         n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574,
         n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
         n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590,
         n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598,
         n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606,
         n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614,
         n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
         n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630,
         n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638,
         n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646,
         n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654,
         n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
         n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670,
         n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
         n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686,
         n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
         n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702,
         n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710,
         n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
         n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
         n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734,
         n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742,
         n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
         n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758,
         n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
         n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774,
         n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782,
         n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
         n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798,
         n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806,
         n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814,
         n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
         n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830,
         n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
         n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846,
         n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854,
         n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862,
         n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
         n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878,
         n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
         n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
         n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902,
         n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
         n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918,
         n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
         n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934,
         n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
         n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950,
         n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
         n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
         n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974,
         n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
         n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990,
         n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998,
         n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006,
         n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
         n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022,
         n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030,
         n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038,
         n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046,
         n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
         n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
         n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070,
         n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078,
         n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086,
         n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094,
         n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102,
         n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110,
         n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118,
         n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
         n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
         n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142,
         n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
         n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
         n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
         n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174,
         n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
         n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190,
         n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
         n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
         n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214,
         n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222,
         n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
         n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238,
         n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246,
         n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
         n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
         n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
         n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278,
         n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286,
         n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294,
         n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
         n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310,
         n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318,
         n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326,
         n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334,
         n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
         n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350,
         n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358,
         n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366,
         n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374,
         n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382,
         n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390,
         n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
         n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406,
         n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
         n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422,
         n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430,
         n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438,
         n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446,
         n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454,
         n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462,
         n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470,
         n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478,
         n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486,
         n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494,
         n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502,
         n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510,
         n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518,
         n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526,
         n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534,
         n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542,
         n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550,
         n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558,
         n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566,
         n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574,
         n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582,
         n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590,
         n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598,
         n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606,
         n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614,
         n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622,
         n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630,
         n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638,
         n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646,
         n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654,
         n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662,
         n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670,
         n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678,
         n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686,
         n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694,
         n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702,
         n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
         n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718,
         n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726,
         n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734,
         n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742,
         n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750,
         n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758,
         n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766,
         n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
         n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782,
         n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790,
         n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798,
         n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
         n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814,
         n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822,
         n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830,
         n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838,
         n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
         n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854,
         n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862,
         n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870,
         n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
         n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886,
         n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894,
         n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902,
         n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910,
         n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
         n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926,
         n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934,
         n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
         n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950,
         n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958,
         n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966,
         n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
         n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982,
         n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990,
         n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998,
         n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006,
         n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014,
         n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022,
         n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030,
         n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038,
         n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046,
         n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054,
         n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062,
         n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070,
         n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078,
         n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
         n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094,
         n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102,
         n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110,
         n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
         n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126,
         n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
         n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142,
         n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150,
         n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158,
         n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166,
         n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174,
         n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182,
         n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190,
         n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198,
         n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206,
         n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214,
         n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222,
         n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
         n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238,
         n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246,
         n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254,
         n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262,
         n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270,
         n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
         n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286,
         n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294,
         n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302,
         n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310,
         n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318,
         n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326,
         n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334,
         n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342,
         n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350,
         n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358,
         n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366,
         n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
         n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382,
         n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390,
         n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398,
         n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406,
         n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414,
         n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422,
         n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430,
         n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438,
         n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
         n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454,
         n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462,
         n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470,
         n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
         n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486,
         n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494,
         n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502,
         n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510,
         n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518,
         n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526,
         n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534,
         n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542,
         n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550,
         n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558,
         n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566,
         n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574,
         n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582,
         n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590,
         n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
         n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606,
         n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614,
         n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622,
         n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630,
         n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638,
         n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646,
         n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654,
         n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662,
         n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670,
         n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678,
         n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686,
         n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694,
         n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702,
         n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710,
         n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718,
         n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726,
         n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734,
         n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742,
         n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750,
         n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758,
         n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
         n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774,
         n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
         n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790,
         n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798,
         n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
         n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814,
         n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822,
         n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830,
         n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838,
         n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846,
         n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
         n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862,
         n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870,
         n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
         n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886,
         n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894,
         n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902,
         n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
         n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918,
         n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
         n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934,
         n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942,
         n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950,
         n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958,
         n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966,
         n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974,
         n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982,
         n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990,
         n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998,
         n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006,
         n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014,
         n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022,
         n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030,
         n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038,
         n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046,
         n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054,
         n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062,
         n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070,
         n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078,
         n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086,
         n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094,
         n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
         n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110,
         n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118,
         n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126,
         n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134,
         n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142,
         n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150,
         n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158,
         n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166,
         n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174,
         n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182,
         n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190,
         n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198,
         n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206,
         n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214,
         n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222,
         n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230,
         n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238,
         n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246,
         n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254,
         n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262,
         n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270,
         n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278,
         n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286,
         n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
         n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
         n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310,
         n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318,
         n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326,
         n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334,
         n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
         n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350,
         n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358,
         n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366,
         n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374,
         n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382,
         n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390,
         n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398,
         n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406,
         n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
         n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422,
         n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430,
         n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
         n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446,
         n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
         n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
         n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470,
         n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478,
         n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486,
         n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494,
         n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
         n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
         n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518,
         n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526,
         n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534,
         n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542,
         n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550,
         n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558,
         n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566,
         n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
         n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582,
         n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590,
         n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598,
         n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606,
         n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614,
         n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622,
         n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630,
         n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638,
         n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
         n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654,
         n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662,
         n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670,
         n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678,
         n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686,
         n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694,
         n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
         n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710,
         n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
         n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726,
         n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734,
         n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742,
         n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750,
         n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758,
         n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766,
         n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
         n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782,
         n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
         n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798,
         n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806,
         n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814,
         n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822,
         n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830,
         n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838,
         n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846,
         n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854,
         n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
         n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870,
         n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878,
         n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886,
         n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894,
         n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902,
         n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910,
         n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918,
         n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
         n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934,
         n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942,
         n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950,
         n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958,
         n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
         n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974,
         n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982,
         n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990,
         n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
         n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006,
         n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014,
         n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022,
         n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030,
         n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038,
         n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046,
         n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054,
         n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
         n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
         n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
         n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086,
         n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094,
         n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102,
         n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
         n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118,
         n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126,
         n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
         n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142,
         n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150,
         n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158,
         n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166,
         n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
         n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182,
         n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190,
         n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198,
         n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
         n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
         n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
         n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
         n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238,
         n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
         n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
         n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262,
         n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270,
         n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
         n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
         n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
         n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302,
         n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310,
         n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318,
         n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326,
         n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334,
         n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342,
         n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
         n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358,
         n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
         n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374,
         n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382,
         n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390,
         n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398,
         n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406,
         n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414,
         n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
         n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430,
         n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
         n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446,
         n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454,
         n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
         n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
         n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478,
         n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
         n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
         n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502,
         n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510,
         n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518,
         n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526,
         n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534,
         n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542,
         n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550,
         n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558,
         n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
         n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574,
         n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582,
         n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590,
         n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598,
         n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606,
         n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614,
         n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622,
         n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630,
         n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
         n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646,
         n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654,
         n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
         n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670,
         n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678,
         n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686,
         n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694,
         n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702,
         n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
         n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
         n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
         n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742,
         n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
         n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758,
         n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766,
         n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774,
         n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
         n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790,
         n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
         n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806,
         n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814,
         n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822,
         n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
         n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
         n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862,
         n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
         n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
         n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886,
         n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894,
         n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
         n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
         n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918,
         n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
         n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934,
         n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
         n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950,
         n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958,
         n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
         n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
         n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982,
         n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
         n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
         n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006,
         n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
         n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022,
         n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030,
         n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
         n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046,
         n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
         n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062,
         n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
         n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
         n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
         n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
         n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102,
         n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
         n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
         n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126,
         n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
         n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
         n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150,
         n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
         n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166,
         n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174,
         n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
         n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
         n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198,
         n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
         n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
         n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222,
         n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
         n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238,
         n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246,
         n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
         n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
         n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270,
         n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278,
         n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
         n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294,
         n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
         n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310,
         n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318,
         n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326,
         n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
         n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342,
         n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350,
         n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
         n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366,
         n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
         n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
         n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390,
         n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
         n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
         n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414,
         n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
         n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
         n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438,
         n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
         n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
         n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462,
         n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470,
         n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478,
         n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
         n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
         n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510,
         n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
         n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526,
         n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534,
         n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
         n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
         n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
         n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566,
         n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
         n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582,
         n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
         n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598,
         n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606,
         n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
         n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
         n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630,
         n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638,
         n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
         n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654,
         n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662,
         n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670,
         n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678,
         n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686,
         n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694,
         n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702,
         n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710,
         n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
         n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726,
         n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
         n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742,
         n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750,
         n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758,
         n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766,
         n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774,
         n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782,
         n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
         n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798,
         n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
         n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814,
         n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822,
         n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
         n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
         n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846,
         n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854,
         n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
         n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870,
         n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878,
         n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886,
         n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894,
         n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902,
         n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910,
         n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918,
         n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926,
         n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
         n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942,
         n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950,
         n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958,
         n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966,
         n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974,
         n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982,
         n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990,
         n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998,
         n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006,
         n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014,
         n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022,
         n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030,
         n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038,
         n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046,
         n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
         n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062,
         n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070,
         n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
         n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086,
         n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
         n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110,
         n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118,
         n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
         n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134,
         n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142,
         n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150,
         n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158,
         n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166,
         n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174,
         n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182,
         n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190,
         n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
         n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206,
         n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214,
         n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
         n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230,
         n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
         n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246,
         n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254,
         n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262,
         n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270,
         n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278,
         n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286,
         n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294,
         n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302,
         n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
         n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318,
         n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326,
         n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
         n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342,
         n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350,
         n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358,
         n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366,
         n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374,
         n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382,
         n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390,
         n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398,
         n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406,
         n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414,
         n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422,
         n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430,
         n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
         n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446,
         n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454,
         n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462,
         n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470,
         n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
         n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
         n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494,
         n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502,
         n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
         n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518,
         n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
         n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
         n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542,
         n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
         n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
         n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566,
         n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574,
         n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582,
         n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590,
         n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
         n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606,
         n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614,
         n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622,
         n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630,
         n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638,
         n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646,
         n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
         n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662,
         n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
         n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678,
         n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686,
         n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694,
         n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702,
         n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710,
         n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718,
         n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726,
         n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734,
         n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
         n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750,
         n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758,
         n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766,
         n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
         n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782,
         n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790,
         n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798,
         n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806,
         n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814,
         n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822,
         n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830,
         n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838,
         n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846,
         n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854,
         n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862,
         n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870,
         n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878,
         n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886,
         n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894,
         n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902,
         n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910,
         n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918,
         n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926,
         n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934,
         n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942,
         n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950,
         n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
         n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966,
         n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
         n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
         n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990,
         n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998,
         n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006,
         n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
         n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
         n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
         n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
         n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046,
         n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054,
         n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062,
         n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070,
         n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078,
         n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
         n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094,
         n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
         n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110,
         n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118,
         n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126,
         n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134,
         n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142,
         n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150,
         n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
         n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166,
         n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
         n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182,
         n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190,
         n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198,
         n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206,
         n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214,
         n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222,
         n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
         n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238,
         n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
         n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254,
         n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262,
         n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270,
         n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278,
         n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286,
         n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294,
         n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
         n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310,
         n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318,
         n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
         n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334,
         n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342,
         n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350,
         n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358,
         n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366,
         n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
         n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382,
         n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
         n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398,
         n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406,
         n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414,
         n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422,
         n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430,
         n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
         n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446,
         n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454,
         n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462,
         n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470,
         n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478,
         n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486,
         n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494,
         n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502,
         n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
         n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
         n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526,
         n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534,
         n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542,
         n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550,
         n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558,
         n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566,
         n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574,
         n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
         n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590,
         n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598,
         n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606,
         n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614,
         n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622,
         n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630,
         n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638,
         n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646,
         n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654,
         n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662,
         n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670,
         n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
         n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
         n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694,
         n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
         n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
         n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718,
         n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
         n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
         n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742,
         n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
         n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
         n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766,
         n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
         n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
         n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
         n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
         n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
         n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
         n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
         n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
         n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
         n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
         n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
         n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
         n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030,
         n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
         n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
         n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054,
         n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
         n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
         n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
         n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
         n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102,
         n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
         n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
         n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
         n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
         n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
         n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
         n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158,
         n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
         n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174,
         n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
         n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
         n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198,
         n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
         n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
         n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222,
         n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230,
         n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
         n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
         n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
         n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
         n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270,
         n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
         n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
         n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294,
         n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
         n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
         n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
         n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342,
         n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
         n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
         n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366,
         n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
         n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
         n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390,
         n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
         n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
         n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
         n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
         n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
         n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446,
         n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462,
         n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
         n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
         n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486,
         n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
         n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
         n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
         n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
         n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
         n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534,
         n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
         n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
         n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
         n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
         n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
         n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
         n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590,
         n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
         n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182,
         n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
         n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
         n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206,
         n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
         n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
         n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230,
         n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238,
         n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
         n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254,
         n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
         n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
         n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278,
         n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
         n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
         n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302,
         n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310,
         n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
         n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326,
         n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
         n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
         n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350,
         n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
         n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366,
         n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374,
         n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382,
         n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
         n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398,
         n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
         n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
         n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422,
         n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
         n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
         n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446,
         n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454,
         n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
         n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470,
         n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
         n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
         n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494,
         n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
         n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
         n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518,
         n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
         n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
         n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542,
         n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
         n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558,
         n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566,
         n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
         n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582,
         n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590,
         n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
         n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
         n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614,
         n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
         n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
         n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638,
         n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646,
         n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654,
         n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662,
         n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670,
         n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
         n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686,
         n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
         n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702,
         n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710,
         n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718,
         n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726,
         n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734,
         n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742,
         n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
         n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758,
         n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
         n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774,
         n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782,
         n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790,
         n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798,
         n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806,
         n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814,
         n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
         n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830,
         n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
         n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846,
         n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854,
         n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862,
         n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
         n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878,
         n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886,
         n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
         n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902,
         n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
         n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918,
         n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926,
         n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
         n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
         n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950,
         n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958,
         n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
         n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974,
         n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
         n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990,
         n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
         n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
         n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014,
         n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022,
         n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030,
         n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
         n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046,
         n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
         n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
         n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
         n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
         n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
         n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
         n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102,
         n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
         n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
         n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
         n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134,
         n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142,
         n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
         n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158,
         n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166,
         n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
         n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
         n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190,
         n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
         n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206,
         n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214,
         n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
         n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230,
         n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238,
         n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246,
         n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
         n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262,
         n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
         n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278,
         n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286,
         n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294,
         n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
         n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310,
         n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318,
         n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
         n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334,
         n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
         n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350,
         n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358,
         n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
         n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374,
         n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382,
         n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390,
         n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
         n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406,
         n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
         n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422,
         n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430,
         n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
         n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
         n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454,
         n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462,
         n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
         n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478,
         n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
         n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
         n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502,
         n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
         n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518,
         n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526,
         n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534,
         n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
         n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550,
         n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
         n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
         n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574,
         n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
         n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590,
         n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598,
         n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606,
         n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
         n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622,
         n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
         n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638,
         n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646,
         n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
         n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662,
         n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670,
         n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678,
         n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
         n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694,
         n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
         n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
         n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718,
         n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726,
         n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734,
         n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742,
         n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
         n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
         n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766,
         n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
         n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
         n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790,
         n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798,
         n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806,
         n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814,
         n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
         n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838,
         n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
         n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
         n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862,
         n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870,
         n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878,
         n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886,
         n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
         n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
         n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910,
         n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
         n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926,
         n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934,
         n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942,
         n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
         n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958,
         n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
         n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
         n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982,
         n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
         n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022,
         n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
         n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038,
         n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
         n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054,
         n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
         n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
         n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
         n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
         n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
         n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102,
         n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110,
         n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
         n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126,
         n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
         n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142,
         n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150,
         n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158,
         n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166,
         n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174,
         n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182,
         n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
         n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198,
         n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
         n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214,
         n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222,
         n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230,
         n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238,
         n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246,
         n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254,
         n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
         n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270,
         n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
         n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286,
         n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294,
         n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302,
         n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
         n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318,
         n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326,
         n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
         n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342,
         n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
         n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358,
         n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366,
         n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374,
         n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
         n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390,
         n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398,
         n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
         n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
         n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
         n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
         n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438,
         n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446,
         n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
         n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486,
         n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
         n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502,
         n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510,
         n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
         n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
         n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534,
         n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542,
         n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
         n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558,
         n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
         n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574,
         n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582,
         n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590,
         n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
         n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606,
         n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614,
         n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
         n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
         n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
         n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646,
         n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654,
         n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662,
         n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
         n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678,
         n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686,
         n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
         n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
         n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
         n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718,
         n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726,
         n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
         n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742,
         n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750,
         n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758,
         n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
         n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
         n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
         n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790,
         n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798,
         n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
         n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
         n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822,
         n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830,
         n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
         n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846,
         n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
         n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
         n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
         n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
         n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886,
         n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894,
         n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902,
         n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
         n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918,
         n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
         n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
         n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942,
         n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
         n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958,
         n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966,
         n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974,
         n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
         n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990,
         n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
         n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006,
         n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014,
         n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
         n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030,
         n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
         n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046,
         n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
         n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062,
         n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
         n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
         n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086,
         n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
         n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102,
         n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110,
         n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118,
         n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
         n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134,
         n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
         n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
         n37151, n37152, n37153, n37154, n37155, n37156;
  wire   [4095:0] reg_file;

  DFFPOSX1 reg_file_reg_0__0_ ( .D(n25128), .CLK(clk), .Q(reg_file[0]) );
  DFFPOSX1 reg_file_reg_0__1_ ( .D(n25127), .CLK(clk), .Q(reg_file[1]) );
  DFFPOSX1 reg_file_reg_0__2_ ( .D(n25126), .CLK(clk), .Q(reg_file[2]) );
  DFFPOSX1 reg_file_reg_0__3_ ( .D(n25125), .CLK(clk), .Q(reg_file[3]) );
  DFFPOSX1 reg_file_reg_0__4_ ( .D(n25124), .CLK(clk), .Q(reg_file[4]) );
  DFFPOSX1 reg_file_reg_0__5_ ( .D(n25123), .CLK(clk), .Q(reg_file[5]) );
  DFFPOSX1 reg_file_reg_0__6_ ( .D(n25122), .CLK(clk), .Q(reg_file[6]) );
  DFFPOSX1 reg_file_reg_0__7_ ( .D(n25121), .CLK(clk), .Q(reg_file[7]) );
  DFFPOSX1 reg_file_reg_0__8_ ( .D(n25120), .CLK(clk), .Q(reg_file[8]) );
  DFFPOSX1 reg_file_reg_0__9_ ( .D(n25119), .CLK(clk), .Q(reg_file[9]) );
  DFFPOSX1 reg_file_reg_0__10_ ( .D(n25118), .CLK(clk), .Q(reg_file[10]) );
  DFFPOSX1 reg_file_reg_0__11_ ( .D(n25117), .CLK(clk), .Q(reg_file[11]) );
  DFFPOSX1 reg_file_reg_0__12_ ( .D(n25116), .CLK(clk), .Q(reg_file[12]) );
  DFFPOSX1 reg_file_reg_0__13_ ( .D(n25115), .CLK(clk), .Q(reg_file[13]) );
  DFFPOSX1 reg_file_reg_0__14_ ( .D(n25114), .CLK(clk), .Q(reg_file[14]) );
  DFFPOSX1 reg_file_reg_0__15_ ( .D(n25113), .CLK(clk), .Q(reg_file[15]) );
  DFFPOSX1 reg_file_reg_0__16_ ( .D(n25112), .CLK(clk), .Q(reg_file[16]) );
  DFFPOSX1 reg_file_reg_0__17_ ( .D(n25111), .CLK(clk), .Q(reg_file[17]) );
  DFFPOSX1 reg_file_reg_0__18_ ( .D(n25110), .CLK(clk), .Q(reg_file[18]) );
  DFFPOSX1 reg_file_reg_0__19_ ( .D(n25109), .CLK(clk), .Q(reg_file[19]) );
  DFFPOSX1 reg_file_reg_0__20_ ( .D(n25108), .CLK(clk), .Q(reg_file[20]) );
  DFFPOSX1 reg_file_reg_0__21_ ( .D(n25107), .CLK(clk), .Q(reg_file[21]) );
  DFFPOSX1 reg_file_reg_0__22_ ( .D(n25106), .CLK(clk), .Q(reg_file[22]) );
  DFFPOSX1 reg_file_reg_0__23_ ( .D(n25105), .CLK(clk), .Q(reg_file[23]) );
  DFFPOSX1 reg_file_reg_0__24_ ( .D(n25104), .CLK(clk), .Q(reg_file[24]) );
  DFFPOSX1 reg_file_reg_0__25_ ( .D(n25103), .CLK(clk), .Q(reg_file[25]) );
  DFFPOSX1 reg_file_reg_0__26_ ( .D(n25102), .CLK(clk), .Q(reg_file[26]) );
  DFFPOSX1 reg_file_reg_0__27_ ( .D(n25101), .CLK(clk), .Q(reg_file[27]) );
  DFFPOSX1 reg_file_reg_0__28_ ( .D(n25100), .CLK(clk), .Q(reg_file[28]) );
  DFFPOSX1 reg_file_reg_0__29_ ( .D(n25099), .CLK(clk), .Q(reg_file[29]) );
  DFFPOSX1 reg_file_reg_0__30_ ( .D(n25098), .CLK(clk), .Q(reg_file[30]) );
  DFFPOSX1 reg_file_reg_0__31_ ( .D(n25097), .CLK(clk), .Q(reg_file[31]) );
  DFFPOSX1 reg_file_reg_0__32_ ( .D(n25096), .CLK(clk), .Q(reg_file[32]) );
  DFFPOSX1 reg_file_reg_0__33_ ( .D(n25095), .CLK(clk), .Q(reg_file[33]) );
  DFFPOSX1 reg_file_reg_0__34_ ( .D(n25094), .CLK(clk), .Q(reg_file[34]) );
  DFFPOSX1 reg_file_reg_0__35_ ( .D(n25093), .CLK(clk), .Q(reg_file[35]) );
  DFFPOSX1 reg_file_reg_0__36_ ( .D(n25092), .CLK(clk), .Q(reg_file[36]) );
  DFFPOSX1 reg_file_reg_0__37_ ( .D(n25091), .CLK(clk), .Q(reg_file[37]) );
  DFFPOSX1 reg_file_reg_0__38_ ( .D(n25090), .CLK(clk), .Q(reg_file[38]) );
  DFFPOSX1 reg_file_reg_0__39_ ( .D(n25089), .CLK(clk), .Q(reg_file[39]) );
  DFFPOSX1 reg_file_reg_0__40_ ( .D(n25088), .CLK(clk), .Q(reg_file[40]) );
  DFFPOSX1 reg_file_reg_0__41_ ( .D(n25087), .CLK(clk), .Q(reg_file[41]) );
  DFFPOSX1 reg_file_reg_0__42_ ( .D(n25086), .CLK(clk), .Q(reg_file[42]) );
  DFFPOSX1 reg_file_reg_0__43_ ( .D(n25085), .CLK(clk), .Q(reg_file[43]) );
  DFFPOSX1 reg_file_reg_0__44_ ( .D(n25084), .CLK(clk), .Q(reg_file[44]) );
  DFFPOSX1 reg_file_reg_0__45_ ( .D(n25083), .CLK(clk), .Q(reg_file[45]) );
  DFFPOSX1 reg_file_reg_0__46_ ( .D(n25082), .CLK(clk), .Q(reg_file[46]) );
  DFFPOSX1 reg_file_reg_0__47_ ( .D(n25081), .CLK(clk), .Q(reg_file[47]) );
  DFFPOSX1 reg_file_reg_0__48_ ( .D(n25080), .CLK(clk), .Q(reg_file[48]) );
  DFFPOSX1 reg_file_reg_0__49_ ( .D(n25079), .CLK(clk), .Q(reg_file[49]) );
  DFFPOSX1 reg_file_reg_0__50_ ( .D(n25078), .CLK(clk), .Q(reg_file[50]) );
  DFFPOSX1 reg_file_reg_0__51_ ( .D(n25077), .CLK(clk), .Q(reg_file[51]) );
  DFFPOSX1 reg_file_reg_0__52_ ( .D(n25076), .CLK(clk), .Q(reg_file[52]) );
  DFFPOSX1 reg_file_reg_0__53_ ( .D(n25075), .CLK(clk), .Q(reg_file[53]) );
  DFFPOSX1 reg_file_reg_0__54_ ( .D(n25074), .CLK(clk), .Q(reg_file[54]) );
  DFFPOSX1 reg_file_reg_0__55_ ( .D(n25073), .CLK(clk), .Q(reg_file[55]) );
  DFFPOSX1 reg_file_reg_0__56_ ( .D(n25072), .CLK(clk), .Q(reg_file[56]) );
  DFFPOSX1 reg_file_reg_0__57_ ( .D(n25071), .CLK(clk), .Q(reg_file[57]) );
  DFFPOSX1 reg_file_reg_0__58_ ( .D(n25070), .CLK(clk), .Q(reg_file[58]) );
  DFFPOSX1 reg_file_reg_0__59_ ( .D(n25069), .CLK(clk), .Q(reg_file[59]) );
  DFFPOSX1 reg_file_reg_0__60_ ( .D(n25068), .CLK(clk), .Q(reg_file[60]) );
  DFFPOSX1 reg_file_reg_0__61_ ( .D(n25067), .CLK(clk), .Q(reg_file[61]) );
  DFFPOSX1 reg_file_reg_0__62_ ( .D(n25066), .CLK(clk), .Q(reg_file[62]) );
  DFFPOSX1 reg_file_reg_0__63_ ( .D(n25065), .CLK(clk), .Q(reg_file[63]) );
  DFFPOSX1 reg_file_reg_0__64_ ( .D(n25064), .CLK(clk), .Q(reg_file[64]) );
  DFFPOSX1 reg_file_reg_0__65_ ( .D(n25063), .CLK(clk), .Q(reg_file[65]) );
  DFFPOSX1 reg_file_reg_0__66_ ( .D(n25062), .CLK(clk), .Q(reg_file[66]) );
  DFFPOSX1 reg_file_reg_0__67_ ( .D(n25061), .CLK(clk), .Q(reg_file[67]) );
  DFFPOSX1 reg_file_reg_0__68_ ( .D(n25060), .CLK(clk), .Q(reg_file[68]) );
  DFFPOSX1 reg_file_reg_0__69_ ( .D(n25059), .CLK(clk), .Q(reg_file[69]) );
  DFFPOSX1 reg_file_reg_0__70_ ( .D(n25058), .CLK(clk), .Q(reg_file[70]) );
  DFFPOSX1 reg_file_reg_0__71_ ( .D(n25057), .CLK(clk), .Q(reg_file[71]) );
  DFFPOSX1 reg_file_reg_0__72_ ( .D(n25056), .CLK(clk), .Q(reg_file[72]) );
  DFFPOSX1 reg_file_reg_0__73_ ( .D(n25055), .CLK(clk), .Q(reg_file[73]) );
  DFFPOSX1 reg_file_reg_0__74_ ( .D(n25054), .CLK(clk), .Q(reg_file[74]) );
  DFFPOSX1 reg_file_reg_0__75_ ( .D(n25053), .CLK(clk), .Q(reg_file[75]) );
  DFFPOSX1 reg_file_reg_0__76_ ( .D(n25052), .CLK(clk), .Q(reg_file[76]) );
  DFFPOSX1 reg_file_reg_0__77_ ( .D(n25051), .CLK(clk), .Q(reg_file[77]) );
  DFFPOSX1 reg_file_reg_0__78_ ( .D(n25050), .CLK(clk), .Q(reg_file[78]) );
  DFFPOSX1 reg_file_reg_0__79_ ( .D(n25049), .CLK(clk), .Q(reg_file[79]) );
  DFFPOSX1 reg_file_reg_0__80_ ( .D(n25048), .CLK(clk), .Q(reg_file[80]) );
  DFFPOSX1 reg_file_reg_0__81_ ( .D(n25047), .CLK(clk), .Q(reg_file[81]) );
  DFFPOSX1 reg_file_reg_0__82_ ( .D(n25046), .CLK(clk), .Q(reg_file[82]) );
  DFFPOSX1 reg_file_reg_0__83_ ( .D(n25045), .CLK(clk), .Q(reg_file[83]) );
  DFFPOSX1 reg_file_reg_0__84_ ( .D(n25044), .CLK(clk), .Q(reg_file[84]) );
  DFFPOSX1 reg_file_reg_0__85_ ( .D(n25043), .CLK(clk), .Q(reg_file[85]) );
  DFFPOSX1 reg_file_reg_0__86_ ( .D(n25042), .CLK(clk), .Q(reg_file[86]) );
  DFFPOSX1 reg_file_reg_0__87_ ( .D(n25041), .CLK(clk), .Q(reg_file[87]) );
  DFFPOSX1 reg_file_reg_0__88_ ( .D(n25040), .CLK(clk), .Q(reg_file[88]) );
  DFFPOSX1 reg_file_reg_0__89_ ( .D(n25039), .CLK(clk), .Q(reg_file[89]) );
  DFFPOSX1 reg_file_reg_0__90_ ( .D(n25038), .CLK(clk), .Q(reg_file[90]) );
  DFFPOSX1 reg_file_reg_0__91_ ( .D(n25037), .CLK(clk), .Q(reg_file[91]) );
  DFFPOSX1 reg_file_reg_0__92_ ( .D(n25036), .CLK(clk), .Q(reg_file[92]) );
  DFFPOSX1 reg_file_reg_0__93_ ( .D(n25035), .CLK(clk), .Q(reg_file[93]) );
  DFFPOSX1 reg_file_reg_0__94_ ( .D(n25034), .CLK(clk), .Q(reg_file[94]) );
  DFFPOSX1 reg_file_reg_0__95_ ( .D(n25033), .CLK(clk), .Q(reg_file[95]) );
  DFFPOSX1 reg_file_reg_0__96_ ( .D(n25032), .CLK(clk), .Q(reg_file[96]) );
  DFFPOSX1 reg_file_reg_0__97_ ( .D(n25031), .CLK(clk), .Q(reg_file[97]) );
  DFFPOSX1 reg_file_reg_0__98_ ( .D(n25030), .CLK(clk), .Q(reg_file[98]) );
  DFFPOSX1 reg_file_reg_0__99_ ( .D(n25029), .CLK(clk), .Q(reg_file[99]) );
  DFFPOSX1 reg_file_reg_0__100_ ( .D(n25028), .CLK(clk), .Q(reg_file[100]) );
  DFFPOSX1 reg_file_reg_0__101_ ( .D(n25027), .CLK(clk), .Q(reg_file[101]) );
  DFFPOSX1 reg_file_reg_0__102_ ( .D(n25026), .CLK(clk), .Q(reg_file[102]) );
  DFFPOSX1 reg_file_reg_0__103_ ( .D(n25025), .CLK(clk), .Q(reg_file[103]) );
  DFFPOSX1 reg_file_reg_0__104_ ( .D(n25024), .CLK(clk), .Q(reg_file[104]) );
  DFFPOSX1 reg_file_reg_0__105_ ( .D(n25023), .CLK(clk), .Q(reg_file[105]) );
  DFFPOSX1 reg_file_reg_0__106_ ( .D(n25022), .CLK(clk), .Q(reg_file[106]) );
  DFFPOSX1 reg_file_reg_0__107_ ( .D(n25021), .CLK(clk), .Q(reg_file[107]) );
  DFFPOSX1 reg_file_reg_0__108_ ( .D(n25020), .CLK(clk), .Q(reg_file[108]) );
  DFFPOSX1 reg_file_reg_0__109_ ( .D(n25019), .CLK(clk), .Q(reg_file[109]) );
  DFFPOSX1 reg_file_reg_0__110_ ( .D(n25018), .CLK(clk), .Q(reg_file[110]) );
  DFFPOSX1 reg_file_reg_0__111_ ( .D(n25017), .CLK(clk), .Q(reg_file[111]) );
  DFFPOSX1 reg_file_reg_0__112_ ( .D(n25016), .CLK(clk), .Q(reg_file[112]) );
  DFFPOSX1 reg_file_reg_0__113_ ( .D(n25015), .CLK(clk), .Q(reg_file[113]) );
  DFFPOSX1 reg_file_reg_0__114_ ( .D(n25014), .CLK(clk), .Q(reg_file[114]) );
  DFFPOSX1 reg_file_reg_0__115_ ( .D(n25013), .CLK(clk), .Q(reg_file[115]) );
  DFFPOSX1 reg_file_reg_0__116_ ( .D(n25012), .CLK(clk), .Q(reg_file[116]) );
  DFFPOSX1 reg_file_reg_0__117_ ( .D(n25011), .CLK(clk), .Q(reg_file[117]) );
  DFFPOSX1 reg_file_reg_0__118_ ( .D(n25010), .CLK(clk), .Q(reg_file[118]) );
  DFFPOSX1 reg_file_reg_0__119_ ( .D(n25009), .CLK(clk), .Q(reg_file[119]) );
  DFFPOSX1 reg_file_reg_0__120_ ( .D(n25008), .CLK(clk), .Q(reg_file[120]) );
  DFFPOSX1 reg_file_reg_0__121_ ( .D(n25007), .CLK(clk), .Q(reg_file[121]) );
  DFFPOSX1 reg_file_reg_0__122_ ( .D(n25006), .CLK(clk), .Q(reg_file[122]) );
  DFFPOSX1 reg_file_reg_0__123_ ( .D(n25005), .CLK(clk), .Q(reg_file[123]) );
  DFFPOSX1 reg_file_reg_0__124_ ( .D(n25004), .CLK(clk), .Q(reg_file[124]) );
  DFFPOSX1 reg_file_reg_0__125_ ( .D(n25003), .CLK(clk), .Q(reg_file[125]) );
  DFFPOSX1 reg_file_reg_0__126_ ( .D(n25002), .CLK(clk), .Q(reg_file[126]) );
  DFFPOSX1 reg_file_reg_0__127_ ( .D(n25001), .CLK(clk), .Q(reg_file[127]) );
  DFFPOSX1 reg_file_reg_1__0_ ( .D(n25000), .CLK(clk), .Q(reg_file[128]) );
  DFFPOSX1 reg_file_reg_1__1_ ( .D(n24999), .CLK(clk), .Q(reg_file[129]) );
  DFFPOSX1 reg_file_reg_1__2_ ( .D(n24998), .CLK(clk), .Q(reg_file[130]) );
  DFFPOSX1 reg_file_reg_1__3_ ( .D(n24997), .CLK(clk), .Q(reg_file[131]) );
  DFFPOSX1 reg_file_reg_1__4_ ( .D(n24996), .CLK(clk), .Q(reg_file[132]) );
  DFFPOSX1 reg_file_reg_1__5_ ( .D(n24995), .CLK(clk), .Q(reg_file[133]) );
  DFFPOSX1 reg_file_reg_1__6_ ( .D(n24994), .CLK(clk), .Q(reg_file[134]) );
  DFFPOSX1 reg_file_reg_1__7_ ( .D(n24993), .CLK(clk), .Q(reg_file[135]) );
  DFFPOSX1 reg_file_reg_1__8_ ( .D(n24992), .CLK(clk), .Q(reg_file[136]) );
  DFFPOSX1 reg_file_reg_1__9_ ( .D(n24991), .CLK(clk), .Q(reg_file[137]) );
  DFFPOSX1 reg_file_reg_1__10_ ( .D(n24990), .CLK(clk), .Q(reg_file[138]) );
  DFFPOSX1 reg_file_reg_1__11_ ( .D(n24989), .CLK(clk), .Q(reg_file[139]) );
  DFFPOSX1 reg_file_reg_1__12_ ( .D(n24988), .CLK(clk), .Q(reg_file[140]) );
  DFFPOSX1 reg_file_reg_1__13_ ( .D(n24987), .CLK(clk), .Q(reg_file[141]) );
  DFFPOSX1 reg_file_reg_1__14_ ( .D(n24986), .CLK(clk), .Q(reg_file[142]) );
  DFFPOSX1 reg_file_reg_1__15_ ( .D(n24985), .CLK(clk), .Q(reg_file[143]) );
  DFFPOSX1 reg_file_reg_1__16_ ( .D(n24984), .CLK(clk), .Q(reg_file[144]) );
  DFFPOSX1 reg_file_reg_1__17_ ( .D(n24983), .CLK(clk), .Q(reg_file[145]) );
  DFFPOSX1 reg_file_reg_1__18_ ( .D(n24982), .CLK(clk), .Q(reg_file[146]) );
  DFFPOSX1 reg_file_reg_1__19_ ( .D(n24981), .CLK(clk), .Q(reg_file[147]) );
  DFFPOSX1 reg_file_reg_1__20_ ( .D(n24980), .CLK(clk), .Q(reg_file[148]) );
  DFFPOSX1 reg_file_reg_1__21_ ( .D(n24979), .CLK(clk), .Q(reg_file[149]) );
  DFFPOSX1 reg_file_reg_1__22_ ( .D(n24978), .CLK(clk), .Q(reg_file[150]) );
  DFFPOSX1 reg_file_reg_1__23_ ( .D(n24977), .CLK(clk), .Q(reg_file[151]) );
  DFFPOSX1 reg_file_reg_1__24_ ( .D(n24976), .CLK(clk), .Q(reg_file[152]) );
  DFFPOSX1 reg_file_reg_1__25_ ( .D(n24975), .CLK(clk), .Q(reg_file[153]) );
  DFFPOSX1 reg_file_reg_1__26_ ( .D(n24974), .CLK(clk), .Q(reg_file[154]) );
  DFFPOSX1 reg_file_reg_1__27_ ( .D(n24973), .CLK(clk), .Q(reg_file[155]) );
  DFFPOSX1 reg_file_reg_1__28_ ( .D(n24972), .CLK(clk), .Q(reg_file[156]) );
  DFFPOSX1 reg_file_reg_1__29_ ( .D(n24971), .CLK(clk), .Q(reg_file[157]) );
  DFFPOSX1 reg_file_reg_1__30_ ( .D(n24970), .CLK(clk), .Q(reg_file[158]) );
  DFFPOSX1 reg_file_reg_1__31_ ( .D(n24969), .CLK(clk), .Q(reg_file[159]) );
  DFFPOSX1 reg_file_reg_1__32_ ( .D(n24968), .CLK(clk), .Q(reg_file[160]) );
  DFFPOSX1 reg_file_reg_1__33_ ( .D(n24967), .CLK(clk), .Q(reg_file[161]) );
  DFFPOSX1 reg_file_reg_1__34_ ( .D(n24966), .CLK(clk), .Q(reg_file[162]) );
  DFFPOSX1 reg_file_reg_1__35_ ( .D(n24965), .CLK(clk), .Q(reg_file[163]) );
  DFFPOSX1 reg_file_reg_1__36_ ( .D(n24964), .CLK(clk), .Q(reg_file[164]) );
  DFFPOSX1 reg_file_reg_1__37_ ( .D(n24963), .CLK(clk), .Q(reg_file[165]) );
  DFFPOSX1 reg_file_reg_1__38_ ( .D(n24962), .CLK(clk), .Q(reg_file[166]) );
  DFFPOSX1 reg_file_reg_1__39_ ( .D(n24961), .CLK(clk), .Q(reg_file[167]) );
  DFFPOSX1 reg_file_reg_1__40_ ( .D(n24960), .CLK(clk), .Q(reg_file[168]) );
  DFFPOSX1 reg_file_reg_1__41_ ( .D(n24959), .CLK(clk), .Q(reg_file[169]) );
  DFFPOSX1 reg_file_reg_1__42_ ( .D(n24958), .CLK(clk), .Q(reg_file[170]) );
  DFFPOSX1 reg_file_reg_1__43_ ( .D(n24957), .CLK(clk), .Q(reg_file[171]) );
  DFFPOSX1 reg_file_reg_1__44_ ( .D(n24956), .CLK(clk), .Q(reg_file[172]) );
  DFFPOSX1 reg_file_reg_1__45_ ( .D(n24955), .CLK(clk), .Q(reg_file[173]) );
  DFFPOSX1 reg_file_reg_1__46_ ( .D(n24954), .CLK(clk), .Q(reg_file[174]) );
  DFFPOSX1 reg_file_reg_1__47_ ( .D(n24953), .CLK(clk), .Q(reg_file[175]) );
  DFFPOSX1 reg_file_reg_1__48_ ( .D(n24952), .CLK(clk), .Q(reg_file[176]) );
  DFFPOSX1 reg_file_reg_1__49_ ( .D(n24951), .CLK(clk), .Q(reg_file[177]) );
  DFFPOSX1 reg_file_reg_1__50_ ( .D(n24950), .CLK(clk), .Q(reg_file[178]) );
  DFFPOSX1 reg_file_reg_1__51_ ( .D(n24949), .CLK(clk), .Q(reg_file[179]) );
  DFFPOSX1 reg_file_reg_1__52_ ( .D(n24948), .CLK(clk), .Q(reg_file[180]) );
  DFFPOSX1 reg_file_reg_1__53_ ( .D(n24947), .CLK(clk), .Q(reg_file[181]) );
  DFFPOSX1 reg_file_reg_1__54_ ( .D(n24946), .CLK(clk), .Q(reg_file[182]) );
  DFFPOSX1 reg_file_reg_1__55_ ( .D(n24945), .CLK(clk), .Q(reg_file[183]) );
  DFFPOSX1 reg_file_reg_1__56_ ( .D(n24944), .CLK(clk), .Q(reg_file[184]) );
  DFFPOSX1 reg_file_reg_1__57_ ( .D(n24943), .CLK(clk), .Q(reg_file[185]) );
  DFFPOSX1 reg_file_reg_1__58_ ( .D(n24942), .CLK(clk), .Q(reg_file[186]) );
  DFFPOSX1 reg_file_reg_1__59_ ( .D(n24941), .CLK(clk), .Q(reg_file[187]) );
  DFFPOSX1 reg_file_reg_1__60_ ( .D(n24940), .CLK(clk), .Q(reg_file[188]) );
  DFFPOSX1 reg_file_reg_1__61_ ( .D(n24939), .CLK(clk), .Q(reg_file[189]) );
  DFFPOSX1 reg_file_reg_1__62_ ( .D(n24938), .CLK(clk), .Q(reg_file[190]) );
  DFFPOSX1 reg_file_reg_1__63_ ( .D(n24937), .CLK(clk), .Q(reg_file[191]) );
  DFFPOSX1 reg_file_reg_1__64_ ( .D(n24936), .CLK(clk), .Q(reg_file[192]) );
  DFFPOSX1 reg_file_reg_1__65_ ( .D(n24935), .CLK(clk), .Q(reg_file[193]) );
  DFFPOSX1 reg_file_reg_1__66_ ( .D(n24934), .CLK(clk), .Q(reg_file[194]) );
  DFFPOSX1 reg_file_reg_1__67_ ( .D(n24933), .CLK(clk), .Q(reg_file[195]) );
  DFFPOSX1 reg_file_reg_1__68_ ( .D(n24932), .CLK(clk), .Q(reg_file[196]) );
  DFFPOSX1 reg_file_reg_1__69_ ( .D(n24931), .CLK(clk), .Q(reg_file[197]) );
  DFFPOSX1 reg_file_reg_1__70_ ( .D(n24930), .CLK(clk), .Q(reg_file[198]) );
  DFFPOSX1 reg_file_reg_1__71_ ( .D(n24929), .CLK(clk), .Q(reg_file[199]) );
  DFFPOSX1 reg_file_reg_1__72_ ( .D(n24928), .CLK(clk), .Q(reg_file[200]) );
  DFFPOSX1 reg_file_reg_1__73_ ( .D(n24927), .CLK(clk), .Q(reg_file[201]) );
  DFFPOSX1 reg_file_reg_1__74_ ( .D(n24926), .CLK(clk), .Q(reg_file[202]) );
  DFFPOSX1 reg_file_reg_1__75_ ( .D(n24925), .CLK(clk), .Q(reg_file[203]) );
  DFFPOSX1 reg_file_reg_1__76_ ( .D(n24924), .CLK(clk), .Q(reg_file[204]) );
  DFFPOSX1 reg_file_reg_1__77_ ( .D(n24923), .CLK(clk), .Q(reg_file[205]) );
  DFFPOSX1 reg_file_reg_1__78_ ( .D(n24922), .CLK(clk), .Q(reg_file[206]) );
  DFFPOSX1 reg_file_reg_1__79_ ( .D(n24921), .CLK(clk), .Q(reg_file[207]) );
  DFFPOSX1 reg_file_reg_1__80_ ( .D(n24920), .CLK(clk), .Q(reg_file[208]) );
  DFFPOSX1 reg_file_reg_1__81_ ( .D(n24919), .CLK(clk), .Q(reg_file[209]) );
  DFFPOSX1 reg_file_reg_1__82_ ( .D(n24918), .CLK(clk), .Q(reg_file[210]) );
  DFFPOSX1 reg_file_reg_1__83_ ( .D(n24917), .CLK(clk), .Q(reg_file[211]) );
  DFFPOSX1 reg_file_reg_1__84_ ( .D(n24916), .CLK(clk), .Q(reg_file[212]) );
  DFFPOSX1 reg_file_reg_1__85_ ( .D(n24915), .CLK(clk), .Q(reg_file[213]) );
  DFFPOSX1 reg_file_reg_1__86_ ( .D(n24914), .CLK(clk), .Q(reg_file[214]) );
  DFFPOSX1 reg_file_reg_1__87_ ( .D(n24913), .CLK(clk), .Q(reg_file[215]) );
  DFFPOSX1 reg_file_reg_1__88_ ( .D(n24912), .CLK(clk), .Q(reg_file[216]) );
  DFFPOSX1 reg_file_reg_1__89_ ( .D(n24911), .CLK(clk), .Q(reg_file[217]) );
  DFFPOSX1 reg_file_reg_1__90_ ( .D(n24910), .CLK(clk), .Q(reg_file[218]) );
  DFFPOSX1 reg_file_reg_1__91_ ( .D(n24909), .CLK(clk), .Q(reg_file[219]) );
  DFFPOSX1 reg_file_reg_1__92_ ( .D(n24908), .CLK(clk), .Q(reg_file[220]) );
  DFFPOSX1 reg_file_reg_1__93_ ( .D(n24907), .CLK(clk), .Q(reg_file[221]) );
  DFFPOSX1 reg_file_reg_1__94_ ( .D(n24906), .CLK(clk), .Q(reg_file[222]) );
  DFFPOSX1 reg_file_reg_1__95_ ( .D(n24905), .CLK(clk), .Q(reg_file[223]) );
  DFFPOSX1 reg_file_reg_1__96_ ( .D(n24904), .CLK(clk), .Q(reg_file[224]) );
  DFFPOSX1 reg_file_reg_1__97_ ( .D(n24903), .CLK(clk), .Q(reg_file[225]) );
  DFFPOSX1 reg_file_reg_1__98_ ( .D(n24902), .CLK(clk), .Q(reg_file[226]) );
  DFFPOSX1 reg_file_reg_1__99_ ( .D(n24901), .CLK(clk), .Q(reg_file[227]) );
  DFFPOSX1 reg_file_reg_1__100_ ( .D(n24900), .CLK(clk), .Q(reg_file[228]) );
  DFFPOSX1 reg_file_reg_1__101_ ( .D(n24899), .CLK(clk), .Q(reg_file[229]) );
  DFFPOSX1 reg_file_reg_1__102_ ( .D(n24898), .CLK(clk), .Q(reg_file[230]) );
  DFFPOSX1 reg_file_reg_1__103_ ( .D(n24897), .CLK(clk), .Q(reg_file[231]) );
  DFFPOSX1 reg_file_reg_1__104_ ( .D(n24896), .CLK(clk), .Q(reg_file[232]) );
  DFFPOSX1 reg_file_reg_1__105_ ( .D(n24895), .CLK(clk), .Q(reg_file[233]) );
  DFFPOSX1 reg_file_reg_1__106_ ( .D(n24894), .CLK(clk), .Q(reg_file[234]) );
  DFFPOSX1 reg_file_reg_1__107_ ( .D(n24893), .CLK(clk), .Q(reg_file[235]) );
  DFFPOSX1 reg_file_reg_1__108_ ( .D(n24892), .CLK(clk), .Q(reg_file[236]) );
  DFFPOSX1 reg_file_reg_1__109_ ( .D(n24891), .CLK(clk), .Q(reg_file[237]) );
  DFFPOSX1 reg_file_reg_1__110_ ( .D(n24890), .CLK(clk), .Q(reg_file[238]) );
  DFFPOSX1 reg_file_reg_1__111_ ( .D(n24889), .CLK(clk), .Q(reg_file[239]) );
  DFFPOSX1 reg_file_reg_1__112_ ( .D(n24888), .CLK(clk), .Q(reg_file[240]) );
  DFFPOSX1 reg_file_reg_1__113_ ( .D(n24887), .CLK(clk), .Q(reg_file[241]) );
  DFFPOSX1 reg_file_reg_1__114_ ( .D(n24886), .CLK(clk), .Q(reg_file[242]) );
  DFFPOSX1 reg_file_reg_1__115_ ( .D(n24885), .CLK(clk), .Q(reg_file[243]) );
  DFFPOSX1 reg_file_reg_1__116_ ( .D(n24884), .CLK(clk), .Q(reg_file[244]) );
  DFFPOSX1 reg_file_reg_1__117_ ( .D(n24883), .CLK(clk), .Q(reg_file[245]) );
  DFFPOSX1 reg_file_reg_1__118_ ( .D(n24882), .CLK(clk), .Q(reg_file[246]) );
  DFFPOSX1 reg_file_reg_1__119_ ( .D(n24881), .CLK(clk), .Q(reg_file[247]) );
  DFFPOSX1 reg_file_reg_1__120_ ( .D(n24880), .CLK(clk), .Q(reg_file[248]) );
  DFFPOSX1 reg_file_reg_1__121_ ( .D(n24879), .CLK(clk), .Q(reg_file[249]) );
  DFFPOSX1 reg_file_reg_1__122_ ( .D(n24878), .CLK(clk), .Q(reg_file[250]) );
  DFFPOSX1 reg_file_reg_1__123_ ( .D(n24877), .CLK(clk), .Q(reg_file[251]) );
  DFFPOSX1 reg_file_reg_1__124_ ( .D(n24876), .CLK(clk), .Q(reg_file[252]) );
  DFFPOSX1 reg_file_reg_1__125_ ( .D(n24875), .CLK(clk), .Q(reg_file[253]) );
  DFFPOSX1 reg_file_reg_1__126_ ( .D(n24874), .CLK(clk), .Q(reg_file[254]) );
  DFFPOSX1 reg_file_reg_1__127_ ( .D(n24873), .CLK(clk), .Q(reg_file[255]) );
  DFFPOSX1 reg_file_reg_2__0_ ( .D(n24872), .CLK(clk), .Q(reg_file[256]) );
  DFFPOSX1 reg_file_reg_2__1_ ( .D(n24871), .CLK(clk), .Q(reg_file[257]) );
  DFFPOSX1 reg_file_reg_2__2_ ( .D(n24870), .CLK(clk), .Q(reg_file[258]) );
  DFFPOSX1 reg_file_reg_2__3_ ( .D(n24869), .CLK(clk), .Q(reg_file[259]) );
  DFFPOSX1 reg_file_reg_2__4_ ( .D(n24868), .CLK(clk), .Q(reg_file[260]) );
  DFFPOSX1 reg_file_reg_2__5_ ( .D(n24867), .CLK(clk), .Q(reg_file[261]) );
  DFFPOSX1 reg_file_reg_2__6_ ( .D(n24866), .CLK(clk), .Q(reg_file[262]) );
  DFFPOSX1 reg_file_reg_2__7_ ( .D(n24865), .CLK(clk), .Q(reg_file[263]) );
  DFFPOSX1 reg_file_reg_2__8_ ( .D(n24864), .CLK(clk), .Q(reg_file[264]) );
  DFFPOSX1 reg_file_reg_2__9_ ( .D(n24863), .CLK(clk), .Q(reg_file[265]) );
  DFFPOSX1 reg_file_reg_2__10_ ( .D(n24862), .CLK(clk), .Q(reg_file[266]) );
  DFFPOSX1 reg_file_reg_2__11_ ( .D(n24861), .CLK(clk), .Q(reg_file[267]) );
  DFFPOSX1 reg_file_reg_2__12_ ( .D(n24860), .CLK(clk), .Q(reg_file[268]) );
  DFFPOSX1 reg_file_reg_2__13_ ( .D(n24859), .CLK(clk), .Q(reg_file[269]) );
  DFFPOSX1 reg_file_reg_2__14_ ( .D(n24858), .CLK(clk), .Q(reg_file[270]) );
  DFFPOSX1 reg_file_reg_2__15_ ( .D(n24857), .CLK(clk), .Q(reg_file[271]) );
  DFFPOSX1 reg_file_reg_2__16_ ( .D(n24856), .CLK(clk), .Q(reg_file[272]) );
  DFFPOSX1 reg_file_reg_2__17_ ( .D(n24855), .CLK(clk), .Q(reg_file[273]) );
  DFFPOSX1 reg_file_reg_2__18_ ( .D(n24854), .CLK(clk), .Q(reg_file[274]) );
  DFFPOSX1 reg_file_reg_2__19_ ( .D(n24853), .CLK(clk), .Q(reg_file[275]) );
  DFFPOSX1 reg_file_reg_2__20_ ( .D(n24852), .CLK(clk), .Q(reg_file[276]) );
  DFFPOSX1 reg_file_reg_2__21_ ( .D(n24851), .CLK(clk), .Q(reg_file[277]) );
  DFFPOSX1 reg_file_reg_2__22_ ( .D(n24850), .CLK(clk), .Q(reg_file[278]) );
  DFFPOSX1 reg_file_reg_2__23_ ( .D(n24849), .CLK(clk), .Q(reg_file[279]) );
  DFFPOSX1 reg_file_reg_2__24_ ( .D(n24848), .CLK(clk), .Q(reg_file[280]) );
  DFFPOSX1 reg_file_reg_2__25_ ( .D(n24847), .CLK(clk), .Q(reg_file[281]) );
  DFFPOSX1 reg_file_reg_2__26_ ( .D(n24846), .CLK(clk), .Q(reg_file[282]) );
  DFFPOSX1 reg_file_reg_2__27_ ( .D(n24845), .CLK(clk), .Q(reg_file[283]) );
  DFFPOSX1 reg_file_reg_2__28_ ( .D(n24844), .CLK(clk), .Q(reg_file[284]) );
  DFFPOSX1 reg_file_reg_2__29_ ( .D(n24843), .CLK(clk), .Q(reg_file[285]) );
  DFFPOSX1 reg_file_reg_2__30_ ( .D(n24842), .CLK(clk), .Q(reg_file[286]) );
  DFFPOSX1 reg_file_reg_2__31_ ( .D(n24841), .CLK(clk), .Q(reg_file[287]) );
  DFFPOSX1 reg_file_reg_2__32_ ( .D(n24840), .CLK(clk), .Q(reg_file[288]) );
  DFFPOSX1 reg_file_reg_2__33_ ( .D(n24839), .CLK(clk), .Q(reg_file[289]) );
  DFFPOSX1 reg_file_reg_2__34_ ( .D(n24838), .CLK(clk), .Q(reg_file[290]) );
  DFFPOSX1 reg_file_reg_2__35_ ( .D(n24837), .CLK(clk), .Q(reg_file[291]) );
  DFFPOSX1 reg_file_reg_2__36_ ( .D(n24836), .CLK(clk), .Q(reg_file[292]) );
  DFFPOSX1 reg_file_reg_2__37_ ( .D(n24835), .CLK(clk), .Q(reg_file[293]) );
  DFFPOSX1 reg_file_reg_2__38_ ( .D(n24834), .CLK(clk), .Q(reg_file[294]) );
  DFFPOSX1 reg_file_reg_2__39_ ( .D(n24833), .CLK(clk), .Q(reg_file[295]) );
  DFFPOSX1 reg_file_reg_2__40_ ( .D(n24832), .CLK(clk), .Q(reg_file[296]) );
  DFFPOSX1 reg_file_reg_2__41_ ( .D(n24831), .CLK(clk), .Q(reg_file[297]) );
  DFFPOSX1 reg_file_reg_2__42_ ( .D(n24830), .CLK(clk), .Q(reg_file[298]) );
  DFFPOSX1 reg_file_reg_2__43_ ( .D(n24829), .CLK(clk), .Q(reg_file[299]) );
  DFFPOSX1 reg_file_reg_2__44_ ( .D(n24828), .CLK(clk), .Q(reg_file[300]) );
  DFFPOSX1 reg_file_reg_2__45_ ( .D(n24827), .CLK(clk), .Q(reg_file[301]) );
  DFFPOSX1 reg_file_reg_2__46_ ( .D(n24826), .CLK(clk), .Q(reg_file[302]) );
  DFFPOSX1 reg_file_reg_2__47_ ( .D(n24825), .CLK(clk), .Q(reg_file[303]) );
  DFFPOSX1 reg_file_reg_2__48_ ( .D(n24824), .CLK(clk), .Q(reg_file[304]) );
  DFFPOSX1 reg_file_reg_2__49_ ( .D(n24823), .CLK(clk), .Q(reg_file[305]) );
  DFFPOSX1 reg_file_reg_2__50_ ( .D(n24822), .CLK(clk), .Q(reg_file[306]) );
  DFFPOSX1 reg_file_reg_2__51_ ( .D(n24821), .CLK(clk), .Q(reg_file[307]) );
  DFFPOSX1 reg_file_reg_2__52_ ( .D(n24820), .CLK(clk), .Q(reg_file[308]) );
  DFFPOSX1 reg_file_reg_2__53_ ( .D(n24819), .CLK(clk), .Q(reg_file[309]) );
  DFFPOSX1 reg_file_reg_2__54_ ( .D(n24818), .CLK(clk), .Q(reg_file[310]) );
  DFFPOSX1 reg_file_reg_2__55_ ( .D(n24817), .CLK(clk), .Q(reg_file[311]) );
  DFFPOSX1 reg_file_reg_2__56_ ( .D(n24816), .CLK(clk), .Q(reg_file[312]) );
  DFFPOSX1 reg_file_reg_2__57_ ( .D(n24815), .CLK(clk), .Q(reg_file[313]) );
  DFFPOSX1 reg_file_reg_2__58_ ( .D(n24814), .CLK(clk), .Q(reg_file[314]) );
  DFFPOSX1 reg_file_reg_2__59_ ( .D(n24813), .CLK(clk), .Q(reg_file[315]) );
  DFFPOSX1 reg_file_reg_2__60_ ( .D(n24812), .CLK(clk), .Q(reg_file[316]) );
  DFFPOSX1 reg_file_reg_2__61_ ( .D(n24811), .CLK(clk), .Q(reg_file[317]) );
  DFFPOSX1 reg_file_reg_2__62_ ( .D(n24810), .CLK(clk), .Q(reg_file[318]) );
  DFFPOSX1 reg_file_reg_2__63_ ( .D(n24809), .CLK(clk), .Q(reg_file[319]) );
  DFFPOSX1 reg_file_reg_2__64_ ( .D(n24808), .CLK(clk), .Q(reg_file[320]) );
  DFFPOSX1 reg_file_reg_2__65_ ( .D(n24807), .CLK(clk), .Q(reg_file[321]) );
  DFFPOSX1 reg_file_reg_2__66_ ( .D(n24806), .CLK(clk), .Q(reg_file[322]) );
  DFFPOSX1 reg_file_reg_2__67_ ( .D(n24805), .CLK(clk), .Q(reg_file[323]) );
  DFFPOSX1 reg_file_reg_2__68_ ( .D(n24804), .CLK(clk), .Q(reg_file[324]) );
  DFFPOSX1 reg_file_reg_2__69_ ( .D(n24803), .CLK(clk), .Q(reg_file[325]) );
  DFFPOSX1 reg_file_reg_2__70_ ( .D(n24802), .CLK(clk), .Q(reg_file[326]) );
  DFFPOSX1 reg_file_reg_2__71_ ( .D(n24801), .CLK(clk), .Q(reg_file[327]) );
  DFFPOSX1 reg_file_reg_2__72_ ( .D(n24800), .CLK(clk), .Q(reg_file[328]) );
  DFFPOSX1 reg_file_reg_2__73_ ( .D(n24799), .CLK(clk), .Q(reg_file[329]) );
  DFFPOSX1 reg_file_reg_2__74_ ( .D(n24798), .CLK(clk), .Q(reg_file[330]) );
  DFFPOSX1 reg_file_reg_2__75_ ( .D(n24797), .CLK(clk), .Q(reg_file[331]) );
  DFFPOSX1 reg_file_reg_2__76_ ( .D(n24796), .CLK(clk), .Q(reg_file[332]) );
  DFFPOSX1 reg_file_reg_2__77_ ( .D(n24795), .CLK(clk), .Q(reg_file[333]) );
  DFFPOSX1 reg_file_reg_2__78_ ( .D(n24794), .CLK(clk), .Q(reg_file[334]) );
  DFFPOSX1 reg_file_reg_2__79_ ( .D(n24793), .CLK(clk), .Q(reg_file[335]) );
  DFFPOSX1 reg_file_reg_2__80_ ( .D(n24792), .CLK(clk), .Q(reg_file[336]) );
  DFFPOSX1 reg_file_reg_2__81_ ( .D(n24791), .CLK(clk), .Q(reg_file[337]) );
  DFFPOSX1 reg_file_reg_2__82_ ( .D(n24790), .CLK(clk), .Q(reg_file[338]) );
  DFFPOSX1 reg_file_reg_2__83_ ( .D(n24789), .CLK(clk), .Q(reg_file[339]) );
  DFFPOSX1 reg_file_reg_2__84_ ( .D(n24788), .CLK(clk), .Q(reg_file[340]) );
  DFFPOSX1 reg_file_reg_2__85_ ( .D(n24787), .CLK(clk), .Q(reg_file[341]) );
  DFFPOSX1 reg_file_reg_2__86_ ( .D(n24786), .CLK(clk), .Q(reg_file[342]) );
  DFFPOSX1 reg_file_reg_2__87_ ( .D(n24785), .CLK(clk), .Q(reg_file[343]) );
  DFFPOSX1 reg_file_reg_2__88_ ( .D(n24784), .CLK(clk), .Q(reg_file[344]) );
  DFFPOSX1 reg_file_reg_2__89_ ( .D(n24783), .CLK(clk), .Q(reg_file[345]) );
  DFFPOSX1 reg_file_reg_2__90_ ( .D(n24782), .CLK(clk), .Q(reg_file[346]) );
  DFFPOSX1 reg_file_reg_2__91_ ( .D(n24781), .CLK(clk), .Q(reg_file[347]) );
  DFFPOSX1 reg_file_reg_2__92_ ( .D(n24780), .CLK(clk), .Q(reg_file[348]) );
  DFFPOSX1 reg_file_reg_2__93_ ( .D(n24779), .CLK(clk), .Q(reg_file[349]) );
  DFFPOSX1 reg_file_reg_2__94_ ( .D(n24778), .CLK(clk), .Q(reg_file[350]) );
  DFFPOSX1 reg_file_reg_2__95_ ( .D(n24777), .CLK(clk), .Q(reg_file[351]) );
  DFFPOSX1 reg_file_reg_2__96_ ( .D(n24776), .CLK(clk), .Q(reg_file[352]) );
  DFFPOSX1 reg_file_reg_2__97_ ( .D(n24775), .CLK(clk), .Q(reg_file[353]) );
  DFFPOSX1 reg_file_reg_2__98_ ( .D(n24774), .CLK(clk), .Q(reg_file[354]) );
  DFFPOSX1 reg_file_reg_2__99_ ( .D(n24773), .CLK(clk), .Q(reg_file[355]) );
  DFFPOSX1 reg_file_reg_2__100_ ( .D(n24772), .CLK(clk), .Q(reg_file[356]) );
  DFFPOSX1 reg_file_reg_2__101_ ( .D(n24771), .CLK(clk), .Q(reg_file[357]) );
  DFFPOSX1 reg_file_reg_2__102_ ( .D(n24770), .CLK(clk), .Q(reg_file[358]) );
  DFFPOSX1 reg_file_reg_2__103_ ( .D(n24769), .CLK(clk), .Q(reg_file[359]) );
  DFFPOSX1 reg_file_reg_2__104_ ( .D(n24768), .CLK(clk), .Q(reg_file[360]) );
  DFFPOSX1 reg_file_reg_2__105_ ( .D(n24767), .CLK(clk), .Q(reg_file[361]) );
  DFFPOSX1 reg_file_reg_2__106_ ( .D(n24766), .CLK(clk), .Q(reg_file[362]) );
  DFFPOSX1 reg_file_reg_2__107_ ( .D(n24765), .CLK(clk), .Q(reg_file[363]) );
  DFFPOSX1 reg_file_reg_2__108_ ( .D(n24764), .CLK(clk), .Q(reg_file[364]) );
  DFFPOSX1 reg_file_reg_2__109_ ( .D(n24763), .CLK(clk), .Q(reg_file[365]) );
  DFFPOSX1 reg_file_reg_2__110_ ( .D(n24762), .CLK(clk), .Q(reg_file[366]) );
  DFFPOSX1 reg_file_reg_2__111_ ( .D(n24761), .CLK(clk), .Q(reg_file[367]) );
  DFFPOSX1 reg_file_reg_2__112_ ( .D(n24760), .CLK(clk), .Q(reg_file[368]) );
  DFFPOSX1 reg_file_reg_2__113_ ( .D(n24759), .CLK(clk), .Q(reg_file[369]) );
  DFFPOSX1 reg_file_reg_2__114_ ( .D(n24758), .CLK(clk), .Q(reg_file[370]) );
  DFFPOSX1 reg_file_reg_2__115_ ( .D(n24757), .CLK(clk), .Q(reg_file[371]) );
  DFFPOSX1 reg_file_reg_2__116_ ( .D(n24756), .CLK(clk), .Q(reg_file[372]) );
  DFFPOSX1 reg_file_reg_2__117_ ( .D(n24755), .CLK(clk), .Q(reg_file[373]) );
  DFFPOSX1 reg_file_reg_2__118_ ( .D(n24754), .CLK(clk), .Q(reg_file[374]) );
  DFFPOSX1 reg_file_reg_2__119_ ( .D(n24753), .CLK(clk), .Q(reg_file[375]) );
  DFFPOSX1 reg_file_reg_2__120_ ( .D(n24752), .CLK(clk), .Q(reg_file[376]) );
  DFFPOSX1 reg_file_reg_2__121_ ( .D(n24751), .CLK(clk), .Q(reg_file[377]) );
  DFFPOSX1 reg_file_reg_2__122_ ( .D(n24750), .CLK(clk), .Q(reg_file[378]) );
  DFFPOSX1 reg_file_reg_2__123_ ( .D(n24749), .CLK(clk), .Q(reg_file[379]) );
  DFFPOSX1 reg_file_reg_2__124_ ( .D(n24748), .CLK(clk), .Q(reg_file[380]) );
  DFFPOSX1 reg_file_reg_2__125_ ( .D(n24747), .CLK(clk), .Q(reg_file[381]) );
  DFFPOSX1 reg_file_reg_2__126_ ( .D(n24746), .CLK(clk), .Q(reg_file[382]) );
  DFFPOSX1 reg_file_reg_2__127_ ( .D(n24745), .CLK(clk), .Q(reg_file[383]) );
  DFFPOSX1 reg_file_reg_3__0_ ( .D(n24744), .CLK(clk), .Q(reg_file[384]) );
  DFFPOSX1 reg_file_reg_3__1_ ( .D(n24743), .CLK(clk), .Q(reg_file[385]) );
  DFFPOSX1 reg_file_reg_3__2_ ( .D(n24742), .CLK(clk), .Q(reg_file[386]) );
  DFFPOSX1 reg_file_reg_3__3_ ( .D(n24741), .CLK(clk), .Q(reg_file[387]) );
  DFFPOSX1 reg_file_reg_3__4_ ( .D(n24740), .CLK(clk), .Q(reg_file[388]) );
  DFFPOSX1 reg_file_reg_3__5_ ( .D(n24739), .CLK(clk), .Q(reg_file[389]) );
  DFFPOSX1 reg_file_reg_3__6_ ( .D(n24738), .CLK(clk), .Q(reg_file[390]) );
  DFFPOSX1 reg_file_reg_3__7_ ( .D(n24737), .CLK(clk), .Q(reg_file[391]) );
  DFFPOSX1 reg_file_reg_3__8_ ( .D(n24736), .CLK(clk), .Q(reg_file[392]) );
  DFFPOSX1 reg_file_reg_3__9_ ( .D(n24735), .CLK(clk), .Q(reg_file[393]) );
  DFFPOSX1 reg_file_reg_3__10_ ( .D(n24734), .CLK(clk), .Q(reg_file[394]) );
  DFFPOSX1 reg_file_reg_3__11_ ( .D(n24733), .CLK(clk), .Q(reg_file[395]) );
  DFFPOSX1 reg_file_reg_3__12_ ( .D(n24732), .CLK(clk), .Q(reg_file[396]) );
  DFFPOSX1 reg_file_reg_3__13_ ( .D(n24731), .CLK(clk), .Q(reg_file[397]) );
  DFFPOSX1 reg_file_reg_3__14_ ( .D(n24730), .CLK(clk), .Q(reg_file[398]) );
  DFFPOSX1 reg_file_reg_3__15_ ( .D(n24729), .CLK(clk), .Q(reg_file[399]) );
  DFFPOSX1 reg_file_reg_3__16_ ( .D(n24728), .CLK(clk), .Q(reg_file[400]) );
  DFFPOSX1 reg_file_reg_3__17_ ( .D(n24727), .CLK(clk), .Q(reg_file[401]) );
  DFFPOSX1 reg_file_reg_3__18_ ( .D(n24726), .CLK(clk), .Q(reg_file[402]) );
  DFFPOSX1 reg_file_reg_3__19_ ( .D(n24725), .CLK(clk), .Q(reg_file[403]) );
  DFFPOSX1 reg_file_reg_3__20_ ( .D(n24724), .CLK(clk), .Q(reg_file[404]) );
  DFFPOSX1 reg_file_reg_3__21_ ( .D(n24723), .CLK(clk), .Q(reg_file[405]) );
  DFFPOSX1 reg_file_reg_3__22_ ( .D(n24722), .CLK(clk), .Q(reg_file[406]) );
  DFFPOSX1 reg_file_reg_3__23_ ( .D(n24721), .CLK(clk), .Q(reg_file[407]) );
  DFFPOSX1 reg_file_reg_3__24_ ( .D(n24720), .CLK(clk), .Q(reg_file[408]) );
  DFFPOSX1 reg_file_reg_3__25_ ( .D(n24719), .CLK(clk), .Q(reg_file[409]) );
  DFFPOSX1 reg_file_reg_3__26_ ( .D(n24718), .CLK(clk), .Q(reg_file[410]) );
  DFFPOSX1 reg_file_reg_3__27_ ( .D(n24717), .CLK(clk), .Q(reg_file[411]) );
  DFFPOSX1 reg_file_reg_3__28_ ( .D(n24716), .CLK(clk), .Q(reg_file[412]) );
  DFFPOSX1 reg_file_reg_3__29_ ( .D(n24715), .CLK(clk), .Q(reg_file[413]) );
  DFFPOSX1 reg_file_reg_3__30_ ( .D(n24714), .CLK(clk), .Q(reg_file[414]) );
  DFFPOSX1 reg_file_reg_3__31_ ( .D(n24713), .CLK(clk), .Q(reg_file[415]) );
  DFFPOSX1 reg_file_reg_3__32_ ( .D(n24712), .CLK(clk), .Q(reg_file[416]) );
  DFFPOSX1 reg_file_reg_3__33_ ( .D(n24711), .CLK(clk), .Q(reg_file[417]) );
  DFFPOSX1 reg_file_reg_3__34_ ( .D(n24710), .CLK(clk), .Q(reg_file[418]) );
  DFFPOSX1 reg_file_reg_3__35_ ( .D(n24709), .CLK(clk), .Q(reg_file[419]) );
  DFFPOSX1 reg_file_reg_3__36_ ( .D(n24708), .CLK(clk), .Q(reg_file[420]) );
  DFFPOSX1 reg_file_reg_3__37_ ( .D(n24707), .CLK(clk), .Q(reg_file[421]) );
  DFFPOSX1 reg_file_reg_3__38_ ( .D(n24706), .CLK(clk), .Q(reg_file[422]) );
  DFFPOSX1 reg_file_reg_3__39_ ( .D(n24705), .CLK(clk), .Q(reg_file[423]) );
  DFFPOSX1 reg_file_reg_3__40_ ( .D(n24704), .CLK(clk), .Q(reg_file[424]) );
  DFFPOSX1 reg_file_reg_3__41_ ( .D(n24703), .CLK(clk), .Q(reg_file[425]) );
  DFFPOSX1 reg_file_reg_3__42_ ( .D(n24702), .CLK(clk), .Q(reg_file[426]) );
  DFFPOSX1 reg_file_reg_3__43_ ( .D(n24701), .CLK(clk), .Q(reg_file[427]) );
  DFFPOSX1 reg_file_reg_3__44_ ( .D(n24700), .CLK(clk), .Q(reg_file[428]) );
  DFFPOSX1 reg_file_reg_3__45_ ( .D(n24699), .CLK(clk), .Q(reg_file[429]) );
  DFFPOSX1 reg_file_reg_3__46_ ( .D(n24698), .CLK(clk), .Q(reg_file[430]) );
  DFFPOSX1 reg_file_reg_3__47_ ( .D(n24697), .CLK(clk), .Q(reg_file[431]) );
  DFFPOSX1 reg_file_reg_3__48_ ( .D(n24696), .CLK(clk), .Q(reg_file[432]) );
  DFFPOSX1 reg_file_reg_3__49_ ( .D(n24695), .CLK(clk), .Q(reg_file[433]) );
  DFFPOSX1 reg_file_reg_3__50_ ( .D(n24694), .CLK(clk), .Q(reg_file[434]) );
  DFFPOSX1 reg_file_reg_3__51_ ( .D(n24693), .CLK(clk), .Q(reg_file[435]) );
  DFFPOSX1 reg_file_reg_3__52_ ( .D(n24692), .CLK(clk), .Q(reg_file[436]) );
  DFFPOSX1 reg_file_reg_3__53_ ( .D(n24691), .CLK(clk), .Q(reg_file[437]) );
  DFFPOSX1 reg_file_reg_3__54_ ( .D(n24690), .CLK(clk), .Q(reg_file[438]) );
  DFFPOSX1 reg_file_reg_3__55_ ( .D(n24689), .CLK(clk), .Q(reg_file[439]) );
  DFFPOSX1 reg_file_reg_3__56_ ( .D(n24688), .CLK(clk), .Q(reg_file[440]) );
  DFFPOSX1 reg_file_reg_3__57_ ( .D(n24687), .CLK(clk), .Q(reg_file[441]) );
  DFFPOSX1 reg_file_reg_3__58_ ( .D(n24686), .CLK(clk), .Q(reg_file[442]) );
  DFFPOSX1 reg_file_reg_3__59_ ( .D(n24685), .CLK(clk), .Q(reg_file[443]) );
  DFFPOSX1 reg_file_reg_3__60_ ( .D(n24684), .CLK(clk), .Q(reg_file[444]) );
  DFFPOSX1 reg_file_reg_3__61_ ( .D(n24683), .CLK(clk), .Q(reg_file[445]) );
  DFFPOSX1 reg_file_reg_3__62_ ( .D(n24682), .CLK(clk), .Q(reg_file[446]) );
  DFFPOSX1 reg_file_reg_3__63_ ( .D(n24681), .CLK(clk), .Q(reg_file[447]) );
  DFFPOSX1 reg_file_reg_3__64_ ( .D(n24680), .CLK(clk), .Q(reg_file[448]) );
  DFFPOSX1 reg_file_reg_3__65_ ( .D(n24679), .CLK(clk), .Q(reg_file[449]) );
  DFFPOSX1 reg_file_reg_3__66_ ( .D(n24678), .CLK(clk), .Q(reg_file[450]) );
  DFFPOSX1 reg_file_reg_3__67_ ( .D(n24677), .CLK(clk), .Q(reg_file[451]) );
  DFFPOSX1 reg_file_reg_3__68_ ( .D(n24676), .CLK(clk), .Q(reg_file[452]) );
  DFFPOSX1 reg_file_reg_3__69_ ( .D(n24675), .CLK(clk), .Q(reg_file[453]) );
  DFFPOSX1 reg_file_reg_3__70_ ( .D(n24674), .CLK(clk), .Q(reg_file[454]) );
  DFFPOSX1 reg_file_reg_3__71_ ( .D(n24673), .CLK(clk), .Q(reg_file[455]) );
  DFFPOSX1 reg_file_reg_3__72_ ( .D(n24672), .CLK(clk), .Q(reg_file[456]) );
  DFFPOSX1 reg_file_reg_3__73_ ( .D(n24671), .CLK(clk), .Q(reg_file[457]) );
  DFFPOSX1 reg_file_reg_3__74_ ( .D(n24670), .CLK(clk), .Q(reg_file[458]) );
  DFFPOSX1 reg_file_reg_3__75_ ( .D(n24669), .CLK(clk), .Q(reg_file[459]) );
  DFFPOSX1 reg_file_reg_3__76_ ( .D(n24668), .CLK(clk), .Q(reg_file[460]) );
  DFFPOSX1 reg_file_reg_3__77_ ( .D(n24667), .CLK(clk), .Q(reg_file[461]) );
  DFFPOSX1 reg_file_reg_3__78_ ( .D(n24666), .CLK(clk), .Q(reg_file[462]) );
  DFFPOSX1 reg_file_reg_3__79_ ( .D(n24665), .CLK(clk), .Q(reg_file[463]) );
  DFFPOSX1 reg_file_reg_3__80_ ( .D(n24664), .CLK(clk), .Q(reg_file[464]) );
  DFFPOSX1 reg_file_reg_3__81_ ( .D(n24663), .CLK(clk), .Q(reg_file[465]) );
  DFFPOSX1 reg_file_reg_3__82_ ( .D(n24662), .CLK(clk), .Q(reg_file[466]) );
  DFFPOSX1 reg_file_reg_3__83_ ( .D(n24661), .CLK(clk), .Q(reg_file[467]) );
  DFFPOSX1 reg_file_reg_3__84_ ( .D(n24660), .CLK(clk), .Q(reg_file[468]) );
  DFFPOSX1 reg_file_reg_3__85_ ( .D(n24659), .CLK(clk), .Q(reg_file[469]) );
  DFFPOSX1 reg_file_reg_3__86_ ( .D(n24658), .CLK(clk), .Q(reg_file[470]) );
  DFFPOSX1 reg_file_reg_3__87_ ( .D(n24657), .CLK(clk), .Q(reg_file[471]) );
  DFFPOSX1 reg_file_reg_3__88_ ( .D(n24656), .CLK(clk), .Q(reg_file[472]) );
  DFFPOSX1 reg_file_reg_3__89_ ( .D(n24655), .CLK(clk), .Q(reg_file[473]) );
  DFFPOSX1 reg_file_reg_3__90_ ( .D(n24654), .CLK(clk), .Q(reg_file[474]) );
  DFFPOSX1 reg_file_reg_3__91_ ( .D(n24653), .CLK(clk), .Q(reg_file[475]) );
  DFFPOSX1 reg_file_reg_3__92_ ( .D(n24652), .CLK(clk), .Q(reg_file[476]) );
  DFFPOSX1 reg_file_reg_3__93_ ( .D(n24651), .CLK(clk), .Q(reg_file[477]) );
  DFFPOSX1 reg_file_reg_3__94_ ( .D(n24650), .CLK(clk), .Q(reg_file[478]) );
  DFFPOSX1 reg_file_reg_3__95_ ( .D(n24649), .CLK(clk), .Q(reg_file[479]) );
  DFFPOSX1 reg_file_reg_3__96_ ( .D(n24648), .CLK(clk), .Q(reg_file[480]) );
  DFFPOSX1 reg_file_reg_3__97_ ( .D(n24647), .CLK(clk), .Q(reg_file[481]) );
  DFFPOSX1 reg_file_reg_3__98_ ( .D(n24646), .CLK(clk), .Q(reg_file[482]) );
  DFFPOSX1 reg_file_reg_3__99_ ( .D(n24645), .CLK(clk), .Q(reg_file[483]) );
  DFFPOSX1 reg_file_reg_3__100_ ( .D(n24644), .CLK(clk), .Q(reg_file[484]) );
  DFFPOSX1 reg_file_reg_3__101_ ( .D(n24643), .CLK(clk), .Q(reg_file[485]) );
  DFFPOSX1 reg_file_reg_3__102_ ( .D(n24642), .CLK(clk), .Q(reg_file[486]) );
  DFFPOSX1 reg_file_reg_3__103_ ( .D(n24641), .CLK(clk), .Q(reg_file[487]) );
  DFFPOSX1 reg_file_reg_3__104_ ( .D(n24640), .CLK(clk), .Q(reg_file[488]) );
  DFFPOSX1 reg_file_reg_3__105_ ( .D(n24639), .CLK(clk), .Q(reg_file[489]) );
  DFFPOSX1 reg_file_reg_3__106_ ( .D(n24638), .CLK(clk), .Q(reg_file[490]) );
  DFFPOSX1 reg_file_reg_3__107_ ( .D(n24637), .CLK(clk), .Q(reg_file[491]) );
  DFFPOSX1 reg_file_reg_3__108_ ( .D(n24636), .CLK(clk), .Q(reg_file[492]) );
  DFFPOSX1 reg_file_reg_3__109_ ( .D(n24635), .CLK(clk), .Q(reg_file[493]) );
  DFFPOSX1 reg_file_reg_3__110_ ( .D(n24634), .CLK(clk), .Q(reg_file[494]) );
  DFFPOSX1 reg_file_reg_3__111_ ( .D(n24633), .CLK(clk), .Q(reg_file[495]) );
  DFFPOSX1 reg_file_reg_3__112_ ( .D(n24632), .CLK(clk), .Q(reg_file[496]) );
  DFFPOSX1 reg_file_reg_3__113_ ( .D(n24631), .CLK(clk), .Q(reg_file[497]) );
  DFFPOSX1 reg_file_reg_3__114_ ( .D(n24630), .CLK(clk), .Q(reg_file[498]) );
  DFFPOSX1 reg_file_reg_3__115_ ( .D(n24629), .CLK(clk), .Q(reg_file[499]) );
  DFFPOSX1 reg_file_reg_3__116_ ( .D(n24628), .CLK(clk), .Q(reg_file[500]) );
  DFFPOSX1 reg_file_reg_3__117_ ( .D(n24627), .CLK(clk), .Q(reg_file[501]) );
  DFFPOSX1 reg_file_reg_3__118_ ( .D(n24626), .CLK(clk), .Q(reg_file[502]) );
  DFFPOSX1 reg_file_reg_3__119_ ( .D(n24625), .CLK(clk), .Q(reg_file[503]) );
  DFFPOSX1 reg_file_reg_3__120_ ( .D(n24624), .CLK(clk), .Q(reg_file[504]) );
  DFFPOSX1 reg_file_reg_3__121_ ( .D(n24623), .CLK(clk), .Q(reg_file[505]) );
  DFFPOSX1 reg_file_reg_3__122_ ( .D(n24622), .CLK(clk), .Q(reg_file[506]) );
  DFFPOSX1 reg_file_reg_3__123_ ( .D(n24621), .CLK(clk), .Q(reg_file[507]) );
  DFFPOSX1 reg_file_reg_3__124_ ( .D(n24620), .CLK(clk), .Q(reg_file[508]) );
  DFFPOSX1 reg_file_reg_3__125_ ( .D(n24619), .CLK(clk), .Q(reg_file[509]) );
  DFFPOSX1 reg_file_reg_3__126_ ( .D(n24618), .CLK(clk), .Q(reg_file[510]) );
  DFFPOSX1 reg_file_reg_3__127_ ( .D(n24617), .CLK(clk), .Q(reg_file[511]) );
  DFFPOSX1 reg_file_reg_4__0_ ( .D(n24616), .CLK(clk), .Q(reg_file[512]) );
  DFFPOSX1 reg_file_reg_4__1_ ( .D(n24615), .CLK(clk), .Q(reg_file[513]) );
  DFFPOSX1 reg_file_reg_4__2_ ( .D(n24614), .CLK(clk), .Q(reg_file[514]) );
  DFFPOSX1 reg_file_reg_4__3_ ( .D(n24613), .CLK(clk), .Q(reg_file[515]) );
  DFFPOSX1 reg_file_reg_4__4_ ( .D(n24612), .CLK(clk), .Q(reg_file[516]) );
  DFFPOSX1 reg_file_reg_4__5_ ( .D(n24611), .CLK(clk), .Q(reg_file[517]) );
  DFFPOSX1 reg_file_reg_4__6_ ( .D(n24610), .CLK(clk), .Q(reg_file[518]) );
  DFFPOSX1 reg_file_reg_4__7_ ( .D(n24609), .CLK(clk), .Q(reg_file[519]) );
  DFFPOSX1 reg_file_reg_4__8_ ( .D(n24608), .CLK(clk), .Q(reg_file[520]) );
  DFFPOSX1 reg_file_reg_4__9_ ( .D(n24607), .CLK(clk), .Q(reg_file[521]) );
  DFFPOSX1 reg_file_reg_4__10_ ( .D(n24606), .CLK(clk), .Q(reg_file[522]) );
  DFFPOSX1 reg_file_reg_4__11_ ( .D(n24605), .CLK(clk), .Q(reg_file[523]) );
  DFFPOSX1 reg_file_reg_4__12_ ( .D(n24604), .CLK(clk), .Q(reg_file[524]) );
  DFFPOSX1 reg_file_reg_4__13_ ( .D(n24603), .CLK(clk), .Q(reg_file[525]) );
  DFFPOSX1 reg_file_reg_4__14_ ( .D(n24602), .CLK(clk), .Q(reg_file[526]) );
  DFFPOSX1 reg_file_reg_4__15_ ( .D(n24601), .CLK(clk), .Q(reg_file[527]) );
  DFFPOSX1 reg_file_reg_4__16_ ( .D(n24600), .CLK(clk), .Q(reg_file[528]) );
  DFFPOSX1 reg_file_reg_4__17_ ( .D(n24599), .CLK(clk), .Q(reg_file[529]) );
  DFFPOSX1 reg_file_reg_4__18_ ( .D(n24598), .CLK(clk), .Q(reg_file[530]) );
  DFFPOSX1 reg_file_reg_4__19_ ( .D(n24597), .CLK(clk), .Q(reg_file[531]) );
  DFFPOSX1 reg_file_reg_4__20_ ( .D(n24596), .CLK(clk), .Q(reg_file[532]) );
  DFFPOSX1 reg_file_reg_4__21_ ( .D(n24595), .CLK(clk), .Q(reg_file[533]) );
  DFFPOSX1 reg_file_reg_4__22_ ( .D(n24594), .CLK(clk), .Q(reg_file[534]) );
  DFFPOSX1 reg_file_reg_4__23_ ( .D(n24593), .CLK(clk), .Q(reg_file[535]) );
  DFFPOSX1 reg_file_reg_4__24_ ( .D(n24592), .CLK(clk), .Q(reg_file[536]) );
  DFFPOSX1 reg_file_reg_4__25_ ( .D(n24591), .CLK(clk), .Q(reg_file[537]) );
  DFFPOSX1 reg_file_reg_4__26_ ( .D(n24590), .CLK(clk), .Q(reg_file[538]) );
  DFFPOSX1 reg_file_reg_4__27_ ( .D(n24589), .CLK(clk), .Q(reg_file[539]) );
  DFFPOSX1 reg_file_reg_4__28_ ( .D(n24588), .CLK(clk), .Q(reg_file[540]) );
  DFFPOSX1 reg_file_reg_4__29_ ( .D(n24587), .CLK(clk), .Q(reg_file[541]) );
  DFFPOSX1 reg_file_reg_4__30_ ( .D(n24586), .CLK(clk), .Q(reg_file[542]) );
  DFFPOSX1 reg_file_reg_4__31_ ( .D(n24585), .CLK(clk), .Q(reg_file[543]) );
  DFFPOSX1 reg_file_reg_4__32_ ( .D(n24584), .CLK(clk), .Q(reg_file[544]) );
  DFFPOSX1 reg_file_reg_4__33_ ( .D(n24583), .CLK(clk), .Q(reg_file[545]) );
  DFFPOSX1 reg_file_reg_4__34_ ( .D(n24582), .CLK(clk), .Q(reg_file[546]) );
  DFFPOSX1 reg_file_reg_4__35_ ( .D(n24581), .CLK(clk), .Q(reg_file[547]) );
  DFFPOSX1 reg_file_reg_4__36_ ( .D(n24580), .CLK(clk), .Q(reg_file[548]) );
  DFFPOSX1 reg_file_reg_4__37_ ( .D(n24579), .CLK(clk), .Q(reg_file[549]) );
  DFFPOSX1 reg_file_reg_4__38_ ( .D(n24578), .CLK(clk), .Q(reg_file[550]) );
  DFFPOSX1 reg_file_reg_4__39_ ( .D(n24577), .CLK(clk), .Q(reg_file[551]) );
  DFFPOSX1 reg_file_reg_4__40_ ( .D(n24576), .CLK(clk), .Q(reg_file[552]) );
  DFFPOSX1 reg_file_reg_4__41_ ( .D(n24575), .CLK(clk), .Q(reg_file[553]) );
  DFFPOSX1 reg_file_reg_4__42_ ( .D(n24574), .CLK(clk), .Q(reg_file[554]) );
  DFFPOSX1 reg_file_reg_4__43_ ( .D(n24573), .CLK(clk), .Q(reg_file[555]) );
  DFFPOSX1 reg_file_reg_4__44_ ( .D(n24572), .CLK(clk), .Q(reg_file[556]) );
  DFFPOSX1 reg_file_reg_4__45_ ( .D(n24571), .CLK(clk), .Q(reg_file[557]) );
  DFFPOSX1 reg_file_reg_4__46_ ( .D(n24570), .CLK(clk), .Q(reg_file[558]) );
  DFFPOSX1 reg_file_reg_4__47_ ( .D(n24569), .CLK(clk), .Q(reg_file[559]) );
  DFFPOSX1 reg_file_reg_4__48_ ( .D(n24568), .CLK(clk), .Q(reg_file[560]) );
  DFFPOSX1 reg_file_reg_4__49_ ( .D(n24567), .CLK(clk), .Q(reg_file[561]) );
  DFFPOSX1 reg_file_reg_4__50_ ( .D(n24566), .CLK(clk), .Q(reg_file[562]) );
  DFFPOSX1 reg_file_reg_4__51_ ( .D(n24565), .CLK(clk), .Q(reg_file[563]) );
  DFFPOSX1 reg_file_reg_4__52_ ( .D(n24564), .CLK(clk), .Q(reg_file[564]) );
  DFFPOSX1 reg_file_reg_4__53_ ( .D(n24563), .CLK(clk), .Q(reg_file[565]) );
  DFFPOSX1 reg_file_reg_4__54_ ( .D(n24562), .CLK(clk), .Q(reg_file[566]) );
  DFFPOSX1 reg_file_reg_4__55_ ( .D(n24561), .CLK(clk), .Q(reg_file[567]) );
  DFFPOSX1 reg_file_reg_4__56_ ( .D(n24560), .CLK(clk), .Q(reg_file[568]) );
  DFFPOSX1 reg_file_reg_4__57_ ( .D(n24559), .CLK(clk), .Q(reg_file[569]) );
  DFFPOSX1 reg_file_reg_4__58_ ( .D(n24558), .CLK(clk), .Q(reg_file[570]) );
  DFFPOSX1 reg_file_reg_4__59_ ( .D(n24557), .CLK(clk), .Q(reg_file[571]) );
  DFFPOSX1 reg_file_reg_4__60_ ( .D(n24556), .CLK(clk), .Q(reg_file[572]) );
  DFFPOSX1 reg_file_reg_4__61_ ( .D(n24555), .CLK(clk), .Q(reg_file[573]) );
  DFFPOSX1 reg_file_reg_4__62_ ( .D(n24554), .CLK(clk), .Q(reg_file[574]) );
  DFFPOSX1 reg_file_reg_4__63_ ( .D(n24553), .CLK(clk), .Q(reg_file[575]) );
  DFFPOSX1 reg_file_reg_4__64_ ( .D(n24552), .CLK(clk), .Q(reg_file[576]) );
  DFFPOSX1 reg_file_reg_4__65_ ( .D(n24551), .CLK(clk), .Q(reg_file[577]) );
  DFFPOSX1 reg_file_reg_4__66_ ( .D(n24550), .CLK(clk), .Q(reg_file[578]) );
  DFFPOSX1 reg_file_reg_4__67_ ( .D(n24549), .CLK(clk), .Q(reg_file[579]) );
  DFFPOSX1 reg_file_reg_4__68_ ( .D(n24548), .CLK(clk), .Q(reg_file[580]) );
  DFFPOSX1 reg_file_reg_4__69_ ( .D(n24547), .CLK(clk), .Q(reg_file[581]) );
  DFFPOSX1 reg_file_reg_4__70_ ( .D(n24546), .CLK(clk), .Q(reg_file[582]) );
  DFFPOSX1 reg_file_reg_4__71_ ( .D(n24545), .CLK(clk), .Q(reg_file[583]) );
  DFFPOSX1 reg_file_reg_4__72_ ( .D(n24544), .CLK(clk), .Q(reg_file[584]) );
  DFFPOSX1 reg_file_reg_4__73_ ( .D(n24543), .CLK(clk), .Q(reg_file[585]) );
  DFFPOSX1 reg_file_reg_4__74_ ( .D(n24542), .CLK(clk), .Q(reg_file[586]) );
  DFFPOSX1 reg_file_reg_4__75_ ( .D(n24541), .CLK(clk), .Q(reg_file[587]) );
  DFFPOSX1 reg_file_reg_4__76_ ( .D(n24540), .CLK(clk), .Q(reg_file[588]) );
  DFFPOSX1 reg_file_reg_4__77_ ( .D(n24539), .CLK(clk), .Q(reg_file[589]) );
  DFFPOSX1 reg_file_reg_4__78_ ( .D(n24538), .CLK(clk), .Q(reg_file[590]) );
  DFFPOSX1 reg_file_reg_4__79_ ( .D(n24537), .CLK(clk), .Q(reg_file[591]) );
  DFFPOSX1 reg_file_reg_4__80_ ( .D(n24536), .CLK(clk), .Q(reg_file[592]) );
  DFFPOSX1 reg_file_reg_4__81_ ( .D(n24535), .CLK(clk), .Q(reg_file[593]) );
  DFFPOSX1 reg_file_reg_4__82_ ( .D(n24534), .CLK(clk), .Q(reg_file[594]) );
  DFFPOSX1 reg_file_reg_4__83_ ( .D(n24533), .CLK(clk), .Q(reg_file[595]) );
  DFFPOSX1 reg_file_reg_4__84_ ( .D(n24532), .CLK(clk), .Q(reg_file[596]) );
  DFFPOSX1 reg_file_reg_4__85_ ( .D(n24531), .CLK(clk), .Q(reg_file[597]) );
  DFFPOSX1 reg_file_reg_4__86_ ( .D(n24530), .CLK(clk), .Q(reg_file[598]) );
  DFFPOSX1 reg_file_reg_4__87_ ( .D(n24529), .CLK(clk), .Q(reg_file[599]) );
  DFFPOSX1 reg_file_reg_4__88_ ( .D(n24528), .CLK(clk), .Q(reg_file[600]) );
  DFFPOSX1 reg_file_reg_4__89_ ( .D(n24527), .CLK(clk), .Q(reg_file[601]) );
  DFFPOSX1 reg_file_reg_4__90_ ( .D(n24526), .CLK(clk), .Q(reg_file[602]) );
  DFFPOSX1 reg_file_reg_4__91_ ( .D(n24525), .CLK(clk), .Q(reg_file[603]) );
  DFFPOSX1 reg_file_reg_4__92_ ( .D(n24524), .CLK(clk), .Q(reg_file[604]) );
  DFFPOSX1 reg_file_reg_4__93_ ( .D(n24523), .CLK(clk), .Q(reg_file[605]) );
  DFFPOSX1 reg_file_reg_4__94_ ( .D(n24522), .CLK(clk), .Q(reg_file[606]) );
  DFFPOSX1 reg_file_reg_4__95_ ( .D(n24521), .CLK(clk), .Q(reg_file[607]) );
  DFFPOSX1 reg_file_reg_4__96_ ( .D(n24520), .CLK(clk), .Q(reg_file[608]) );
  DFFPOSX1 reg_file_reg_4__97_ ( .D(n24519), .CLK(clk), .Q(reg_file[609]) );
  DFFPOSX1 reg_file_reg_4__98_ ( .D(n24518), .CLK(clk), .Q(reg_file[610]) );
  DFFPOSX1 reg_file_reg_4__99_ ( .D(n24517), .CLK(clk), .Q(reg_file[611]) );
  DFFPOSX1 reg_file_reg_4__100_ ( .D(n24516), .CLK(clk), .Q(reg_file[612]) );
  DFFPOSX1 reg_file_reg_4__101_ ( .D(n24515), .CLK(clk), .Q(reg_file[613]) );
  DFFPOSX1 reg_file_reg_4__102_ ( .D(n24514), .CLK(clk), .Q(reg_file[614]) );
  DFFPOSX1 reg_file_reg_4__103_ ( .D(n24513), .CLK(clk), .Q(reg_file[615]) );
  DFFPOSX1 reg_file_reg_4__104_ ( .D(n24512), .CLK(clk), .Q(reg_file[616]) );
  DFFPOSX1 reg_file_reg_4__105_ ( .D(n24511), .CLK(clk), .Q(reg_file[617]) );
  DFFPOSX1 reg_file_reg_4__106_ ( .D(n24510), .CLK(clk), .Q(reg_file[618]) );
  DFFPOSX1 reg_file_reg_4__107_ ( .D(n24509), .CLK(clk), .Q(reg_file[619]) );
  DFFPOSX1 reg_file_reg_4__108_ ( .D(n24508), .CLK(clk), .Q(reg_file[620]) );
  DFFPOSX1 reg_file_reg_4__109_ ( .D(n24507), .CLK(clk), .Q(reg_file[621]) );
  DFFPOSX1 reg_file_reg_4__110_ ( .D(n24506), .CLK(clk), .Q(reg_file[622]) );
  DFFPOSX1 reg_file_reg_4__111_ ( .D(n24505), .CLK(clk), .Q(reg_file[623]) );
  DFFPOSX1 reg_file_reg_4__112_ ( .D(n24504), .CLK(clk), .Q(reg_file[624]) );
  DFFPOSX1 reg_file_reg_4__113_ ( .D(n24503), .CLK(clk), .Q(reg_file[625]) );
  DFFPOSX1 reg_file_reg_4__114_ ( .D(n24502), .CLK(clk), .Q(reg_file[626]) );
  DFFPOSX1 reg_file_reg_4__115_ ( .D(n24501), .CLK(clk), .Q(reg_file[627]) );
  DFFPOSX1 reg_file_reg_4__116_ ( .D(n24500), .CLK(clk), .Q(reg_file[628]) );
  DFFPOSX1 reg_file_reg_4__117_ ( .D(n24499), .CLK(clk), .Q(reg_file[629]) );
  DFFPOSX1 reg_file_reg_4__118_ ( .D(n24498), .CLK(clk), .Q(reg_file[630]) );
  DFFPOSX1 reg_file_reg_4__119_ ( .D(n24497), .CLK(clk), .Q(reg_file[631]) );
  DFFPOSX1 reg_file_reg_4__120_ ( .D(n24496), .CLK(clk), .Q(reg_file[632]) );
  DFFPOSX1 reg_file_reg_4__121_ ( .D(n24495), .CLK(clk), .Q(reg_file[633]) );
  DFFPOSX1 reg_file_reg_4__122_ ( .D(n24494), .CLK(clk), .Q(reg_file[634]) );
  DFFPOSX1 reg_file_reg_4__123_ ( .D(n24493), .CLK(clk), .Q(reg_file[635]) );
  DFFPOSX1 reg_file_reg_4__124_ ( .D(n24492), .CLK(clk), .Q(reg_file[636]) );
  DFFPOSX1 reg_file_reg_4__125_ ( .D(n24491), .CLK(clk), .Q(reg_file[637]) );
  DFFPOSX1 reg_file_reg_4__126_ ( .D(n24490), .CLK(clk), .Q(reg_file[638]) );
  DFFPOSX1 reg_file_reg_4__127_ ( .D(n24489), .CLK(clk), .Q(reg_file[639]) );
  DFFPOSX1 reg_file_reg_5__0_ ( .D(n24488), .CLK(clk), .Q(reg_file[640]) );
  DFFPOSX1 reg_file_reg_5__1_ ( .D(n24487), .CLK(clk), .Q(reg_file[641]) );
  DFFPOSX1 reg_file_reg_5__2_ ( .D(n24486), .CLK(clk), .Q(reg_file[642]) );
  DFFPOSX1 reg_file_reg_5__3_ ( .D(n24485), .CLK(clk), .Q(reg_file[643]) );
  DFFPOSX1 reg_file_reg_5__4_ ( .D(n24484), .CLK(clk), .Q(reg_file[644]) );
  DFFPOSX1 reg_file_reg_5__5_ ( .D(n24483), .CLK(clk), .Q(reg_file[645]) );
  DFFPOSX1 reg_file_reg_5__6_ ( .D(n24482), .CLK(clk), .Q(reg_file[646]) );
  DFFPOSX1 reg_file_reg_5__7_ ( .D(n24481), .CLK(clk), .Q(reg_file[647]) );
  DFFPOSX1 reg_file_reg_5__8_ ( .D(n24480), .CLK(clk), .Q(reg_file[648]) );
  DFFPOSX1 reg_file_reg_5__9_ ( .D(n24479), .CLK(clk), .Q(reg_file[649]) );
  DFFPOSX1 reg_file_reg_5__10_ ( .D(n24478), .CLK(clk), .Q(reg_file[650]) );
  DFFPOSX1 reg_file_reg_5__11_ ( .D(n24477), .CLK(clk), .Q(reg_file[651]) );
  DFFPOSX1 reg_file_reg_5__12_ ( .D(n24476), .CLK(clk), .Q(reg_file[652]) );
  DFFPOSX1 reg_file_reg_5__13_ ( .D(n24475), .CLK(clk), .Q(reg_file[653]) );
  DFFPOSX1 reg_file_reg_5__14_ ( .D(n24474), .CLK(clk), .Q(reg_file[654]) );
  DFFPOSX1 reg_file_reg_5__15_ ( .D(n24473), .CLK(clk), .Q(reg_file[655]) );
  DFFPOSX1 reg_file_reg_5__16_ ( .D(n24472), .CLK(clk), .Q(reg_file[656]) );
  DFFPOSX1 reg_file_reg_5__17_ ( .D(n24471), .CLK(clk), .Q(reg_file[657]) );
  DFFPOSX1 reg_file_reg_5__18_ ( .D(n24470), .CLK(clk), .Q(reg_file[658]) );
  DFFPOSX1 reg_file_reg_5__19_ ( .D(n24469), .CLK(clk), .Q(reg_file[659]) );
  DFFPOSX1 reg_file_reg_5__20_ ( .D(n24468), .CLK(clk), .Q(reg_file[660]) );
  DFFPOSX1 reg_file_reg_5__21_ ( .D(n24467), .CLK(clk), .Q(reg_file[661]) );
  DFFPOSX1 reg_file_reg_5__22_ ( .D(n24466), .CLK(clk), .Q(reg_file[662]) );
  DFFPOSX1 reg_file_reg_5__23_ ( .D(n24465), .CLK(clk), .Q(reg_file[663]) );
  DFFPOSX1 reg_file_reg_5__24_ ( .D(n24464), .CLK(clk), .Q(reg_file[664]) );
  DFFPOSX1 reg_file_reg_5__25_ ( .D(n24463), .CLK(clk), .Q(reg_file[665]) );
  DFFPOSX1 reg_file_reg_5__26_ ( .D(n24462), .CLK(clk), .Q(reg_file[666]) );
  DFFPOSX1 reg_file_reg_5__27_ ( .D(n24461), .CLK(clk), .Q(reg_file[667]) );
  DFFPOSX1 reg_file_reg_5__28_ ( .D(n24460), .CLK(clk), .Q(reg_file[668]) );
  DFFPOSX1 reg_file_reg_5__29_ ( .D(n24459), .CLK(clk), .Q(reg_file[669]) );
  DFFPOSX1 reg_file_reg_5__30_ ( .D(n24458), .CLK(clk), .Q(reg_file[670]) );
  DFFPOSX1 reg_file_reg_5__31_ ( .D(n24457), .CLK(clk), .Q(reg_file[671]) );
  DFFPOSX1 reg_file_reg_5__32_ ( .D(n24456), .CLK(clk), .Q(reg_file[672]) );
  DFFPOSX1 reg_file_reg_5__33_ ( .D(n24455), .CLK(clk), .Q(reg_file[673]) );
  DFFPOSX1 reg_file_reg_5__34_ ( .D(n24454), .CLK(clk), .Q(reg_file[674]) );
  DFFPOSX1 reg_file_reg_5__35_ ( .D(n24453), .CLK(clk), .Q(reg_file[675]) );
  DFFPOSX1 reg_file_reg_5__36_ ( .D(n24452), .CLK(clk), .Q(reg_file[676]) );
  DFFPOSX1 reg_file_reg_5__37_ ( .D(n24451), .CLK(clk), .Q(reg_file[677]) );
  DFFPOSX1 reg_file_reg_5__38_ ( .D(n24450), .CLK(clk), .Q(reg_file[678]) );
  DFFPOSX1 reg_file_reg_5__39_ ( .D(n24449), .CLK(clk), .Q(reg_file[679]) );
  DFFPOSX1 reg_file_reg_5__40_ ( .D(n24448), .CLK(clk), .Q(reg_file[680]) );
  DFFPOSX1 reg_file_reg_5__41_ ( .D(n24447), .CLK(clk), .Q(reg_file[681]) );
  DFFPOSX1 reg_file_reg_5__42_ ( .D(n24446), .CLK(clk), .Q(reg_file[682]) );
  DFFPOSX1 reg_file_reg_5__43_ ( .D(n24445), .CLK(clk), .Q(reg_file[683]) );
  DFFPOSX1 reg_file_reg_5__44_ ( .D(n24444), .CLK(clk), .Q(reg_file[684]) );
  DFFPOSX1 reg_file_reg_5__45_ ( .D(n24443), .CLK(clk), .Q(reg_file[685]) );
  DFFPOSX1 reg_file_reg_5__46_ ( .D(n24442), .CLK(clk), .Q(reg_file[686]) );
  DFFPOSX1 reg_file_reg_5__47_ ( .D(n24441), .CLK(clk), .Q(reg_file[687]) );
  DFFPOSX1 reg_file_reg_5__48_ ( .D(n24440), .CLK(clk), .Q(reg_file[688]) );
  DFFPOSX1 reg_file_reg_5__49_ ( .D(n24439), .CLK(clk), .Q(reg_file[689]) );
  DFFPOSX1 reg_file_reg_5__50_ ( .D(n24438), .CLK(clk), .Q(reg_file[690]) );
  DFFPOSX1 reg_file_reg_5__51_ ( .D(n24437), .CLK(clk), .Q(reg_file[691]) );
  DFFPOSX1 reg_file_reg_5__52_ ( .D(n24436), .CLK(clk), .Q(reg_file[692]) );
  DFFPOSX1 reg_file_reg_5__53_ ( .D(n24435), .CLK(clk), .Q(reg_file[693]) );
  DFFPOSX1 reg_file_reg_5__54_ ( .D(n24434), .CLK(clk), .Q(reg_file[694]) );
  DFFPOSX1 reg_file_reg_5__55_ ( .D(n24433), .CLK(clk), .Q(reg_file[695]) );
  DFFPOSX1 reg_file_reg_5__56_ ( .D(n24432), .CLK(clk), .Q(reg_file[696]) );
  DFFPOSX1 reg_file_reg_5__57_ ( .D(n24431), .CLK(clk), .Q(reg_file[697]) );
  DFFPOSX1 reg_file_reg_5__58_ ( .D(n24430), .CLK(clk), .Q(reg_file[698]) );
  DFFPOSX1 reg_file_reg_5__59_ ( .D(n24429), .CLK(clk), .Q(reg_file[699]) );
  DFFPOSX1 reg_file_reg_5__60_ ( .D(n24428), .CLK(clk), .Q(reg_file[700]) );
  DFFPOSX1 reg_file_reg_5__61_ ( .D(n24427), .CLK(clk), .Q(reg_file[701]) );
  DFFPOSX1 reg_file_reg_5__62_ ( .D(n24426), .CLK(clk), .Q(reg_file[702]) );
  DFFPOSX1 reg_file_reg_5__63_ ( .D(n24425), .CLK(clk), .Q(reg_file[703]) );
  DFFPOSX1 reg_file_reg_5__64_ ( .D(n24424), .CLK(clk), .Q(reg_file[704]) );
  DFFPOSX1 reg_file_reg_5__65_ ( .D(n24423), .CLK(clk), .Q(reg_file[705]) );
  DFFPOSX1 reg_file_reg_5__66_ ( .D(n24422), .CLK(clk), .Q(reg_file[706]) );
  DFFPOSX1 reg_file_reg_5__67_ ( .D(n24421), .CLK(clk), .Q(reg_file[707]) );
  DFFPOSX1 reg_file_reg_5__68_ ( .D(n24420), .CLK(clk), .Q(reg_file[708]) );
  DFFPOSX1 reg_file_reg_5__69_ ( .D(n24419), .CLK(clk), .Q(reg_file[709]) );
  DFFPOSX1 reg_file_reg_5__70_ ( .D(n24418), .CLK(clk), .Q(reg_file[710]) );
  DFFPOSX1 reg_file_reg_5__71_ ( .D(n24417), .CLK(clk), .Q(reg_file[711]) );
  DFFPOSX1 reg_file_reg_5__72_ ( .D(n24416), .CLK(clk), .Q(reg_file[712]) );
  DFFPOSX1 reg_file_reg_5__73_ ( .D(n24415), .CLK(clk), .Q(reg_file[713]) );
  DFFPOSX1 reg_file_reg_5__74_ ( .D(n24414), .CLK(clk), .Q(reg_file[714]) );
  DFFPOSX1 reg_file_reg_5__75_ ( .D(n24413), .CLK(clk), .Q(reg_file[715]) );
  DFFPOSX1 reg_file_reg_5__76_ ( .D(n24412), .CLK(clk), .Q(reg_file[716]) );
  DFFPOSX1 reg_file_reg_5__77_ ( .D(n24411), .CLK(clk), .Q(reg_file[717]) );
  DFFPOSX1 reg_file_reg_5__78_ ( .D(n24410), .CLK(clk), .Q(reg_file[718]) );
  DFFPOSX1 reg_file_reg_5__79_ ( .D(n24409), .CLK(clk), .Q(reg_file[719]) );
  DFFPOSX1 reg_file_reg_5__80_ ( .D(n24408), .CLK(clk), .Q(reg_file[720]) );
  DFFPOSX1 reg_file_reg_5__81_ ( .D(n24407), .CLK(clk), .Q(reg_file[721]) );
  DFFPOSX1 reg_file_reg_5__82_ ( .D(n24406), .CLK(clk), .Q(reg_file[722]) );
  DFFPOSX1 reg_file_reg_5__83_ ( .D(n24405), .CLK(clk), .Q(reg_file[723]) );
  DFFPOSX1 reg_file_reg_5__84_ ( .D(n24404), .CLK(clk), .Q(reg_file[724]) );
  DFFPOSX1 reg_file_reg_5__85_ ( .D(n24403), .CLK(clk), .Q(reg_file[725]) );
  DFFPOSX1 reg_file_reg_5__86_ ( .D(n24402), .CLK(clk), .Q(reg_file[726]) );
  DFFPOSX1 reg_file_reg_5__87_ ( .D(n24401), .CLK(clk), .Q(reg_file[727]) );
  DFFPOSX1 reg_file_reg_5__88_ ( .D(n24400), .CLK(clk), .Q(reg_file[728]) );
  DFFPOSX1 reg_file_reg_5__89_ ( .D(n24399), .CLK(clk), .Q(reg_file[729]) );
  DFFPOSX1 reg_file_reg_5__90_ ( .D(n24398), .CLK(clk), .Q(reg_file[730]) );
  DFFPOSX1 reg_file_reg_5__91_ ( .D(n24397), .CLK(clk), .Q(reg_file[731]) );
  DFFPOSX1 reg_file_reg_5__92_ ( .D(n24396), .CLK(clk), .Q(reg_file[732]) );
  DFFPOSX1 reg_file_reg_5__93_ ( .D(n24395), .CLK(clk), .Q(reg_file[733]) );
  DFFPOSX1 reg_file_reg_5__94_ ( .D(n24394), .CLK(clk), .Q(reg_file[734]) );
  DFFPOSX1 reg_file_reg_5__95_ ( .D(n24393), .CLK(clk), .Q(reg_file[735]) );
  DFFPOSX1 reg_file_reg_5__96_ ( .D(n24392), .CLK(clk), .Q(reg_file[736]) );
  DFFPOSX1 reg_file_reg_5__97_ ( .D(n24391), .CLK(clk), .Q(reg_file[737]) );
  DFFPOSX1 reg_file_reg_5__98_ ( .D(n24390), .CLK(clk), .Q(reg_file[738]) );
  DFFPOSX1 reg_file_reg_5__99_ ( .D(n24389), .CLK(clk), .Q(reg_file[739]) );
  DFFPOSX1 reg_file_reg_5__100_ ( .D(n24388), .CLK(clk), .Q(reg_file[740]) );
  DFFPOSX1 reg_file_reg_5__101_ ( .D(n24387), .CLK(clk), .Q(reg_file[741]) );
  DFFPOSX1 reg_file_reg_5__102_ ( .D(n24386), .CLK(clk), .Q(reg_file[742]) );
  DFFPOSX1 reg_file_reg_5__103_ ( .D(n24385), .CLK(clk), .Q(reg_file[743]) );
  DFFPOSX1 reg_file_reg_5__104_ ( .D(n24384), .CLK(clk), .Q(reg_file[744]) );
  DFFPOSX1 reg_file_reg_5__105_ ( .D(n24383), .CLK(clk), .Q(reg_file[745]) );
  DFFPOSX1 reg_file_reg_5__106_ ( .D(n24382), .CLK(clk), .Q(reg_file[746]) );
  DFFPOSX1 reg_file_reg_5__107_ ( .D(n24381), .CLK(clk), .Q(reg_file[747]) );
  DFFPOSX1 reg_file_reg_5__108_ ( .D(n24380), .CLK(clk), .Q(reg_file[748]) );
  DFFPOSX1 reg_file_reg_5__109_ ( .D(n24379), .CLK(clk), .Q(reg_file[749]) );
  DFFPOSX1 reg_file_reg_5__110_ ( .D(n24378), .CLK(clk), .Q(reg_file[750]) );
  DFFPOSX1 reg_file_reg_5__111_ ( .D(n24377), .CLK(clk), .Q(reg_file[751]) );
  DFFPOSX1 reg_file_reg_5__112_ ( .D(n24376), .CLK(clk), .Q(reg_file[752]) );
  DFFPOSX1 reg_file_reg_5__113_ ( .D(n24375), .CLK(clk), .Q(reg_file[753]) );
  DFFPOSX1 reg_file_reg_5__114_ ( .D(n24374), .CLK(clk), .Q(reg_file[754]) );
  DFFPOSX1 reg_file_reg_5__115_ ( .D(n24373), .CLK(clk), .Q(reg_file[755]) );
  DFFPOSX1 reg_file_reg_5__116_ ( .D(n24372), .CLK(clk), .Q(reg_file[756]) );
  DFFPOSX1 reg_file_reg_5__117_ ( .D(n24371), .CLK(clk), .Q(reg_file[757]) );
  DFFPOSX1 reg_file_reg_5__118_ ( .D(n24370), .CLK(clk), .Q(reg_file[758]) );
  DFFPOSX1 reg_file_reg_5__119_ ( .D(n24369), .CLK(clk), .Q(reg_file[759]) );
  DFFPOSX1 reg_file_reg_5__120_ ( .D(n24368), .CLK(clk), .Q(reg_file[760]) );
  DFFPOSX1 reg_file_reg_5__121_ ( .D(n24367), .CLK(clk), .Q(reg_file[761]) );
  DFFPOSX1 reg_file_reg_5__122_ ( .D(n24366), .CLK(clk), .Q(reg_file[762]) );
  DFFPOSX1 reg_file_reg_5__123_ ( .D(n24365), .CLK(clk), .Q(reg_file[763]) );
  DFFPOSX1 reg_file_reg_5__124_ ( .D(n24364), .CLK(clk), .Q(reg_file[764]) );
  DFFPOSX1 reg_file_reg_5__125_ ( .D(n24363), .CLK(clk), .Q(reg_file[765]) );
  DFFPOSX1 reg_file_reg_5__126_ ( .D(n24362), .CLK(clk), .Q(reg_file[766]) );
  DFFPOSX1 reg_file_reg_5__127_ ( .D(n24361), .CLK(clk), .Q(reg_file[767]) );
  DFFPOSX1 reg_file_reg_6__0_ ( .D(n24360), .CLK(clk), .Q(reg_file[768]) );
  DFFPOSX1 reg_file_reg_6__1_ ( .D(n24359), .CLK(clk), .Q(reg_file[769]) );
  DFFPOSX1 reg_file_reg_6__2_ ( .D(n24358), .CLK(clk), .Q(reg_file[770]) );
  DFFPOSX1 reg_file_reg_6__3_ ( .D(n24357), .CLK(clk), .Q(reg_file[771]) );
  DFFPOSX1 reg_file_reg_6__4_ ( .D(n24356), .CLK(clk), .Q(reg_file[772]) );
  DFFPOSX1 reg_file_reg_6__5_ ( .D(n24355), .CLK(clk), .Q(reg_file[773]) );
  DFFPOSX1 reg_file_reg_6__6_ ( .D(n24354), .CLK(clk), .Q(reg_file[774]) );
  DFFPOSX1 reg_file_reg_6__7_ ( .D(n24353), .CLK(clk), .Q(reg_file[775]) );
  DFFPOSX1 reg_file_reg_6__8_ ( .D(n24352), .CLK(clk), .Q(reg_file[776]) );
  DFFPOSX1 reg_file_reg_6__9_ ( .D(n24351), .CLK(clk), .Q(reg_file[777]) );
  DFFPOSX1 reg_file_reg_6__10_ ( .D(n24350), .CLK(clk), .Q(reg_file[778]) );
  DFFPOSX1 reg_file_reg_6__11_ ( .D(n24349), .CLK(clk), .Q(reg_file[779]) );
  DFFPOSX1 reg_file_reg_6__12_ ( .D(n24348), .CLK(clk), .Q(reg_file[780]) );
  DFFPOSX1 reg_file_reg_6__13_ ( .D(n24347), .CLK(clk), .Q(reg_file[781]) );
  DFFPOSX1 reg_file_reg_6__14_ ( .D(n24346), .CLK(clk), .Q(reg_file[782]) );
  DFFPOSX1 reg_file_reg_6__15_ ( .D(n24345), .CLK(clk), .Q(reg_file[783]) );
  DFFPOSX1 reg_file_reg_6__16_ ( .D(n24344), .CLK(clk), .Q(reg_file[784]) );
  DFFPOSX1 reg_file_reg_6__17_ ( .D(n24343), .CLK(clk), .Q(reg_file[785]) );
  DFFPOSX1 reg_file_reg_6__18_ ( .D(n24342), .CLK(clk), .Q(reg_file[786]) );
  DFFPOSX1 reg_file_reg_6__19_ ( .D(n24341), .CLK(clk), .Q(reg_file[787]) );
  DFFPOSX1 reg_file_reg_6__20_ ( .D(n24340), .CLK(clk), .Q(reg_file[788]) );
  DFFPOSX1 reg_file_reg_6__21_ ( .D(n24339), .CLK(clk), .Q(reg_file[789]) );
  DFFPOSX1 reg_file_reg_6__22_ ( .D(n24338), .CLK(clk), .Q(reg_file[790]) );
  DFFPOSX1 reg_file_reg_6__23_ ( .D(n24337), .CLK(clk), .Q(reg_file[791]) );
  DFFPOSX1 reg_file_reg_6__24_ ( .D(n24336), .CLK(clk), .Q(reg_file[792]) );
  DFFPOSX1 reg_file_reg_6__25_ ( .D(n24335), .CLK(clk), .Q(reg_file[793]) );
  DFFPOSX1 reg_file_reg_6__26_ ( .D(n24334), .CLK(clk), .Q(reg_file[794]) );
  DFFPOSX1 reg_file_reg_6__27_ ( .D(n24333), .CLK(clk), .Q(reg_file[795]) );
  DFFPOSX1 reg_file_reg_6__28_ ( .D(n24332), .CLK(clk), .Q(reg_file[796]) );
  DFFPOSX1 reg_file_reg_6__29_ ( .D(n24331), .CLK(clk), .Q(reg_file[797]) );
  DFFPOSX1 reg_file_reg_6__30_ ( .D(n24330), .CLK(clk), .Q(reg_file[798]) );
  DFFPOSX1 reg_file_reg_6__31_ ( .D(n24329), .CLK(clk), .Q(reg_file[799]) );
  DFFPOSX1 reg_file_reg_6__32_ ( .D(n24328), .CLK(clk), .Q(reg_file[800]) );
  DFFPOSX1 reg_file_reg_6__33_ ( .D(n24327), .CLK(clk), .Q(reg_file[801]) );
  DFFPOSX1 reg_file_reg_6__34_ ( .D(n24326), .CLK(clk), .Q(reg_file[802]) );
  DFFPOSX1 reg_file_reg_6__35_ ( .D(n24325), .CLK(clk), .Q(reg_file[803]) );
  DFFPOSX1 reg_file_reg_6__36_ ( .D(n24324), .CLK(clk), .Q(reg_file[804]) );
  DFFPOSX1 reg_file_reg_6__37_ ( .D(n24323), .CLK(clk), .Q(reg_file[805]) );
  DFFPOSX1 reg_file_reg_6__38_ ( .D(n24322), .CLK(clk), .Q(reg_file[806]) );
  DFFPOSX1 reg_file_reg_6__39_ ( .D(n24321), .CLK(clk), .Q(reg_file[807]) );
  DFFPOSX1 reg_file_reg_6__40_ ( .D(n24320), .CLK(clk), .Q(reg_file[808]) );
  DFFPOSX1 reg_file_reg_6__41_ ( .D(n24319), .CLK(clk), .Q(reg_file[809]) );
  DFFPOSX1 reg_file_reg_6__42_ ( .D(n24318), .CLK(clk), .Q(reg_file[810]) );
  DFFPOSX1 reg_file_reg_6__43_ ( .D(n24317), .CLK(clk), .Q(reg_file[811]) );
  DFFPOSX1 reg_file_reg_6__44_ ( .D(n24316), .CLK(clk), .Q(reg_file[812]) );
  DFFPOSX1 reg_file_reg_6__45_ ( .D(n24315), .CLK(clk), .Q(reg_file[813]) );
  DFFPOSX1 reg_file_reg_6__46_ ( .D(n24314), .CLK(clk), .Q(reg_file[814]) );
  DFFPOSX1 reg_file_reg_6__47_ ( .D(n24313), .CLK(clk), .Q(reg_file[815]) );
  DFFPOSX1 reg_file_reg_6__48_ ( .D(n24312), .CLK(clk), .Q(reg_file[816]) );
  DFFPOSX1 reg_file_reg_6__49_ ( .D(n24311), .CLK(clk), .Q(reg_file[817]) );
  DFFPOSX1 reg_file_reg_6__50_ ( .D(n24310), .CLK(clk), .Q(reg_file[818]) );
  DFFPOSX1 reg_file_reg_6__51_ ( .D(n24309), .CLK(clk), .Q(reg_file[819]) );
  DFFPOSX1 reg_file_reg_6__52_ ( .D(n24308), .CLK(clk), .Q(reg_file[820]) );
  DFFPOSX1 reg_file_reg_6__53_ ( .D(n24307), .CLK(clk), .Q(reg_file[821]) );
  DFFPOSX1 reg_file_reg_6__54_ ( .D(n24306), .CLK(clk), .Q(reg_file[822]) );
  DFFPOSX1 reg_file_reg_6__55_ ( .D(n24305), .CLK(clk), .Q(reg_file[823]) );
  DFFPOSX1 reg_file_reg_6__56_ ( .D(n24304), .CLK(clk), .Q(reg_file[824]) );
  DFFPOSX1 reg_file_reg_6__57_ ( .D(n24303), .CLK(clk), .Q(reg_file[825]) );
  DFFPOSX1 reg_file_reg_6__58_ ( .D(n24302), .CLK(clk), .Q(reg_file[826]) );
  DFFPOSX1 reg_file_reg_6__59_ ( .D(n24301), .CLK(clk), .Q(reg_file[827]) );
  DFFPOSX1 reg_file_reg_6__60_ ( .D(n24300), .CLK(clk), .Q(reg_file[828]) );
  DFFPOSX1 reg_file_reg_6__61_ ( .D(n24299), .CLK(clk), .Q(reg_file[829]) );
  DFFPOSX1 reg_file_reg_6__62_ ( .D(n24298), .CLK(clk), .Q(reg_file[830]) );
  DFFPOSX1 reg_file_reg_6__63_ ( .D(n24297), .CLK(clk), .Q(reg_file[831]) );
  DFFPOSX1 reg_file_reg_6__64_ ( .D(n24296), .CLK(clk), .Q(reg_file[832]) );
  DFFPOSX1 reg_file_reg_6__65_ ( .D(n24295), .CLK(clk), .Q(reg_file[833]) );
  DFFPOSX1 reg_file_reg_6__66_ ( .D(n24294), .CLK(clk), .Q(reg_file[834]) );
  DFFPOSX1 reg_file_reg_6__67_ ( .D(n24293), .CLK(clk), .Q(reg_file[835]) );
  DFFPOSX1 reg_file_reg_6__68_ ( .D(n24292), .CLK(clk), .Q(reg_file[836]) );
  DFFPOSX1 reg_file_reg_6__69_ ( .D(n24291), .CLK(clk), .Q(reg_file[837]) );
  DFFPOSX1 reg_file_reg_6__70_ ( .D(n24290), .CLK(clk), .Q(reg_file[838]) );
  DFFPOSX1 reg_file_reg_6__71_ ( .D(n24289), .CLK(clk), .Q(reg_file[839]) );
  DFFPOSX1 reg_file_reg_6__72_ ( .D(n24288), .CLK(clk), .Q(reg_file[840]) );
  DFFPOSX1 reg_file_reg_6__73_ ( .D(n24287), .CLK(clk), .Q(reg_file[841]) );
  DFFPOSX1 reg_file_reg_6__74_ ( .D(n24286), .CLK(clk), .Q(reg_file[842]) );
  DFFPOSX1 reg_file_reg_6__75_ ( .D(n24285), .CLK(clk), .Q(reg_file[843]) );
  DFFPOSX1 reg_file_reg_6__76_ ( .D(n24284), .CLK(clk), .Q(reg_file[844]) );
  DFFPOSX1 reg_file_reg_6__77_ ( .D(n24283), .CLK(clk), .Q(reg_file[845]) );
  DFFPOSX1 reg_file_reg_6__78_ ( .D(n24282), .CLK(clk), .Q(reg_file[846]) );
  DFFPOSX1 reg_file_reg_6__79_ ( .D(n24281), .CLK(clk), .Q(reg_file[847]) );
  DFFPOSX1 reg_file_reg_6__80_ ( .D(n24280), .CLK(clk), .Q(reg_file[848]) );
  DFFPOSX1 reg_file_reg_6__81_ ( .D(n24279), .CLK(clk), .Q(reg_file[849]) );
  DFFPOSX1 reg_file_reg_6__82_ ( .D(n24278), .CLK(clk), .Q(reg_file[850]) );
  DFFPOSX1 reg_file_reg_6__83_ ( .D(n24277), .CLK(clk), .Q(reg_file[851]) );
  DFFPOSX1 reg_file_reg_6__84_ ( .D(n24276), .CLK(clk), .Q(reg_file[852]) );
  DFFPOSX1 reg_file_reg_6__85_ ( .D(n24275), .CLK(clk), .Q(reg_file[853]) );
  DFFPOSX1 reg_file_reg_6__86_ ( .D(n24274), .CLK(clk), .Q(reg_file[854]) );
  DFFPOSX1 reg_file_reg_6__87_ ( .D(n24273), .CLK(clk), .Q(reg_file[855]) );
  DFFPOSX1 reg_file_reg_6__88_ ( .D(n24272), .CLK(clk), .Q(reg_file[856]) );
  DFFPOSX1 reg_file_reg_6__89_ ( .D(n24271), .CLK(clk), .Q(reg_file[857]) );
  DFFPOSX1 reg_file_reg_6__90_ ( .D(n24270), .CLK(clk), .Q(reg_file[858]) );
  DFFPOSX1 reg_file_reg_6__91_ ( .D(n24269), .CLK(clk), .Q(reg_file[859]) );
  DFFPOSX1 reg_file_reg_6__92_ ( .D(n24268), .CLK(clk), .Q(reg_file[860]) );
  DFFPOSX1 reg_file_reg_6__93_ ( .D(n24267), .CLK(clk), .Q(reg_file[861]) );
  DFFPOSX1 reg_file_reg_6__94_ ( .D(n24266), .CLK(clk), .Q(reg_file[862]) );
  DFFPOSX1 reg_file_reg_6__95_ ( .D(n24265), .CLK(clk), .Q(reg_file[863]) );
  DFFPOSX1 reg_file_reg_6__96_ ( .D(n24264), .CLK(clk), .Q(reg_file[864]) );
  DFFPOSX1 reg_file_reg_6__97_ ( .D(n24263), .CLK(clk), .Q(reg_file[865]) );
  DFFPOSX1 reg_file_reg_6__98_ ( .D(n24262), .CLK(clk), .Q(reg_file[866]) );
  DFFPOSX1 reg_file_reg_6__99_ ( .D(n24261), .CLK(clk), .Q(reg_file[867]) );
  DFFPOSX1 reg_file_reg_6__100_ ( .D(n24260), .CLK(clk), .Q(reg_file[868]) );
  DFFPOSX1 reg_file_reg_6__101_ ( .D(n24259), .CLK(clk), .Q(reg_file[869]) );
  DFFPOSX1 reg_file_reg_6__102_ ( .D(n24258), .CLK(clk), .Q(reg_file[870]) );
  DFFPOSX1 reg_file_reg_6__103_ ( .D(n24257), .CLK(clk), .Q(reg_file[871]) );
  DFFPOSX1 reg_file_reg_6__104_ ( .D(n24256), .CLK(clk), .Q(reg_file[872]) );
  DFFPOSX1 reg_file_reg_6__105_ ( .D(n24255), .CLK(clk), .Q(reg_file[873]) );
  DFFPOSX1 reg_file_reg_6__106_ ( .D(n24254), .CLK(clk), .Q(reg_file[874]) );
  DFFPOSX1 reg_file_reg_6__107_ ( .D(n24253), .CLK(clk), .Q(reg_file[875]) );
  DFFPOSX1 reg_file_reg_6__108_ ( .D(n24252), .CLK(clk), .Q(reg_file[876]) );
  DFFPOSX1 reg_file_reg_6__109_ ( .D(n24251), .CLK(clk), .Q(reg_file[877]) );
  DFFPOSX1 reg_file_reg_6__110_ ( .D(n24250), .CLK(clk), .Q(reg_file[878]) );
  DFFPOSX1 reg_file_reg_6__111_ ( .D(n24249), .CLK(clk), .Q(reg_file[879]) );
  DFFPOSX1 reg_file_reg_6__112_ ( .D(n24248), .CLK(clk), .Q(reg_file[880]) );
  DFFPOSX1 reg_file_reg_6__113_ ( .D(n24247), .CLK(clk), .Q(reg_file[881]) );
  DFFPOSX1 reg_file_reg_6__114_ ( .D(n24246), .CLK(clk), .Q(reg_file[882]) );
  DFFPOSX1 reg_file_reg_6__115_ ( .D(n24245), .CLK(clk), .Q(reg_file[883]) );
  DFFPOSX1 reg_file_reg_6__116_ ( .D(n24244), .CLK(clk), .Q(reg_file[884]) );
  DFFPOSX1 reg_file_reg_6__117_ ( .D(n24243), .CLK(clk), .Q(reg_file[885]) );
  DFFPOSX1 reg_file_reg_6__118_ ( .D(n24242), .CLK(clk), .Q(reg_file[886]) );
  DFFPOSX1 reg_file_reg_6__119_ ( .D(n24241), .CLK(clk), .Q(reg_file[887]) );
  DFFPOSX1 reg_file_reg_6__120_ ( .D(n24240), .CLK(clk), .Q(reg_file[888]) );
  DFFPOSX1 reg_file_reg_6__121_ ( .D(n24239), .CLK(clk), .Q(reg_file[889]) );
  DFFPOSX1 reg_file_reg_6__122_ ( .D(n24238), .CLK(clk), .Q(reg_file[890]) );
  DFFPOSX1 reg_file_reg_6__123_ ( .D(n24237), .CLK(clk), .Q(reg_file[891]) );
  DFFPOSX1 reg_file_reg_6__124_ ( .D(n24236), .CLK(clk), .Q(reg_file[892]) );
  DFFPOSX1 reg_file_reg_6__125_ ( .D(n24235), .CLK(clk), .Q(reg_file[893]) );
  DFFPOSX1 reg_file_reg_6__126_ ( .D(n24234), .CLK(clk), .Q(reg_file[894]) );
  DFFPOSX1 reg_file_reg_6__127_ ( .D(n24233), .CLK(clk), .Q(reg_file[895]) );
  DFFPOSX1 reg_file_reg_7__0_ ( .D(n24232), .CLK(clk), .Q(reg_file[896]) );
  DFFPOSX1 reg_file_reg_7__1_ ( .D(n24231), .CLK(clk), .Q(reg_file[897]) );
  DFFPOSX1 reg_file_reg_7__2_ ( .D(n24230), .CLK(clk), .Q(reg_file[898]) );
  DFFPOSX1 reg_file_reg_7__3_ ( .D(n24229), .CLK(clk), .Q(reg_file[899]) );
  DFFPOSX1 reg_file_reg_7__4_ ( .D(n24228), .CLK(clk), .Q(reg_file[900]) );
  DFFPOSX1 reg_file_reg_7__5_ ( .D(n24227), .CLK(clk), .Q(reg_file[901]) );
  DFFPOSX1 reg_file_reg_7__6_ ( .D(n24226), .CLK(clk), .Q(reg_file[902]) );
  DFFPOSX1 reg_file_reg_7__7_ ( .D(n24225), .CLK(clk), .Q(reg_file[903]) );
  DFFPOSX1 reg_file_reg_7__8_ ( .D(n24224), .CLK(clk), .Q(reg_file[904]) );
  DFFPOSX1 reg_file_reg_7__9_ ( .D(n24223), .CLK(clk), .Q(reg_file[905]) );
  DFFPOSX1 reg_file_reg_7__10_ ( .D(n24222), .CLK(clk), .Q(reg_file[906]) );
  DFFPOSX1 reg_file_reg_7__11_ ( .D(n24221), .CLK(clk), .Q(reg_file[907]) );
  DFFPOSX1 reg_file_reg_7__12_ ( .D(n24220), .CLK(clk), .Q(reg_file[908]) );
  DFFPOSX1 reg_file_reg_7__13_ ( .D(n24219), .CLK(clk), .Q(reg_file[909]) );
  DFFPOSX1 reg_file_reg_7__14_ ( .D(n24218), .CLK(clk), .Q(reg_file[910]) );
  DFFPOSX1 reg_file_reg_7__15_ ( .D(n24217), .CLK(clk), .Q(reg_file[911]) );
  DFFPOSX1 reg_file_reg_7__16_ ( .D(n24216), .CLK(clk), .Q(reg_file[912]) );
  DFFPOSX1 reg_file_reg_7__17_ ( .D(n24215), .CLK(clk), .Q(reg_file[913]) );
  DFFPOSX1 reg_file_reg_7__18_ ( .D(n24214), .CLK(clk), .Q(reg_file[914]) );
  DFFPOSX1 reg_file_reg_7__19_ ( .D(n24213), .CLK(clk), .Q(reg_file[915]) );
  DFFPOSX1 reg_file_reg_7__20_ ( .D(n24212), .CLK(clk), .Q(reg_file[916]) );
  DFFPOSX1 reg_file_reg_7__21_ ( .D(n24211), .CLK(clk), .Q(reg_file[917]) );
  DFFPOSX1 reg_file_reg_7__22_ ( .D(n24210), .CLK(clk), .Q(reg_file[918]) );
  DFFPOSX1 reg_file_reg_7__23_ ( .D(n24209), .CLK(clk), .Q(reg_file[919]) );
  DFFPOSX1 reg_file_reg_7__24_ ( .D(n24208), .CLK(clk), .Q(reg_file[920]) );
  DFFPOSX1 reg_file_reg_7__25_ ( .D(n24207), .CLK(clk), .Q(reg_file[921]) );
  DFFPOSX1 reg_file_reg_7__26_ ( .D(n24206), .CLK(clk), .Q(reg_file[922]) );
  DFFPOSX1 reg_file_reg_7__27_ ( .D(n24205), .CLK(clk), .Q(reg_file[923]) );
  DFFPOSX1 reg_file_reg_7__28_ ( .D(n24204), .CLK(clk), .Q(reg_file[924]) );
  DFFPOSX1 reg_file_reg_7__29_ ( .D(n24203), .CLK(clk), .Q(reg_file[925]) );
  DFFPOSX1 reg_file_reg_7__30_ ( .D(n24202), .CLK(clk), .Q(reg_file[926]) );
  DFFPOSX1 reg_file_reg_7__31_ ( .D(n24201), .CLK(clk), .Q(reg_file[927]) );
  DFFPOSX1 reg_file_reg_7__32_ ( .D(n24200), .CLK(clk), .Q(reg_file[928]) );
  DFFPOSX1 reg_file_reg_7__33_ ( .D(n24199), .CLK(clk), .Q(reg_file[929]) );
  DFFPOSX1 reg_file_reg_7__34_ ( .D(n24198), .CLK(clk), .Q(reg_file[930]) );
  DFFPOSX1 reg_file_reg_7__35_ ( .D(n24197), .CLK(clk), .Q(reg_file[931]) );
  DFFPOSX1 reg_file_reg_7__36_ ( .D(n24196), .CLK(clk), .Q(reg_file[932]) );
  DFFPOSX1 reg_file_reg_7__37_ ( .D(n24195), .CLK(clk), .Q(reg_file[933]) );
  DFFPOSX1 reg_file_reg_7__38_ ( .D(n24194), .CLK(clk), .Q(reg_file[934]) );
  DFFPOSX1 reg_file_reg_7__39_ ( .D(n24193), .CLK(clk), .Q(reg_file[935]) );
  DFFPOSX1 reg_file_reg_7__40_ ( .D(n24192), .CLK(clk), .Q(reg_file[936]) );
  DFFPOSX1 reg_file_reg_7__41_ ( .D(n24191), .CLK(clk), .Q(reg_file[937]) );
  DFFPOSX1 reg_file_reg_7__42_ ( .D(n24190), .CLK(clk), .Q(reg_file[938]) );
  DFFPOSX1 reg_file_reg_7__43_ ( .D(n24189), .CLK(clk), .Q(reg_file[939]) );
  DFFPOSX1 reg_file_reg_7__44_ ( .D(n24188), .CLK(clk), .Q(reg_file[940]) );
  DFFPOSX1 reg_file_reg_7__45_ ( .D(n24187), .CLK(clk), .Q(reg_file[941]) );
  DFFPOSX1 reg_file_reg_7__46_ ( .D(n24186), .CLK(clk), .Q(reg_file[942]) );
  DFFPOSX1 reg_file_reg_7__47_ ( .D(n24185), .CLK(clk), .Q(reg_file[943]) );
  DFFPOSX1 reg_file_reg_7__48_ ( .D(n24184), .CLK(clk), .Q(reg_file[944]) );
  DFFPOSX1 reg_file_reg_7__49_ ( .D(n24183), .CLK(clk), .Q(reg_file[945]) );
  DFFPOSX1 reg_file_reg_7__50_ ( .D(n24182), .CLK(clk), .Q(reg_file[946]) );
  DFFPOSX1 reg_file_reg_7__51_ ( .D(n24181), .CLK(clk), .Q(reg_file[947]) );
  DFFPOSX1 reg_file_reg_7__52_ ( .D(n24180), .CLK(clk), .Q(reg_file[948]) );
  DFFPOSX1 reg_file_reg_7__53_ ( .D(n24179), .CLK(clk), .Q(reg_file[949]) );
  DFFPOSX1 reg_file_reg_7__54_ ( .D(n24178), .CLK(clk), .Q(reg_file[950]) );
  DFFPOSX1 reg_file_reg_7__55_ ( .D(n24177), .CLK(clk), .Q(reg_file[951]) );
  DFFPOSX1 reg_file_reg_7__56_ ( .D(n24176), .CLK(clk), .Q(reg_file[952]) );
  DFFPOSX1 reg_file_reg_7__57_ ( .D(n24175), .CLK(clk), .Q(reg_file[953]) );
  DFFPOSX1 reg_file_reg_7__58_ ( .D(n24174), .CLK(clk), .Q(reg_file[954]) );
  DFFPOSX1 reg_file_reg_7__59_ ( .D(n24173), .CLK(clk), .Q(reg_file[955]) );
  DFFPOSX1 reg_file_reg_7__60_ ( .D(n24172), .CLK(clk), .Q(reg_file[956]) );
  DFFPOSX1 reg_file_reg_7__61_ ( .D(n24171), .CLK(clk), .Q(reg_file[957]) );
  DFFPOSX1 reg_file_reg_7__62_ ( .D(n24170), .CLK(clk), .Q(reg_file[958]) );
  DFFPOSX1 reg_file_reg_7__63_ ( .D(n24169), .CLK(clk), .Q(reg_file[959]) );
  DFFPOSX1 reg_file_reg_7__64_ ( .D(n24168), .CLK(clk), .Q(reg_file[960]) );
  DFFPOSX1 reg_file_reg_7__65_ ( .D(n24167), .CLK(clk), .Q(reg_file[961]) );
  DFFPOSX1 reg_file_reg_7__66_ ( .D(n24166), .CLK(clk), .Q(reg_file[962]) );
  DFFPOSX1 reg_file_reg_7__67_ ( .D(n24165), .CLK(clk), .Q(reg_file[963]) );
  DFFPOSX1 reg_file_reg_7__68_ ( .D(n24164), .CLK(clk), .Q(reg_file[964]) );
  DFFPOSX1 reg_file_reg_7__69_ ( .D(n24163), .CLK(clk), .Q(reg_file[965]) );
  DFFPOSX1 reg_file_reg_7__70_ ( .D(n24162), .CLK(clk), .Q(reg_file[966]) );
  DFFPOSX1 reg_file_reg_7__71_ ( .D(n24161), .CLK(clk), .Q(reg_file[967]) );
  DFFPOSX1 reg_file_reg_7__72_ ( .D(n24160), .CLK(clk), .Q(reg_file[968]) );
  DFFPOSX1 reg_file_reg_7__73_ ( .D(n24159), .CLK(clk), .Q(reg_file[969]) );
  DFFPOSX1 reg_file_reg_7__74_ ( .D(n24158), .CLK(clk), .Q(reg_file[970]) );
  DFFPOSX1 reg_file_reg_7__75_ ( .D(n24157), .CLK(clk), .Q(reg_file[971]) );
  DFFPOSX1 reg_file_reg_7__76_ ( .D(n24156), .CLK(clk), .Q(reg_file[972]) );
  DFFPOSX1 reg_file_reg_7__77_ ( .D(n24155), .CLK(clk), .Q(reg_file[973]) );
  DFFPOSX1 reg_file_reg_7__78_ ( .D(n24154), .CLK(clk), .Q(reg_file[974]) );
  DFFPOSX1 reg_file_reg_7__79_ ( .D(n24153), .CLK(clk), .Q(reg_file[975]) );
  DFFPOSX1 reg_file_reg_7__80_ ( .D(n24152), .CLK(clk), .Q(reg_file[976]) );
  DFFPOSX1 reg_file_reg_7__81_ ( .D(n24151), .CLK(clk), .Q(reg_file[977]) );
  DFFPOSX1 reg_file_reg_7__82_ ( .D(n24150), .CLK(clk), .Q(reg_file[978]) );
  DFFPOSX1 reg_file_reg_7__83_ ( .D(n24149), .CLK(clk), .Q(reg_file[979]) );
  DFFPOSX1 reg_file_reg_7__84_ ( .D(n24148), .CLK(clk), .Q(reg_file[980]) );
  DFFPOSX1 reg_file_reg_7__85_ ( .D(n24147), .CLK(clk), .Q(reg_file[981]) );
  DFFPOSX1 reg_file_reg_7__86_ ( .D(n24146), .CLK(clk), .Q(reg_file[982]) );
  DFFPOSX1 reg_file_reg_7__87_ ( .D(n24145), .CLK(clk), .Q(reg_file[983]) );
  DFFPOSX1 reg_file_reg_7__88_ ( .D(n24144), .CLK(clk), .Q(reg_file[984]) );
  DFFPOSX1 reg_file_reg_7__89_ ( .D(n24143), .CLK(clk), .Q(reg_file[985]) );
  DFFPOSX1 reg_file_reg_7__90_ ( .D(n24142), .CLK(clk), .Q(reg_file[986]) );
  DFFPOSX1 reg_file_reg_7__91_ ( .D(n24141), .CLK(clk), .Q(reg_file[987]) );
  DFFPOSX1 reg_file_reg_7__92_ ( .D(n24140), .CLK(clk), .Q(reg_file[988]) );
  DFFPOSX1 reg_file_reg_7__93_ ( .D(n24139), .CLK(clk), .Q(reg_file[989]) );
  DFFPOSX1 reg_file_reg_7__94_ ( .D(n24138), .CLK(clk), .Q(reg_file[990]) );
  DFFPOSX1 reg_file_reg_7__95_ ( .D(n24137), .CLK(clk), .Q(reg_file[991]) );
  DFFPOSX1 reg_file_reg_7__96_ ( .D(n24136), .CLK(clk), .Q(reg_file[992]) );
  DFFPOSX1 reg_file_reg_7__97_ ( .D(n24135), .CLK(clk), .Q(reg_file[993]) );
  DFFPOSX1 reg_file_reg_7__98_ ( .D(n24134), .CLK(clk), .Q(reg_file[994]) );
  DFFPOSX1 reg_file_reg_7__99_ ( .D(n24133), .CLK(clk), .Q(reg_file[995]) );
  DFFPOSX1 reg_file_reg_7__100_ ( .D(n24132), .CLK(clk), .Q(reg_file[996]) );
  DFFPOSX1 reg_file_reg_7__101_ ( .D(n24131), .CLK(clk), .Q(reg_file[997]) );
  DFFPOSX1 reg_file_reg_7__102_ ( .D(n24130), .CLK(clk), .Q(reg_file[998]) );
  DFFPOSX1 reg_file_reg_7__103_ ( .D(n24129), .CLK(clk), .Q(reg_file[999]) );
  DFFPOSX1 reg_file_reg_7__104_ ( .D(n24128), .CLK(clk), .Q(reg_file[1000]) );
  DFFPOSX1 reg_file_reg_7__105_ ( .D(n24127), .CLK(clk), .Q(reg_file[1001]) );
  DFFPOSX1 reg_file_reg_7__106_ ( .D(n24126), .CLK(clk), .Q(reg_file[1002]) );
  DFFPOSX1 reg_file_reg_7__107_ ( .D(n24125), .CLK(clk), .Q(reg_file[1003]) );
  DFFPOSX1 reg_file_reg_7__108_ ( .D(n24124), .CLK(clk), .Q(reg_file[1004]) );
  DFFPOSX1 reg_file_reg_7__109_ ( .D(n24123), .CLK(clk), .Q(reg_file[1005]) );
  DFFPOSX1 reg_file_reg_7__110_ ( .D(n24122), .CLK(clk), .Q(reg_file[1006]) );
  DFFPOSX1 reg_file_reg_7__111_ ( .D(n24121), .CLK(clk), .Q(reg_file[1007]) );
  DFFPOSX1 reg_file_reg_7__112_ ( .D(n24120), .CLK(clk), .Q(reg_file[1008]) );
  DFFPOSX1 reg_file_reg_7__113_ ( .D(n24119), .CLK(clk), .Q(reg_file[1009]) );
  DFFPOSX1 reg_file_reg_7__114_ ( .D(n24118), .CLK(clk), .Q(reg_file[1010]) );
  DFFPOSX1 reg_file_reg_7__115_ ( .D(n24117), .CLK(clk), .Q(reg_file[1011]) );
  DFFPOSX1 reg_file_reg_7__116_ ( .D(n24116), .CLK(clk), .Q(reg_file[1012]) );
  DFFPOSX1 reg_file_reg_7__117_ ( .D(n24115), .CLK(clk), .Q(reg_file[1013]) );
  DFFPOSX1 reg_file_reg_7__118_ ( .D(n24114), .CLK(clk), .Q(reg_file[1014]) );
  DFFPOSX1 reg_file_reg_7__119_ ( .D(n24113), .CLK(clk), .Q(reg_file[1015]) );
  DFFPOSX1 reg_file_reg_7__120_ ( .D(n24112), .CLK(clk), .Q(reg_file[1016]) );
  DFFPOSX1 reg_file_reg_7__121_ ( .D(n24111), .CLK(clk), .Q(reg_file[1017]) );
  DFFPOSX1 reg_file_reg_7__122_ ( .D(n24110), .CLK(clk), .Q(reg_file[1018]) );
  DFFPOSX1 reg_file_reg_7__123_ ( .D(n24109), .CLK(clk), .Q(reg_file[1019]) );
  DFFPOSX1 reg_file_reg_7__124_ ( .D(n24108), .CLK(clk), .Q(reg_file[1020]) );
  DFFPOSX1 reg_file_reg_7__125_ ( .D(n24107), .CLK(clk), .Q(reg_file[1021]) );
  DFFPOSX1 reg_file_reg_7__126_ ( .D(n24106), .CLK(clk), .Q(reg_file[1022]) );
  DFFPOSX1 reg_file_reg_7__127_ ( .D(n24105), .CLK(clk), .Q(reg_file[1023]) );
  DFFPOSX1 reg_file_reg_8__0_ ( .D(n24104), .CLK(clk), .Q(reg_file[1024]) );
  DFFPOSX1 reg_file_reg_8__1_ ( .D(n24103), .CLK(clk), .Q(reg_file[1025]) );
  DFFPOSX1 reg_file_reg_8__2_ ( .D(n24102), .CLK(clk), .Q(reg_file[1026]) );
  DFFPOSX1 reg_file_reg_8__3_ ( .D(n24101), .CLK(clk), .Q(reg_file[1027]) );
  DFFPOSX1 reg_file_reg_8__4_ ( .D(n24100), .CLK(clk), .Q(reg_file[1028]) );
  DFFPOSX1 reg_file_reg_8__5_ ( .D(n24099), .CLK(clk), .Q(reg_file[1029]) );
  DFFPOSX1 reg_file_reg_8__6_ ( .D(n24098), .CLK(clk), .Q(reg_file[1030]) );
  DFFPOSX1 reg_file_reg_8__7_ ( .D(n24097), .CLK(clk), .Q(reg_file[1031]) );
  DFFPOSX1 reg_file_reg_8__8_ ( .D(n24096), .CLK(clk), .Q(reg_file[1032]) );
  DFFPOSX1 reg_file_reg_8__9_ ( .D(n24095), .CLK(clk), .Q(reg_file[1033]) );
  DFFPOSX1 reg_file_reg_8__10_ ( .D(n24094), .CLK(clk), .Q(reg_file[1034]) );
  DFFPOSX1 reg_file_reg_8__11_ ( .D(n24093), .CLK(clk), .Q(reg_file[1035]) );
  DFFPOSX1 reg_file_reg_8__12_ ( .D(n24092), .CLK(clk), .Q(reg_file[1036]) );
  DFFPOSX1 reg_file_reg_8__13_ ( .D(n24091), .CLK(clk), .Q(reg_file[1037]) );
  DFFPOSX1 reg_file_reg_8__14_ ( .D(n24090), .CLK(clk), .Q(reg_file[1038]) );
  DFFPOSX1 reg_file_reg_8__15_ ( .D(n24089), .CLK(clk), .Q(reg_file[1039]) );
  DFFPOSX1 reg_file_reg_8__16_ ( .D(n24088), .CLK(clk), .Q(reg_file[1040]) );
  DFFPOSX1 reg_file_reg_8__17_ ( .D(n24087), .CLK(clk), .Q(reg_file[1041]) );
  DFFPOSX1 reg_file_reg_8__18_ ( .D(n24086), .CLK(clk), .Q(reg_file[1042]) );
  DFFPOSX1 reg_file_reg_8__19_ ( .D(n24085), .CLK(clk), .Q(reg_file[1043]) );
  DFFPOSX1 reg_file_reg_8__20_ ( .D(n24084), .CLK(clk), .Q(reg_file[1044]) );
  DFFPOSX1 reg_file_reg_8__21_ ( .D(n24083), .CLK(clk), .Q(reg_file[1045]) );
  DFFPOSX1 reg_file_reg_8__22_ ( .D(n24082), .CLK(clk), .Q(reg_file[1046]) );
  DFFPOSX1 reg_file_reg_8__23_ ( .D(n24081), .CLK(clk), .Q(reg_file[1047]) );
  DFFPOSX1 reg_file_reg_8__24_ ( .D(n24080), .CLK(clk), .Q(reg_file[1048]) );
  DFFPOSX1 reg_file_reg_8__25_ ( .D(n24079), .CLK(clk), .Q(reg_file[1049]) );
  DFFPOSX1 reg_file_reg_8__26_ ( .D(n24078), .CLK(clk), .Q(reg_file[1050]) );
  DFFPOSX1 reg_file_reg_8__27_ ( .D(n24077), .CLK(clk), .Q(reg_file[1051]) );
  DFFPOSX1 reg_file_reg_8__28_ ( .D(n24076), .CLK(clk), .Q(reg_file[1052]) );
  DFFPOSX1 reg_file_reg_8__29_ ( .D(n24075), .CLK(clk), .Q(reg_file[1053]) );
  DFFPOSX1 reg_file_reg_8__30_ ( .D(n24074), .CLK(clk), .Q(reg_file[1054]) );
  DFFPOSX1 reg_file_reg_8__31_ ( .D(n24073), .CLK(clk), .Q(reg_file[1055]) );
  DFFPOSX1 reg_file_reg_8__32_ ( .D(n24072), .CLK(clk), .Q(reg_file[1056]) );
  DFFPOSX1 reg_file_reg_8__33_ ( .D(n24071), .CLK(clk), .Q(reg_file[1057]) );
  DFFPOSX1 reg_file_reg_8__34_ ( .D(n24070), .CLK(clk), .Q(reg_file[1058]) );
  DFFPOSX1 reg_file_reg_8__35_ ( .D(n24069), .CLK(clk), .Q(reg_file[1059]) );
  DFFPOSX1 reg_file_reg_8__36_ ( .D(n24068), .CLK(clk), .Q(reg_file[1060]) );
  DFFPOSX1 reg_file_reg_8__37_ ( .D(n24067), .CLK(clk), .Q(reg_file[1061]) );
  DFFPOSX1 reg_file_reg_8__38_ ( .D(n24066), .CLK(clk), .Q(reg_file[1062]) );
  DFFPOSX1 reg_file_reg_8__39_ ( .D(n24065), .CLK(clk), .Q(reg_file[1063]) );
  DFFPOSX1 reg_file_reg_8__40_ ( .D(n24064), .CLK(clk), .Q(reg_file[1064]) );
  DFFPOSX1 reg_file_reg_8__41_ ( .D(n24063), .CLK(clk), .Q(reg_file[1065]) );
  DFFPOSX1 reg_file_reg_8__42_ ( .D(n24062), .CLK(clk), .Q(reg_file[1066]) );
  DFFPOSX1 reg_file_reg_8__43_ ( .D(n24061), .CLK(clk), .Q(reg_file[1067]) );
  DFFPOSX1 reg_file_reg_8__44_ ( .D(n24060), .CLK(clk), .Q(reg_file[1068]) );
  DFFPOSX1 reg_file_reg_8__45_ ( .D(n24059), .CLK(clk), .Q(reg_file[1069]) );
  DFFPOSX1 reg_file_reg_8__46_ ( .D(n24058), .CLK(clk), .Q(reg_file[1070]) );
  DFFPOSX1 reg_file_reg_8__47_ ( .D(n24057), .CLK(clk), .Q(reg_file[1071]) );
  DFFPOSX1 reg_file_reg_8__48_ ( .D(n24056), .CLK(clk), .Q(reg_file[1072]) );
  DFFPOSX1 reg_file_reg_8__49_ ( .D(n24055), .CLK(clk), .Q(reg_file[1073]) );
  DFFPOSX1 reg_file_reg_8__50_ ( .D(n24054), .CLK(clk), .Q(reg_file[1074]) );
  DFFPOSX1 reg_file_reg_8__51_ ( .D(n24053), .CLK(clk), .Q(reg_file[1075]) );
  DFFPOSX1 reg_file_reg_8__52_ ( .D(n24052), .CLK(clk), .Q(reg_file[1076]) );
  DFFPOSX1 reg_file_reg_8__53_ ( .D(n24051), .CLK(clk), .Q(reg_file[1077]) );
  DFFPOSX1 reg_file_reg_8__54_ ( .D(n24050), .CLK(clk), .Q(reg_file[1078]) );
  DFFPOSX1 reg_file_reg_8__55_ ( .D(n24049), .CLK(clk), .Q(reg_file[1079]) );
  DFFPOSX1 reg_file_reg_8__56_ ( .D(n24048), .CLK(clk), .Q(reg_file[1080]) );
  DFFPOSX1 reg_file_reg_8__57_ ( .D(n24047), .CLK(clk), .Q(reg_file[1081]) );
  DFFPOSX1 reg_file_reg_8__58_ ( .D(n24046), .CLK(clk), .Q(reg_file[1082]) );
  DFFPOSX1 reg_file_reg_8__59_ ( .D(n24045), .CLK(clk), .Q(reg_file[1083]) );
  DFFPOSX1 reg_file_reg_8__60_ ( .D(n24044), .CLK(clk), .Q(reg_file[1084]) );
  DFFPOSX1 reg_file_reg_8__61_ ( .D(n24043), .CLK(clk), .Q(reg_file[1085]) );
  DFFPOSX1 reg_file_reg_8__62_ ( .D(n24042), .CLK(clk), .Q(reg_file[1086]) );
  DFFPOSX1 reg_file_reg_8__63_ ( .D(n24041), .CLK(clk), .Q(reg_file[1087]) );
  DFFPOSX1 reg_file_reg_8__64_ ( .D(n24040), .CLK(clk), .Q(reg_file[1088]) );
  DFFPOSX1 reg_file_reg_8__65_ ( .D(n24039), .CLK(clk), .Q(reg_file[1089]) );
  DFFPOSX1 reg_file_reg_8__66_ ( .D(n24038), .CLK(clk), .Q(reg_file[1090]) );
  DFFPOSX1 reg_file_reg_8__67_ ( .D(n24037), .CLK(clk), .Q(reg_file[1091]) );
  DFFPOSX1 reg_file_reg_8__68_ ( .D(n24036), .CLK(clk), .Q(reg_file[1092]) );
  DFFPOSX1 reg_file_reg_8__69_ ( .D(n24035), .CLK(clk), .Q(reg_file[1093]) );
  DFFPOSX1 reg_file_reg_8__70_ ( .D(n24034), .CLK(clk), .Q(reg_file[1094]) );
  DFFPOSX1 reg_file_reg_8__71_ ( .D(n24033), .CLK(clk), .Q(reg_file[1095]) );
  DFFPOSX1 reg_file_reg_8__72_ ( .D(n24032), .CLK(clk), .Q(reg_file[1096]) );
  DFFPOSX1 reg_file_reg_8__73_ ( .D(n24031), .CLK(clk), .Q(reg_file[1097]) );
  DFFPOSX1 reg_file_reg_8__74_ ( .D(n24030), .CLK(clk), .Q(reg_file[1098]) );
  DFFPOSX1 reg_file_reg_8__75_ ( .D(n24029), .CLK(clk), .Q(reg_file[1099]) );
  DFFPOSX1 reg_file_reg_8__76_ ( .D(n24028), .CLK(clk), .Q(reg_file[1100]) );
  DFFPOSX1 reg_file_reg_8__77_ ( .D(n24027), .CLK(clk), .Q(reg_file[1101]) );
  DFFPOSX1 reg_file_reg_8__78_ ( .D(n24026), .CLK(clk), .Q(reg_file[1102]) );
  DFFPOSX1 reg_file_reg_8__79_ ( .D(n24025), .CLK(clk), .Q(reg_file[1103]) );
  DFFPOSX1 reg_file_reg_8__80_ ( .D(n24024), .CLK(clk), .Q(reg_file[1104]) );
  DFFPOSX1 reg_file_reg_8__81_ ( .D(n24023), .CLK(clk), .Q(reg_file[1105]) );
  DFFPOSX1 reg_file_reg_8__82_ ( .D(n24022), .CLK(clk), .Q(reg_file[1106]) );
  DFFPOSX1 reg_file_reg_8__83_ ( .D(n24021), .CLK(clk), .Q(reg_file[1107]) );
  DFFPOSX1 reg_file_reg_8__84_ ( .D(n24020), .CLK(clk), .Q(reg_file[1108]) );
  DFFPOSX1 reg_file_reg_8__85_ ( .D(n24019), .CLK(clk), .Q(reg_file[1109]) );
  DFFPOSX1 reg_file_reg_8__86_ ( .D(n24018), .CLK(clk), .Q(reg_file[1110]) );
  DFFPOSX1 reg_file_reg_8__87_ ( .D(n24017), .CLK(clk), .Q(reg_file[1111]) );
  DFFPOSX1 reg_file_reg_8__88_ ( .D(n24016), .CLK(clk), .Q(reg_file[1112]) );
  DFFPOSX1 reg_file_reg_8__89_ ( .D(n24015), .CLK(clk), .Q(reg_file[1113]) );
  DFFPOSX1 reg_file_reg_8__90_ ( .D(n24014), .CLK(clk), .Q(reg_file[1114]) );
  DFFPOSX1 reg_file_reg_8__91_ ( .D(n24013), .CLK(clk), .Q(reg_file[1115]) );
  DFFPOSX1 reg_file_reg_8__92_ ( .D(n24012), .CLK(clk), .Q(reg_file[1116]) );
  DFFPOSX1 reg_file_reg_8__93_ ( .D(n24011), .CLK(clk), .Q(reg_file[1117]) );
  DFFPOSX1 reg_file_reg_8__94_ ( .D(n24010), .CLK(clk), .Q(reg_file[1118]) );
  DFFPOSX1 reg_file_reg_8__95_ ( .D(n24009), .CLK(clk), .Q(reg_file[1119]) );
  DFFPOSX1 reg_file_reg_8__96_ ( .D(n24008), .CLK(clk), .Q(reg_file[1120]) );
  DFFPOSX1 reg_file_reg_8__97_ ( .D(n24007), .CLK(clk), .Q(reg_file[1121]) );
  DFFPOSX1 reg_file_reg_8__98_ ( .D(n24006), .CLK(clk), .Q(reg_file[1122]) );
  DFFPOSX1 reg_file_reg_8__99_ ( .D(n24005), .CLK(clk), .Q(reg_file[1123]) );
  DFFPOSX1 reg_file_reg_8__100_ ( .D(n24004), .CLK(clk), .Q(reg_file[1124]) );
  DFFPOSX1 reg_file_reg_8__101_ ( .D(n24003), .CLK(clk), .Q(reg_file[1125]) );
  DFFPOSX1 reg_file_reg_8__102_ ( .D(n24002), .CLK(clk), .Q(reg_file[1126]) );
  DFFPOSX1 reg_file_reg_8__103_ ( .D(n24001), .CLK(clk), .Q(reg_file[1127]) );
  DFFPOSX1 reg_file_reg_8__104_ ( .D(n24000), .CLK(clk), .Q(reg_file[1128]) );
  DFFPOSX1 reg_file_reg_8__105_ ( .D(n23999), .CLK(clk), .Q(reg_file[1129]) );
  DFFPOSX1 reg_file_reg_8__106_ ( .D(n23998), .CLK(clk), .Q(reg_file[1130]) );
  DFFPOSX1 reg_file_reg_8__107_ ( .D(n23997), .CLK(clk), .Q(reg_file[1131]) );
  DFFPOSX1 reg_file_reg_8__108_ ( .D(n23996), .CLK(clk), .Q(reg_file[1132]) );
  DFFPOSX1 reg_file_reg_8__109_ ( .D(n23995), .CLK(clk), .Q(reg_file[1133]) );
  DFFPOSX1 reg_file_reg_8__110_ ( .D(n23994), .CLK(clk), .Q(reg_file[1134]) );
  DFFPOSX1 reg_file_reg_8__111_ ( .D(n23993), .CLK(clk), .Q(reg_file[1135]) );
  DFFPOSX1 reg_file_reg_8__112_ ( .D(n23992), .CLK(clk), .Q(reg_file[1136]) );
  DFFPOSX1 reg_file_reg_8__113_ ( .D(n23991), .CLK(clk), .Q(reg_file[1137]) );
  DFFPOSX1 reg_file_reg_8__114_ ( .D(n23990), .CLK(clk), .Q(reg_file[1138]) );
  DFFPOSX1 reg_file_reg_8__115_ ( .D(n23989), .CLK(clk), .Q(reg_file[1139]) );
  DFFPOSX1 reg_file_reg_8__116_ ( .D(n23988), .CLK(clk), .Q(reg_file[1140]) );
  DFFPOSX1 reg_file_reg_8__117_ ( .D(n23987), .CLK(clk), .Q(reg_file[1141]) );
  DFFPOSX1 reg_file_reg_8__118_ ( .D(n23986), .CLK(clk), .Q(reg_file[1142]) );
  DFFPOSX1 reg_file_reg_8__119_ ( .D(n23985), .CLK(clk), .Q(reg_file[1143]) );
  DFFPOSX1 reg_file_reg_8__120_ ( .D(n23984), .CLK(clk), .Q(reg_file[1144]) );
  DFFPOSX1 reg_file_reg_8__121_ ( .D(n23983), .CLK(clk), .Q(reg_file[1145]) );
  DFFPOSX1 reg_file_reg_8__122_ ( .D(n23982), .CLK(clk), .Q(reg_file[1146]) );
  DFFPOSX1 reg_file_reg_8__123_ ( .D(n23981), .CLK(clk), .Q(reg_file[1147]) );
  DFFPOSX1 reg_file_reg_8__124_ ( .D(n23980), .CLK(clk), .Q(reg_file[1148]) );
  DFFPOSX1 reg_file_reg_8__125_ ( .D(n23979), .CLK(clk), .Q(reg_file[1149]) );
  DFFPOSX1 reg_file_reg_8__126_ ( .D(n23978), .CLK(clk), .Q(reg_file[1150]) );
  DFFPOSX1 reg_file_reg_8__127_ ( .D(n23977), .CLK(clk), .Q(reg_file[1151]) );
  DFFPOSX1 reg_file_reg_9__0_ ( .D(n23976), .CLK(clk), .Q(reg_file[1152]) );
  DFFPOSX1 reg_file_reg_9__1_ ( .D(n23975), .CLK(clk), .Q(reg_file[1153]) );
  DFFPOSX1 reg_file_reg_9__2_ ( .D(n23974), .CLK(clk), .Q(reg_file[1154]) );
  DFFPOSX1 reg_file_reg_9__3_ ( .D(n23973), .CLK(clk), .Q(reg_file[1155]) );
  DFFPOSX1 reg_file_reg_9__4_ ( .D(n23972), .CLK(clk), .Q(reg_file[1156]) );
  DFFPOSX1 reg_file_reg_9__5_ ( .D(n23971), .CLK(clk), .Q(reg_file[1157]) );
  DFFPOSX1 reg_file_reg_9__6_ ( .D(n23970), .CLK(clk), .Q(reg_file[1158]) );
  DFFPOSX1 reg_file_reg_9__7_ ( .D(n23969), .CLK(clk), .Q(reg_file[1159]) );
  DFFPOSX1 reg_file_reg_9__8_ ( .D(n23968), .CLK(clk), .Q(reg_file[1160]) );
  DFFPOSX1 reg_file_reg_9__9_ ( .D(n23967), .CLK(clk), .Q(reg_file[1161]) );
  DFFPOSX1 reg_file_reg_9__10_ ( .D(n23966), .CLK(clk), .Q(reg_file[1162]) );
  DFFPOSX1 reg_file_reg_9__11_ ( .D(n23965), .CLK(clk), .Q(reg_file[1163]) );
  DFFPOSX1 reg_file_reg_9__12_ ( .D(n23964), .CLK(clk), .Q(reg_file[1164]) );
  DFFPOSX1 reg_file_reg_9__13_ ( .D(n23963), .CLK(clk), .Q(reg_file[1165]) );
  DFFPOSX1 reg_file_reg_9__14_ ( .D(n23962), .CLK(clk), .Q(reg_file[1166]) );
  DFFPOSX1 reg_file_reg_9__15_ ( .D(n23961), .CLK(clk), .Q(reg_file[1167]) );
  DFFPOSX1 reg_file_reg_9__16_ ( .D(n23960), .CLK(clk), .Q(reg_file[1168]) );
  DFFPOSX1 reg_file_reg_9__17_ ( .D(n23959), .CLK(clk), .Q(reg_file[1169]) );
  DFFPOSX1 reg_file_reg_9__18_ ( .D(n23958), .CLK(clk), .Q(reg_file[1170]) );
  DFFPOSX1 reg_file_reg_9__19_ ( .D(n23957), .CLK(clk), .Q(reg_file[1171]) );
  DFFPOSX1 reg_file_reg_9__20_ ( .D(n23956), .CLK(clk), .Q(reg_file[1172]) );
  DFFPOSX1 reg_file_reg_9__21_ ( .D(n23955), .CLK(clk), .Q(reg_file[1173]) );
  DFFPOSX1 reg_file_reg_9__22_ ( .D(n23954), .CLK(clk), .Q(reg_file[1174]) );
  DFFPOSX1 reg_file_reg_9__23_ ( .D(n23953), .CLK(clk), .Q(reg_file[1175]) );
  DFFPOSX1 reg_file_reg_9__24_ ( .D(n23952), .CLK(clk), .Q(reg_file[1176]) );
  DFFPOSX1 reg_file_reg_9__25_ ( .D(n23951), .CLK(clk), .Q(reg_file[1177]) );
  DFFPOSX1 reg_file_reg_9__26_ ( .D(n23950), .CLK(clk), .Q(reg_file[1178]) );
  DFFPOSX1 reg_file_reg_9__27_ ( .D(n23949), .CLK(clk), .Q(reg_file[1179]) );
  DFFPOSX1 reg_file_reg_9__28_ ( .D(n23948), .CLK(clk), .Q(reg_file[1180]) );
  DFFPOSX1 reg_file_reg_9__29_ ( .D(n23947), .CLK(clk), .Q(reg_file[1181]) );
  DFFPOSX1 reg_file_reg_9__30_ ( .D(n23946), .CLK(clk), .Q(reg_file[1182]) );
  DFFPOSX1 reg_file_reg_9__31_ ( .D(n23945), .CLK(clk), .Q(reg_file[1183]) );
  DFFPOSX1 reg_file_reg_9__32_ ( .D(n23944), .CLK(clk), .Q(reg_file[1184]) );
  DFFPOSX1 reg_file_reg_9__33_ ( .D(n23943), .CLK(clk), .Q(reg_file[1185]) );
  DFFPOSX1 reg_file_reg_9__34_ ( .D(n23942), .CLK(clk), .Q(reg_file[1186]) );
  DFFPOSX1 reg_file_reg_9__35_ ( .D(n23941), .CLK(clk), .Q(reg_file[1187]) );
  DFFPOSX1 reg_file_reg_9__36_ ( .D(n23940), .CLK(clk), .Q(reg_file[1188]) );
  DFFPOSX1 reg_file_reg_9__37_ ( .D(n23939), .CLK(clk), .Q(reg_file[1189]) );
  DFFPOSX1 reg_file_reg_9__38_ ( .D(n23938), .CLK(clk), .Q(reg_file[1190]) );
  DFFPOSX1 reg_file_reg_9__39_ ( .D(n23937), .CLK(clk), .Q(reg_file[1191]) );
  DFFPOSX1 reg_file_reg_9__40_ ( .D(n23936), .CLK(clk), .Q(reg_file[1192]) );
  DFFPOSX1 reg_file_reg_9__41_ ( .D(n23935), .CLK(clk), .Q(reg_file[1193]) );
  DFFPOSX1 reg_file_reg_9__42_ ( .D(n23934), .CLK(clk), .Q(reg_file[1194]) );
  DFFPOSX1 reg_file_reg_9__43_ ( .D(n23933), .CLK(clk), .Q(reg_file[1195]) );
  DFFPOSX1 reg_file_reg_9__44_ ( .D(n23932), .CLK(clk), .Q(reg_file[1196]) );
  DFFPOSX1 reg_file_reg_9__45_ ( .D(n23931), .CLK(clk), .Q(reg_file[1197]) );
  DFFPOSX1 reg_file_reg_9__46_ ( .D(n23930), .CLK(clk), .Q(reg_file[1198]) );
  DFFPOSX1 reg_file_reg_9__47_ ( .D(n23929), .CLK(clk), .Q(reg_file[1199]) );
  DFFPOSX1 reg_file_reg_9__48_ ( .D(n23928), .CLK(clk), .Q(reg_file[1200]) );
  DFFPOSX1 reg_file_reg_9__49_ ( .D(n23927), .CLK(clk), .Q(reg_file[1201]) );
  DFFPOSX1 reg_file_reg_9__50_ ( .D(n23926), .CLK(clk), .Q(reg_file[1202]) );
  DFFPOSX1 reg_file_reg_9__51_ ( .D(n23925), .CLK(clk), .Q(reg_file[1203]) );
  DFFPOSX1 reg_file_reg_9__52_ ( .D(n23924), .CLK(clk), .Q(reg_file[1204]) );
  DFFPOSX1 reg_file_reg_9__53_ ( .D(n23923), .CLK(clk), .Q(reg_file[1205]) );
  DFFPOSX1 reg_file_reg_9__54_ ( .D(n23922), .CLK(clk), .Q(reg_file[1206]) );
  DFFPOSX1 reg_file_reg_9__55_ ( .D(n23921), .CLK(clk), .Q(reg_file[1207]) );
  DFFPOSX1 reg_file_reg_9__56_ ( .D(n23920), .CLK(clk), .Q(reg_file[1208]) );
  DFFPOSX1 reg_file_reg_9__57_ ( .D(n23919), .CLK(clk), .Q(reg_file[1209]) );
  DFFPOSX1 reg_file_reg_9__58_ ( .D(n23918), .CLK(clk), .Q(reg_file[1210]) );
  DFFPOSX1 reg_file_reg_9__59_ ( .D(n23917), .CLK(clk), .Q(reg_file[1211]) );
  DFFPOSX1 reg_file_reg_9__60_ ( .D(n23916), .CLK(clk), .Q(reg_file[1212]) );
  DFFPOSX1 reg_file_reg_9__61_ ( .D(n23915), .CLK(clk), .Q(reg_file[1213]) );
  DFFPOSX1 reg_file_reg_9__62_ ( .D(n23914), .CLK(clk), .Q(reg_file[1214]) );
  DFFPOSX1 reg_file_reg_9__63_ ( .D(n23913), .CLK(clk), .Q(reg_file[1215]) );
  DFFPOSX1 reg_file_reg_9__64_ ( .D(n23912), .CLK(clk), .Q(reg_file[1216]) );
  DFFPOSX1 reg_file_reg_9__65_ ( .D(n23911), .CLK(clk), .Q(reg_file[1217]) );
  DFFPOSX1 reg_file_reg_9__66_ ( .D(n23910), .CLK(clk), .Q(reg_file[1218]) );
  DFFPOSX1 reg_file_reg_9__67_ ( .D(n23909), .CLK(clk), .Q(reg_file[1219]) );
  DFFPOSX1 reg_file_reg_9__68_ ( .D(n23908), .CLK(clk), .Q(reg_file[1220]) );
  DFFPOSX1 reg_file_reg_9__69_ ( .D(n23907), .CLK(clk), .Q(reg_file[1221]) );
  DFFPOSX1 reg_file_reg_9__70_ ( .D(n23906), .CLK(clk), .Q(reg_file[1222]) );
  DFFPOSX1 reg_file_reg_9__71_ ( .D(n23905), .CLK(clk), .Q(reg_file[1223]) );
  DFFPOSX1 reg_file_reg_9__72_ ( .D(n23904), .CLK(clk), .Q(reg_file[1224]) );
  DFFPOSX1 reg_file_reg_9__73_ ( .D(n23903), .CLK(clk), .Q(reg_file[1225]) );
  DFFPOSX1 reg_file_reg_9__74_ ( .D(n23902), .CLK(clk), .Q(reg_file[1226]) );
  DFFPOSX1 reg_file_reg_9__75_ ( .D(n23901), .CLK(clk), .Q(reg_file[1227]) );
  DFFPOSX1 reg_file_reg_9__76_ ( .D(n23900), .CLK(clk), .Q(reg_file[1228]) );
  DFFPOSX1 reg_file_reg_9__77_ ( .D(n23899), .CLK(clk), .Q(reg_file[1229]) );
  DFFPOSX1 reg_file_reg_9__78_ ( .D(n23898), .CLK(clk), .Q(reg_file[1230]) );
  DFFPOSX1 reg_file_reg_9__79_ ( .D(n23897), .CLK(clk), .Q(reg_file[1231]) );
  DFFPOSX1 reg_file_reg_9__80_ ( .D(n23896), .CLK(clk), .Q(reg_file[1232]) );
  DFFPOSX1 reg_file_reg_9__81_ ( .D(n23895), .CLK(clk), .Q(reg_file[1233]) );
  DFFPOSX1 reg_file_reg_9__82_ ( .D(n23894), .CLK(clk), .Q(reg_file[1234]) );
  DFFPOSX1 reg_file_reg_9__83_ ( .D(n23893), .CLK(clk), .Q(reg_file[1235]) );
  DFFPOSX1 reg_file_reg_9__84_ ( .D(n23892), .CLK(clk), .Q(reg_file[1236]) );
  DFFPOSX1 reg_file_reg_9__85_ ( .D(n23891), .CLK(clk), .Q(reg_file[1237]) );
  DFFPOSX1 reg_file_reg_9__86_ ( .D(n23890), .CLK(clk), .Q(reg_file[1238]) );
  DFFPOSX1 reg_file_reg_9__87_ ( .D(n23889), .CLK(clk), .Q(reg_file[1239]) );
  DFFPOSX1 reg_file_reg_9__88_ ( .D(n23888), .CLK(clk), .Q(reg_file[1240]) );
  DFFPOSX1 reg_file_reg_9__89_ ( .D(n23887), .CLK(clk), .Q(reg_file[1241]) );
  DFFPOSX1 reg_file_reg_9__90_ ( .D(n23886), .CLK(clk), .Q(reg_file[1242]) );
  DFFPOSX1 reg_file_reg_9__91_ ( .D(n23885), .CLK(clk), .Q(reg_file[1243]) );
  DFFPOSX1 reg_file_reg_9__92_ ( .D(n23884), .CLK(clk), .Q(reg_file[1244]) );
  DFFPOSX1 reg_file_reg_9__93_ ( .D(n23883), .CLK(clk), .Q(reg_file[1245]) );
  DFFPOSX1 reg_file_reg_9__94_ ( .D(n23882), .CLK(clk), .Q(reg_file[1246]) );
  DFFPOSX1 reg_file_reg_9__95_ ( .D(n23881), .CLK(clk), .Q(reg_file[1247]) );
  DFFPOSX1 reg_file_reg_9__96_ ( .D(n23880), .CLK(clk), .Q(reg_file[1248]) );
  DFFPOSX1 reg_file_reg_9__97_ ( .D(n23879), .CLK(clk), .Q(reg_file[1249]) );
  DFFPOSX1 reg_file_reg_9__98_ ( .D(n23878), .CLK(clk), .Q(reg_file[1250]) );
  DFFPOSX1 reg_file_reg_9__99_ ( .D(n23877), .CLK(clk), .Q(reg_file[1251]) );
  DFFPOSX1 reg_file_reg_9__100_ ( .D(n23876), .CLK(clk), .Q(reg_file[1252]) );
  DFFPOSX1 reg_file_reg_9__101_ ( .D(n23875), .CLK(clk), .Q(reg_file[1253]) );
  DFFPOSX1 reg_file_reg_9__102_ ( .D(n23874), .CLK(clk), .Q(reg_file[1254]) );
  DFFPOSX1 reg_file_reg_9__103_ ( .D(n23873), .CLK(clk), .Q(reg_file[1255]) );
  DFFPOSX1 reg_file_reg_9__104_ ( .D(n23872), .CLK(clk), .Q(reg_file[1256]) );
  DFFPOSX1 reg_file_reg_9__105_ ( .D(n23871), .CLK(clk), .Q(reg_file[1257]) );
  DFFPOSX1 reg_file_reg_9__106_ ( .D(n23870), .CLK(clk), .Q(reg_file[1258]) );
  DFFPOSX1 reg_file_reg_9__107_ ( .D(n23869), .CLK(clk), .Q(reg_file[1259]) );
  DFFPOSX1 reg_file_reg_9__108_ ( .D(n23868), .CLK(clk), .Q(reg_file[1260]) );
  DFFPOSX1 reg_file_reg_9__109_ ( .D(n23867), .CLK(clk), .Q(reg_file[1261]) );
  DFFPOSX1 reg_file_reg_9__110_ ( .D(n23866), .CLK(clk), .Q(reg_file[1262]) );
  DFFPOSX1 reg_file_reg_9__111_ ( .D(n23865), .CLK(clk), .Q(reg_file[1263]) );
  DFFPOSX1 reg_file_reg_9__112_ ( .D(n23864), .CLK(clk), .Q(reg_file[1264]) );
  DFFPOSX1 reg_file_reg_9__113_ ( .D(n23863), .CLK(clk), .Q(reg_file[1265]) );
  DFFPOSX1 reg_file_reg_9__114_ ( .D(n23862), .CLK(clk), .Q(reg_file[1266]) );
  DFFPOSX1 reg_file_reg_9__115_ ( .D(n23861), .CLK(clk), .Q(reg_file[1267]) );
  DFFPOSX1 reg_file_reg_9__116_ ( .D(n23860), .CLK(clk), .Q(reg_file[1268]) );
  DFFPOSX1 reg_file_reg_9__117_ ( .D(n23859), .CLK(clk), .Q(reg_file[1269]) );
  DFFPOSX1 reg_file_reg_9__118_ ( .D(n23858), .CLK(clk), .Q(reg_file[1270]) );
  DFFPOSX1 reg_file_reg_9__119_ ( .D(n23857), .CLK(clk), .Q(reg_file[1271]) );
  DFFPOSX1 reg_file_reg_9__120_ ( .D(n23856), .CLK(clk), .Q(reg_file[1272]) );
  DFFPOSX1 reg_file_reg_9__121_ ( .D(n23855), .CLK(clk), .Q(reg_file[1273]) );
  DFFPOSX1 reg_file_reg_9__122_ ( .D(n23854), .CLK(clk), .Q(reg_file[1274]) );
  DFFPOSX1 reg_file_reg_9__123_ ( .D(n23853), .CLK(clk), .Q(reg_file[1275]) );
  DFFPOSX1 reg_file_reg_9__124_ ( .D(n23852), .CLK(clk), .Q(reg_file[1276]) );
  DFFPOSX1 reg_file_reg_9__125_ ( .D(n23851), .CLK(clk), .Q(reg_file[1277]) );
  DFFPOSX1 reg_file_reg_9__126_ ( .D(n23850), .CLK(clk), .Q(reg_file[1278]) );
  DFFPOSX1 reg_file_reg_9__127_ ( .D(n23849), .CLK(clk), .Q(reg_file[1279]) );
  DFFPOSX1 reg_file_reg_10__0_ ( .D(n23848), .CLK(clk), .Q(reg_file[1280]) );
  DFFPOSX1 reg_file_reg_10__1_ ( .D(n23847), .CLK(clk), .Q(reg_file[1281]) );
  DFFPOSX1 reg_file_reg_10__2_ ( .D(n23846), .CLK(clk), .Q(reg_file[1282]) );
  DFFPOSX1 reg_file_reg_10__3_ ( .D(n23845), .CLK(clk), .Q(reg_file[1283]) );
  DFFPOSX1 reg_file_reg_10__4_ ( .D(n23844), .CLK(clk), .Q(reg_file[1284]) );
  DFFPOSX1 reg_file_reg_10__5_ ( .D(n23843), .CLK(clk), .Q(reg_file[1285]) );
  DFFPOSX1 reg_file_reg_10__6_ ( .D(n23842), .CLK(clk), .Q(reg_file[1286]) );
  DFFPOSX1 reg_file_reg_10__7_ ( .D(n23841), .CLK(clk), .Q(reg_file[1287]) );
  DFFPOSX1 reg_file_reg_10__8_ ( .D(n23840), .CLK(clk), .Q(reg_file[1288]) );
  DFFPOSX1 reg_file_reg_10__9_ ( .D(n23839), .CLK(clk), .Q(reg_file[1289]) );
  DFFPOSX1 reg_file_reg_10__10_ ( .D(n23838), .CLK(clk), .Q(reg_file[1290]) );
  DFFPOSX1 reg_file_reg_10__11_ ( .D(n23837), .CLK(clk), .Q(reg_file[1291]) );
  DFFPOSX1 reg_file_reg_10__12_ ( .D(n23836), .CLK(clk), .Q(reg_file[1292]) );
  DFFPOSX1 reg_file_reg_10__13_ ( .D(n23835), .CLK(clk), .Q(reg_file[1293]) );
  DFFPOSX1 reg_file_reg_10__14_ ( .D(n23834), .CLK(clk), .Q(reg_file[1294]) );
  DFFPOSX1 reg_file_reg_10__15_ ( .D(n23833), .CLK(clk), .Q(reg_file[1295]) );
  DFFPOSX1 reg_file_reg_10__16_ ( .D(n23832), .CLK(clk), .Q(reg_file[1296]) );
  DFFPOSX1 reg_file_reg_10__17_ ( .D(n23831), .CLK(clk), .Q(reg_file[1297]) );
  DFFPOSX1 reg_file_reg_10__18_ ( .D(n23830), .CLK(clk), .Q(reg_file[1298]) );
  DFFPOSX1 reg_file_reg_10__19_ ( .D(n23829), .CLK(clk), .Q(reg_file[1299]) );
  DFFPOSX1 reg_file_reg_10__20_ ( .D(n23828), .CLK(clk), .Q(reg_file[1300]) );
  DFFPOSX1 reg_file_reg_10__21_ ( .D(n23827), .CLK(clk), .Q(reg_file[1301]) );
  DFFPOSX1 reg_file_reg_10__22_ ( .D(n23826), .CLK(clk), .Q(reg_file[1302]) );
  DFFPOSX1 reg_file_reg_10__23_ ( .D(n23825), .CLK(clk), .Q(reg_file[1303]) );
  DFFPOSX1 reg_file_reg_10__24_ ( .D(n23824), .CLK(clk), .Q(reg_file[1304]) );
  DFFPOSX1 reg_file_reg_10__25_ ( .D(n23823), .CLK(clk), .Q(reg_file[1305]) );
  DFFPOSX1 reg_file_reg_10__26_ ( .D(n23822), .CLK(clk), .Q(reg_file[1306]) );
  DFFPOSX1 reg_file_reg_10__27_ ( .D(n23821), .CLK(clk), .Q(reg_file[1307]) );
  DFFPOSX1 reg_file_reg_10__28_ ( .D(n23820), .CLK(clk), .Q(reg_file[1308]) );
  DFFPOSX1 reg_file_reg_10__29_ ( .D(n23819), .CLK(clk), .Q(reg_file[1309]) );
  DFFPOSX1 reg_file_reg_10__30_ ( .D(n23818), .CLK(clk), .Q(reg_file[1310]) );
  DFFPOSX1 reg_file_reg_10__31_ ( .D(n23817), .CLK(clk), .Q(reg_file[1311]) );
  DFFPOSX1 reg_file_reg_10__32_ ( .D(n23816), .CLK(clk), .Q(reg_file[1312]) );
  DFFPOSX1 reg_file_reg_10__33_ ( .D(n23815), .CLK(clk), .Q(reg_file[1313]) );
  DFFPOSX1 reg_file_reg_10__34_ ( .D(n23814), .CLK(clk), .Q(reg_file[1314]) );
  DFFPOSX1 reg_file_reg_10__35_ ( .D(n23813), .CLK(clk), .Q(reg_file[1315]) );
  DFFPOSX1 reg_file_reg_10__36_ ( .D(n23812), .CLK(clk), .Q(reg_file[1316]) );
  DFFPOSX1 reg_file_reg_10__37_ ( .D(n23811), .CLK(clk), .Q(reg_file[1317]) );
  DFFPOSX1 reg_file_reg_10__38_ ( .D(n23810), .CLK(clk), .Q(reg_file[1318]) );
  DFFPOSX1 reg_file_reg_10__39_ ( .D(n23809), .CLK(clk), .Q(reg_file[1319]) );
  DFFPOSX1 reg_file_reg_10__40_ ( .D(n23808), .CLK(clk), .Q(reg_file[1320]) );
  DFFPOSX1 reg_file_reg_10__41_ ( .D(n23807), .CLK(clk), .Q(reg_file[1321]) );
  DFFPOSX1 reg_file_reg_10__42_ ( .D(n23806), .CLK(clk), .Q(reg_file[1322]) );
  DFFPOSX1 reg_file_reg_10__43_ ( .D(n23805), .CLK(clk), .Q(reg_file[1323]) );
  DFFPOSX1 reg_file_reg_10__44_ ( .D(n23804), .CLK(clk), .Q(reg_file[1324]) );
  DFFPOSX1 reg_file_reg_10__45_ ( .D(n23803), .CLK(clk), .Q(reg_file[1325]) );
  DFFPOSX1 reg_file_reg_10__46_ ( .D(n23802), .CLK(clk), .Q(reg_file[1326]) );
  DFFPOSX1 reg_file_reg_10__47_ ( .D(n23801), .CLK(clk), .Q(reg_file[1327]) );
  DFFPOSX1 reg_file_reg_10__48_ ( .D(n23800), .CLK(clk), .Q(reg_file[1328]) );
  DFFPOSX1 reg_file_reg_10__49_ ( .D(n23799), .CLK(clk), .Q(reg_file[1329]) );
  DFFPOSX1 reg_file_reg_10__50_ ( .D(n23798), .CLK(clk), .Q(reg_file[1330]) );
  DFFPOSX1 reg_file_reg_10__51_ ( .D(n23797), .CLK(clk), .Q(reg_file[1331]) );
  DFFPOSX1 reg_file_reg_10__52_ ( .D(n23796), .CLK(clk), .Q(reg_file[1332]) );
  DFFPOSX1 reg_file_reg_10__53_ ( .D(n23795), .CLK(clk), .Q(reg_file[1333]) );
  DFFPOSX1 reg_file_reg_10__54_ ( .D(n23794), .CLK(clk), .Q(reg_file[1334]) );
  DFFPOSX1 reg_file_reg_10__55_ ( .D(n23793), .CLK(clk), .Q(reg_file[1335]) );
  DFFPOSX1 reg_file_reg_10__56_ ( .D(n23792), .CLK(clk), .Q(reg_file[1336]) );
  DFFPOSX1 reg_file_reg_10__57_ ( .D(n23791), .CLK(clk), .Q(reg_file[1337]) );
  DFFPOSX1 reg_file_reg_10__58_ ( .D(n23790), .CLK(clk), .Q(reg_file[1338]) );
  DFFPOSX1 reg_file_reg_10__59_ ( .D(n23789), .CLK(clk), .Q(reg_file[1339]) );
  DFFPOSX1 reg_file_reg_10__60_ ( .D(n23788), .CLK(clk), .Q(reg_file[1340]) );
  DFFPOSX1 reg_file_reg_10__61_ ( .D(n23787), .CLK(clk), .Q(reg_file[1341]) );
  DFFPOSX1 reg_file_reg_10__62_ ( .D(n23786), .CLK(clk), .Q(reg_file[1342]) );
  DFFPOSX1 reg_file_reg_10__63_ ( .D(n23785), .CLK(clk), .Q(reg_file[1343]) );
  DFFPOSX1 reg_file_reg_10__64_ ( .D(n23784), .CLK(clk), .Q(reg_file[1344]) );
  DFFPOSX1 reg_file_reg_10__65_ ( .D(n23783), .CLK(clk), .Q(reg_file[1345]) );
  DFFPOSX1 reg_file_reg_10__66_ ( .D(n23782), .CLK(clk), .Q(reg_file[1346]) );
  DFFPOSX1 reg_file_reg_10__67_ ( .D(n23781), .CLK(clk), .Q(reg_file[1347]) );
  DFFPOSX1 reg_file_reg_10__68_ ( .D(n23780), .CLK(clk), .Q(reg_file[1348]) );
  DFFPOSX1 reg_file_reg_10__69_ ( .D(n23779), .CLK(clk), .Q(reg_file[1349]) );
  DFFPOSX1 reg_file_reg_10__70_ ( .D(n23778), .CLK(clk), .Q(reg_file[1350]) );
  DFFPOSX1 reg_file_reg_10__71_ ( .D(n23777), .CLK(clk), .Q(reg_file[1351]) );
  DFFPOSX1 reg_file_reg_10__72_ ( .D(n23776), .CLK(clk), .Q(reg_file[1352]) );
  DFFPOSX1 reg_file_reg_10__73_ ( .D(n23775), .CLK(clk), .Q(reg_file[1353]) );
  DFFPOSX1 reg_file_reg_10__74_ ( .D(n23774), .CLK(clk), .Q(reg_file[1354]) );
  DFFPOSX1 reg_file_reg_10__75_ ( .D(n23773), .CLK(clk), .Q(reg_file[1355]) );
  DFFPOSX1 reg_file_reg_10__76_ ( .D(n23772), .CLK(clk), .Q(reg_file[1356]) );
  DFFPOSX1 reg_file_reg_10__77_ ( .D(n23771), .CLK(clk), .Q(reg_file[1357]) );
  DFFPOSX1 reg_file_reg_10__78_ ( .D(n23770), .CLK(clk), .Q(reg_file[1358]) );
  DFFPOSX1 reg_file_reg_10__79_ ( .D(n23769), .CLK(clk), .Q(reg_file[1359]) );
  DFFPOSX1 reg_file_reg_10__80_ ( .D(n23768), .CLK(clk), .Q(reg_file[1360]) );
  DFFPOSX1 reg_file_reg_10__81_ ( .D(n23767), .CLK(clk), .Q(reg_file[1361]) );
  DFFPOSX1 reg_file_reg_10__82_ ( .D(n23766), .CLK(clk), .Q(reg_file[1362]) );
  DFFPOSX1 reg_file_reg_10__83_ ( .D(n23765), .CLK(clk), .Q(reg_file[1363]) );
  DFFPOSX1 reg_file_reg_10__84_ ( .D(n23764), .CLK(clk), .Q(reg_file[1364]) );
  DFFPOSX1 reg_file_reg_10__85_ ( .D(n23763), .CLK(clk), .Q(reg_file[1365]) );
  DFFPOSX1 reg_file_reg_10__86_ ( .D(n23762), .CLK(clk), .Q(reg_file[1366]) );
  DFFPOSX1 reg_file_reg_10__87_ ( .D(n23761), .CLK(clk), .Q(reg_file[1367]) );
  DFFPOSX1 reg_file_reg_10__88_ ( .D(n23760), .CLK(clk), .Q(reg_file[1368]) );
  DFFPOSX1 reg_file_reg_10__89_ ( .D(n23759), .CLK(clk), .Q(reg_file[1369]) );
  DFFPOSX1 reg_file_reg_10__90_ ( .D(n23758), .CLK(clk), .Q(reg_file[1370]) );
  DFFPOSX1 reg_file_reg_10__91_ ( .D(n23757), .CLK(clk), .Q(reg_file[1371]) );
  DFFPOSX1 reg_file_reg_10__92_ ( .D(n23756), .CLK(clk), .Q(reg_file[1372]) );
  DFFPOSX1 reg_file_reg_10__93_ ( .D(n23755), .CLK(clk), .Q(reg_file[1373]) );
  DFFPOSX1 reg_file_reg_10__94_ ( .D(n23754), .CLK(clk), .Q(reg_file[1374]) );
  DFFPOSX1 reg_file_reg_10__95_ ( .D(n23753), .CLK(clk), .Q(reg_file[1375]) );
  DFFPOSX1 reg_file_reg_10__96_ ( .D(n23752), .CLK(clk), .Q(reg_file[1376]) );
  DFFPOSX1 reg_file_reg_10__97_ ( .D(n23751), .CLK(clk), .Q(reg_file[1377]) );
  DFFPOSX1 reg_file_reg_10__98_ ( .D(n23750), .CLK(clk), .Q(reg_file[1378]) );
  DFFPOSX1 reg_file_reg_10__99_ ( .D(n23749), .CLK(clk), .Q(reg_file[1379]) );
  DFFPOSX1 reg_file_reg_10__100_ ( .D(n23748), .CLK(clk), .Q(reg_file[1380])
         );
  DFFPOSX1 reg_file_reg_10__101_ ( .D(n23747), .CLK(clk), .Q(reg_file[1381])
         );
  DFFPOSX1 reg_file_reg_10__102_ ( .D(n23746), .CLK(clk), .Q(reg_file[1382])
         );
  DFFPOSX1 reg_file_reg_10__103_ ( .D(n23745), .CLK(clk), .Q(reg_file[1383])
         );
  DFFPOSX1 reg_file_reg_10__104_ ( .D(n23744), .CLK(clk), .Q(reg_file[1384])
         );
  DFFPOSX1 reg_file_reg_10__105_ ( .D(n23743), .CLK(clk), .Q(reg_file[1385])
         );
  DFFPOSX1 reg_file_reg_10__106_ ( .D(n23742), .CLK(clk), .Q(reg_file[1386])
         );
  DFFPOSX1 reg_file_reg_10__107_ ( .D(n23741), .CLK(clk), .Q(reg_file[1387])
         );
  DFFPOSX1 reg_file_reg_10__108_ ( .D(n23740), .CLK(clk), .Q(reg_file[1388])
         );
  DFFPOSX1 reg_file_reg_10__109_ ( .D(n23739), .CLK(clk), .Q(reg_file[1389])
         );
  DFFPOSX1 reg_file_reg_10__110_ ( .D(n23738), .CLK(clk), .Q(reg_file[1390])
         );
  DFFPOSX1 reg_file_reg_10__111_ ( .D(n23737), .CLK(clk), .Q(reg_file[1391])
         );
  DFFPOSX1 reg_file_reg_10__112_ ( .D(n23736), .CLK(clk), .Q(reg_file[1392])
         );
  DFFPOSX1 reg_file_reg_10__113_ ( .D(n23735), .CLK(clk), .Q(reg_file[1393])
         );
  DFFPOSX1 reg_file_reg_10__114_ ( .D(n23734), .CLK(clk), .Q(reg_file[1394])
         );
  DFFPOSX1 reg_file_reg_10__115_ ( .D(n23733), .CLK(clk), .Q(reg_file[1395])
         );
  DFFPOSX1 reg_file_reg_10__116_ ( .D(n23732), .CLK(clk), .Q(reg_file[1396])
         );
  DFFPOSX1 reg_file_reg_10__117_ ( .D(n23731), .CLK(clk), .Q(reg_file[1397])
         );
  DFFPOSX1 reg_file_reg_10__118_ ( .D(n23730), .CLK(clk), .Q(reg_file[1398])
         );
  DFFPOSX1 reg_file_reg_10__119_ ( .D(n23729), .CLK(clk), .Q(reg_file[1399])
         );
  DFFPOSX1 reg_file_reg_10__120_ ( .D(n23728), .CLK(clk), .Q(reg_file[1400])
         );
  DFFPOSX1 reg_file_reg_10__121_ ( .D(n23727), .CLK(clk), .Q(reg_file[1401])
         );
  DFFPOSX1 reg_file_reg_10__122_ ( .D(n23726), .CLK(clk), .Q(reg_file[1402])
         );
  DFFPOSX1 reg_file_reg_10__123_ ( .D(n23725), .CLK(clk), .Q(reg_file[1403])
         );
  DFFPOSX1 reg_file_reg_10__124_ ( .D(n23724), .CLK(clk), .Q(reg_file[1404])
         );
  DFFPOSX1 reg_file_reg_10__125_ ( .D(n23723), .CLK(clk), .Q(reg_file[1405])
         );
  DFFPOSX1 reg_file_reg_10__126_ ( .D(n23722), .CLK(clk), .Q(reg_file[1406])
         );
  DFFPOSX1 reg_file_reg_10__127_ ( .D(n23721), .CLK(clk), .Q(reg_file[1407])
         );
  DFFPOSX1 reg_file_reg_11__0_ ( .D(n23720), .CLK(clk), .Q(reg_file[1408]) );
  DFFPOSX1 reg_file_reg_11__1_ ( .D(n23719), .CLK(clk), .Q(reg_file[1409]) );
  DFFPOSX1 reg_file_reg_11__2_ ( .D(n23718), .CLK(clk), .Q(reg_file[1410]) );
  DFFPOSX1 reg_file_reg_11__3_ ( .D(n23717), .CLK(clk), .Q(reg_file[1411]) );
  DFFPOSX1 reg_file_reg_11__4_ ( .D(n23716), .CLK(clk), .Q(reg_file[1412]) );
  DFFPOSX1 reg_file_reg_11__5_ ( .D(n23715), .CLK(clk), .Q(reg_file[1413]) );
  DFFPOSX1 reg_file_reg_11__6_ ( .D(n23714), .CLK(clk), .Q(reg_file[1414]) );
  DFFPOSX1 reg_file_reg_11__7_ ( .D(n23713), .CLK(clk), .Q(reg_file[1415]) );
  DFFPOSX1 reg_file_reg_11__8_ ( .D(n23712), .CLK(clk), .Q(reg_file[1416]) );
  DFFPOSX1 reg_file_reg_11__9_ ( .D(n23711), .CLK(clk), .Q(reg_file[1417]) );
  DFFPOSX1 reg_file_reg_11__10_ ( .D(n23710), .CLK(clk), .Q(reg_file[1418]) );
  DFFPOSX1 reg_file_reg_11__11_ ( .D(n23709), .CLK(clk), .Q(reg_file[1419]) );
  DFFPOSX1 reg_file_reg_11__12_ ( .D(n23708), .CLK(clk), .Q(reg_file[1420]) );
  DFFPOSX1 reg_file_reg_11__13_ ( .D(n23707), .CLK(clk), .Q(reg_file[1421]) );
  DFFPOSX1 reg_file_reg_11__14_ ( .D(n23706), .CLK(clk), .Q(reg_file[1422]) );
  DFFPOSX1 reg_file_reg_11__15_ ( .D(n23705), .CLK(clk), .Q(reg_file[1423]) );
  DFFPOSX1 reg_file_reg_11__16_ ( .D(n23704), .CLK(clk), .Q(reg_file[1424]) );
  DFFPOSX1 reg_file_reg_11__17_ ( .D(n23703), .CLK(clk), .Q(reg_file[1425]) );
  DFFPOSX1 reg_file_reg_11__18_ ( .D(n23702), .CLK(clk), .Q(reg_file[1426]) );
  DFFPOSX1 reg_file_reg_11__19_ ( .D(n23701), .CLK(clk), .Q(reg_file[1427]) );
  DFFPOSX1 reg_file_reg_11__20_ ( .D(n23700), .CLK(clk), .Q(reg_file[1428]) );
  DFFPOSX1 reg_file_reg_11__21_ ( .D(n23699), .CLK(clk), .Q(reg_file[1429]) );
  DFFPOSX1 reg_file_reg_11__22_ ( .D(n23698), .CLK(clk), .Q(reg_file[1430]) );
  DFFPOSX1 reg_file_reg_11__23_ ( .D(n23697), .CLK(clk), .Q(reg_file[1431]) );
  DFFPOSX1 reg_file_reg_11__24_ ( .D(n23696), .CLK(clk), .Q(reg_file[1432]) );
  DFFPOSX1 reg_file_reg_11__25_ ( .D(n23695), .CLK(clk), .Q(reg_file[1433]) );
  DFFPOSX1 reg_file_reg_11__26_ ( .D(n23694), .CLK(clk), .Q(reg_file[1434]) );
  DFFPOSX1 reg_file_reg_11__27_ ( .D(n23693), .CLK(clk), .Q(reg_file[1435]) );
  DFFPOSX1 reg_file_reg_11__28_ ( .D(n23692), .CLK(clk), .Q(reg_file[1436]) );
  DFFPOSX1 reg_file_reg_11__29_ ( .D(n23691), .CLK(clk), .Q(reg_file[1437]) );
  DFFPOSX1 reg_file_reg_11__30_ ( .D(n23690), .CLK(clk), .Q(reg_file[1438]) );
  DFFPOSX1 reg_file_reg_11__31_ ( .D(n23689), .CLK(clk), .Q(reg_file[1439]) );
  DFFPOSX1 reg_file_reg_11__32_ ( .D(n23688), .CLK(clk), .Q(reg_file[1440]) );
  DFFPOSX1 reg_file_reg_11__33_ ( .D(n23687), .CLK(clk), .Q(reg_file[1441]) );
  DFFPOSX1 reg_file_reg_11__34_ ( .D(n23686), .CLK(clk), .Q(reg_file[1442]) );
  DFFPOSX1 reg_file_reg_11__35_ ( .D(n23685), .CLK(clk), .Q(reg_file[1443]) );
  DFFPOSX1 reg_file_reg_11__36_ ( .D(n23684), .CLK(clk), .Q(reg_file[1444]) );
  DFFPOSX1 reg_file_reg_11__37_ ( .D(n23683), .CLK(clk), .Q(reg_file[1445]) );
  DFFPOSX1 reg_file_reg_11__38_ ( .D(n23682), .CLK(clk), .Q(reg_file[1446]) );
  DFFPOSX1 reg_file_reg_11__39_ ( .D(n23681), .CLK(clk), .Q(reg_file[1447]) );
  DFFPOSX1 reg_file_reg_11__40_ ( .D(n23680), .CLK(clk), .Q(reg_file[1448]) );
  DFFPOSX1 reg_file_reg_11__41_ ( .D(n23679), .CLK(clk), .Q(reg_file[1449]) );
  DFFPOSX1 reg_file_reg_11__42_ ( .D(n23678), .CLK(clk), .Q(reg_file[1450]) );
  DFFPOSX1 reg_file_reg_11__43_ ( .D(n23677), .CLK(clk), .Q(reg_file[1451]) );
  DFFPOSX1 reg_file_reg_11__44_ ( .D(n23676), .CLK(clk), .Q(reg_file[1452]) );
  DFFPOSX1 reg_file_reg_11__45_ ( .D(n23675), .CLK(clk), .Q(reg_file[1453]) );
  DFFPOSX1 reg_file_reg_11__46_ ( .D(n23674), .CLK(clk), .Q(reg_file[1454]) );
  DFFPOSX1 reg_file_reg_11__47_ ( .D(n23673), .CLK(clk), .Q(reg_file[1455]) );
  DFFPOSX1 reg_file_reg_11__48_ ( .D(n23672), .CLK(clk), .Q(reg_file[1456]) );
  DFFPOSX1 reg_file_reg_11__49_ ( .D(n23671), .CLK(clk), .Q(reg_file[1457]) );
  DFFPOSX1 reg_file_reg_11__50_ ( .D(n23670), .CLK(clk), .Q(reg_file[1458]) );
  DFFPOSX1 reg_file_reg_11__51_ ( .D(n23669), .CLK(clk), .Q(reg_file[1459]) );
  DFFPOSX1 reg_file_reg_11__52_ ( .D(n23668), .CLK(clk), .Q(reg_file[1460]) );
  DFFPOSX1 reg_file_reg_11__53_ ( .D(n23667), .CLK(clk), .Q(reg_file[1461]) );
  DFFPOSX1 reg_file_reg_11__54_ ( .D(n23666), .CLK(clk), .Q(reg_file[1462]) );
  DFFPOSX1 reg_file_reg_11__55_ ( .D(n23665), .CLK(clk), .Q(reg_file[1463]) );
  DFFPOSX1 reg_file_reg_11__56_ ( .D(n23664), .CLK(clk), .Q(reg_file[1464]) );
  DFFPOSX1 reg_file_reg_11__57_ ( .D(n23663), .CLK(clk), .Q(reg_file[1465]) );
  DFFPOSX1 reg_file_reg_11__58_ ( .D(n23662), .CLK(clk), .Q(reg_file[1466]) );
  DFFPOSX1 reg_file_reg_11__59_ ( .D(n23661), .CLK(clk), .Q(reg_file[1467]) );
  DFFPOSX1 reg_file_reg_11__60_ ( .D(n23660), .CLK(clk), .Q(reg_file[1468]) );
  DFFPOSX1 reg_file_reg_11__61_ ( .D(n23659), .CLK(clk), .Q(reg_file[1469]) );
  DFFPOSX1 reg_file_reg_11__62_ ( .D(n23658), .CLK(clk), .Q(reg_file[1470]) );
  DFFPOSX1 reg_file_reg_11__63_ ( .D(n23657), .CLK(clk), .Q(reg_file[1471]) );
  DFFPOSX1 reg_file_reg_11__64_ ( .D(n23656), .CLK(clk), .Q(reg_file[1472]) );
  DFFPOSX1 reg_file_reg_11__65_ ( .D(n23655), .CLK(clk), .Q(reg_file[1473]) );
  DFFPOSX1 reg_file_reg_11__66_ ( .D(n23654), .CLK(clk), .Q(reg_file[1474]) );
  DFFPOSX1 reg_file_reg_11__67_ ( .D(n23653), .CLK(clk), .Q(reg_file[1475]) );
  DFFPOSX1 reg_file_reg_11__68_ ( .D(n23652), .CLK(clk), .Q(reg_file[1476]) );
  DFFPOSX1 reg_file_reg_11__69_ ( .D(n23651), .CLK(clk), .Q(reg_file[1477]) );
  DFFPOSX1 reg_file_reg_11__70_ ( .D(n23650), .CLK(clk), .Q(reg_file[1478]) );
  DFFPOSX1 reg_file_reg_11__71_ ( .D(n23649), .CLK(clk), .Q(reg_file[1479]) );
  DFFPOSX1 reg_file_reg_11__72_ ( .D(n23648), .CLK(clk), .Q(reg_file[1480]) );
  DFFPOSX1 reg_file_reg_11__73_ ( .D(n23647), .CLK(clk), .Q(reg_file[1481]) );
  DFFPOSX1 reg_file_reg_11__74_ ( .D(n23646), .CLK(clk), .Q(reg_file[1482]) );
  DFFPOSX1 reg_file_reg_11__75_ ( .D(n23645), .CLK(clk), .Q(reg_file[1483]) );
  DFFPOSX1 reg_file_reg_11__76_ ( .D(n23644), .CLK(clk), .Q(reg_file[1484]) );
  DFFPOSX1 reg_file_reg_11__77_ ( .D(n23643), .CLK(clk), .Q(reg_file[1485]) );
  DFFPOSX1 reg_file_reg_11__78_ ( .D(n23642), .CLK(clk), .Q(reg_file[1486]) );
  DFFPOSX1 reg_file_reg_11__79_ ( .D(n23641), .CLK(clk), .Q(reg_file[1487]) );
  DFFPOSX1 reg_file_reg_11__80_ ( .D(n23640), .CLK(clk), .Q(reg_file[1488]) );
  DFFPOSX1 reg_file_reg_11__81_ ( .D(n23639), .CLK(clk), .Q(reg_file[1489]) );
  DFFPOSX1 reg_file_reg_11__82_ ( .D(n23638), .CLK(clk), .Q(reg_file[1490]) );
  DFFPOSX1 reg_file_reg_11__83_ ( .D(n23637), .CLK(clk), .Q(reg_file[1491]) );
  DFFPOSX1 reg_file_reg_11__84_ ( .D(n23636), .CLK(clk), .Q(reg_file[1492]) );
  DFFPOSX1 reg_file_reg_11__85_ ( .D(n23635), .CLK(clk), .Q(reg_file[1493]) );
  DFFPOSX1 reg_file_reg_11__86_ ( .D(n23634), .CLK(clk), .Q(reg_file[1494]) );
  DFFPOSX1 reg_file_reg_11__87_ ( .D(n23633), .CLK(clk), .Q(reg_file[1495]) );
  DFFPOSX1 reg_file_reg_11__88_ ( .D(n23632), .CLK(clk), .Q(reg_file[1496]) );
  DFFPOSX1 reg_file_reg_11__89_ ( .D(n23631), .CLK(clk), .Q(reg_file[1497]) );
  DFFPOSX1 reg_file_reg_11__90_ ( .D(n23630), .CLK(clk), .Q(reg_file[1498]) );
  DFFPOSX1 reg_file_reg_11__91_ ( .D(n23629), .CLK(clk), .Q(reg_file[1499]) );
  DFFPOSX1 reg_file_reg_11__92_ ( .D(n23628), .CLK(clk), .Q(reg_file[1500]) );
  DFFPOSX1 reg_file_reg_11__93_ ( .D(n23627), .CLK(clk), .Q(reg_file[1501]) );
  DFFPOSX1 reg_file_reg_11__94_ ( .D(n23626), .CLK(clk), .Q(reg_file[1502]) );
  DFFPOSX1 reg_file_reg_11__95_ ( .D(n23625), .CLK(clk), .Q(reg_file[1503]) );
  DFFPOSX1 reg_file_reg_11__96_ ( .D(n23624), .CLK(clk), .Q(reg_file[1504]) );
  DFFPOSX1 reg_file_reg_11__97_ ( .D(n23623), .CLK(clk), .Q(reg_file[1505]) );
  DFFPOSX1 reg_file_reg_11__98_ ( .D(n23622), .CLK(clk), .Q(reg_file[1506]) );
  DFFPOSX1 reg_file_reg_11__99_ ( .D(n23621), .CLK(clk), .Q(reg_file[1507]) );
  DFFPOSX1 reg_file_reg_11__100_ ( .D(n23620), .CLK(clk), .Q(reg_file[1508])
         );
  DFFPOSX1 reg_file_reg_11__101_ ( .D(n23619), .CLK(clk), .Q(reg_file[1509])
         );
  DFFPOSX1 reg_file_reg_11__102_ ( .D(n23618), .CLK(clk), .Q(reg_file[1510])
         );
  DFFPOSX1 reg_file_reg_11__103_ ( .D(n23617), .CLK(clk), .Q(reg_file[1511])
         );
  DFFPOSX1 reg_file_reg_11__104_ ( .D(n23616), .CLK(clk), .Q(reg_file[1512])
         );
  DFFPOSX1 reg_file_reg_11__105_ ( .D(n23615), .CLK(clk), .Q(reg_file[1513])
         );
  DFFPOSX1 reg_file_reg_11__106_ ( .D(n23614), .CLK(clk), .Q(reg_file[1514])
         );
  DFFPOSX1 reg_file_reg_11__107_ ( .D(n23613), .CLK(clk), .Q(reg_file[1515])
         );
  DFFPOSX1 reg_file_reg_11__108_ ( .D(n23612), .CLK(clk), .Q(reg_file[1516])
         );
  DFFPOSX1 reg_file_reg_11__109_ ( .D(n23611), .CLK(clk), .Q(reg_file[1517])
         );
  DFFPOSX1 reg_file_reg_11__110_ ( .D(n23610), .CLK(clk), .Q(reg_file[1518])
         );
  DFFPOSX1 reg_file_reg_11__111_ ( .D(n23609), .CLK(clk), .Q(reg_file[1519])
         );
  DFFPOSX1 reg_file_reg_11__112_ ( .D(n23608), .CLK(clk), .Q(reg_file[1520])
         );
  DFFPOSX1 reg_file_reg_11__113_ ( .D(n23607), .CLK(clk), .Q(reg_file[1521])
         );
  DFFPOSX1 reg_file_reg_11__114_ ( .D(n23606), .CLK(clk), .Q(reg_file[1522])
         );
  DFFPOSX1 reg_file_reg_11__115_ ( .D(n23605), .CLK(clk), .Q(reg_file[1523])
         );
  DFFPOSX1 reg_file_reg_11__116_ ( .D(n23604), .CLK(clk), .Q(reg_file[1524])
         );
  DFFPOSX1 reg_file_reg_11__117_ ( .D(n23603), .CLK(clk), .Q(reg_file[1525])
         );
  DFFPOSX1 reg_file_reg_11__118_ ( .D(n23602), .CLK(clk), .Q(reg_file[1526])
         );
  DFFPOSX1 reg_file_reg_11__119_ ( .D(n23601), .CLK(clk), .Q(reg_file[1527])
         );
  DFFPOSX1 reg_file_reg_11__120_ ( .D(n23600), .CLK(clk), .Q(reg_file[1528])
         );
  DFFPOSX1 reg_file_reg_11__121_ ( .D(n23599), .CLK(clk), .Q(reg_file[1529])
         );
  DFFPOSX1 reg_file_reg_11__122_ ( .D(n23598), .CLK(clk), .Q(reg_file[1530])
         );
  DFFPOSX1 reg_file_reg_11__123_ ( .D(n23597), .CLK(clk), .Q(reg_file[1531])
         );
  DFFPOSX1 reg_file_reg_11__124_ ( .D(n23596), .CLK(clk), .Q(reg_file[1532])
         );
  DFFPOSX1 reg_file_reg_11__125_ ( .D(n23595), .CLK(clk), .Q(reg_file[1533])
         );
  DFFPOSX1 reg_file_reg_11__126_ ( .D(n23594), .CLK(clk), .Q(reg_file[1534])
         );
  DFFPOSX1 reg_file_reg_11__127_ ( .D(n23593), .CLK(clk), .Q(reg_file[1535])
         );
  DFFPOSX1 reg_file_reg_12__0_ ( .D(n23592), .CLK(clk), .Q(reg_file[1536]) );
  DFFPOSX1 reg_file_reg_12__1_ ( .D(n23591), .CLK(clk), .Q(reg_file[1537]) );
  DFFPOSX1 reg_file_reg_12__2_ ( .D(n23590), .CLK(clk), .Q(reg_file[1538]) );
  DFFPOSX1 reg_file_reg_12__3_ ( .D(n23589), .CLK(clk), .Q(reg_file[1539]) );
  DFFPOSX1 reg_file_reg_12__4_ ( .D(n23588), .CLK(clk), .Q(reg_file[1540]) );
  DFFPOSX1 reg_file_reg_12__5_ ( .D(n23587), .CLK(clk), .Q(reg_file[1541]) );
  DFFPOSX1 reg_file_reg_12__6_ ( .D(n23586), .CLK(clk), .Q(reg_file[1542]) );
  DFFPOSX1 reg_file_reg_12__7_ ( .D(n23585), .CLK(clk), .Q(reg_file[1543]) );
  DFFPOSX1 reg_file_reg_12__8_ ( .D(n23584), .CLK(clk), .Q(reg_file[1544]) );
  DFFPOSX1 reg_file_reg_12__9_ ( .D(n23583), .CLK(clk), .Q(reg_file[1545]) );
  DFFPOSX1 reg_file_reg_12__10_ ( .D(n23582), .CLK(clk), .Q(reg_file[1546]) );
  DFFPOSX1 reg_file_reg_12__11_ ( .D(n23581), .CLK(clk), .Q(reg_file[1547]) );
  DFFPOSX1 reg_file_reg_12__12_ ( .D(n23580), .CLK(clk), .Q(reg_file[1548]) );
  DFFPOSX1 reg_file_reg_12__13_ ( .D(n23579), .CLK(clk), .Q(reg_file[1549]) );
  DFFPOSX1 reg_file_reg_12__14_ ( .D(n23578), .CLK(clk), .Q(reg_file[1550]) );
  DFFPOSX1 reg_file_reg_12__15_ ( .D(n23577), .CLK(clk), .Q(reg_file[1551]) );
  DFFPOSX1 reg_file_reg_12__16_ ( .D(n23576), .CLK(clk), .Q(reg_file[1552]) );
  DFFPOSX1 reg_file_reg_12__17_ ( .D(n23575), .CLK(clk), .Q(reg_file[1553]) );
  DFFPOSX1 reg_file_reg_12__18_ ( .D(n23574), .CLK(clk), .Q(reg_file[1554]) );
  DFFPOSX1 reg_file_reg_12__19_ ( .D(n23573), .CLK(clk), .Q(reg_file[1555]) );
  DFFPOSX1 reg_file_reg_12__20_ ( .D(n23572), .CLK(clk), .Q(reg_file[1556]) );
  DFFPOSX1 reg_file_reg_12__21_ ( .D(n23571), .CLK(clk), .Q(reg_file[1557]) );
  DFFPOSX1 reg_file_reg_12__22_ ( .D(n23570), .CLK(clk), .Q(reg_file[1558]) );
  DFFPOSX1 reg_file_reg_12__23_ ( .D(n23569), .CLK(clk), .Q(reg_file[1559]) );
  DFFPOSX1 reg_file_reg_12__24_ ( .D(n23568), .CLK(clk), .Q(reg_file[1560]) );
  DFFPOSX1 reg_file_reg_12__25_ ( .D(n23567), .CLK(clk), .Q(reg_file[1561]) );
  DFFPOSX1 reg_file_reg_12__26_ ( .D(n23566), .CLK(clk), .Q(reg_file[1562]) );
  DFFPOSX1 reg_file_reg_12__27_ ( .D(n23565), .CLK(clk), .Q(reg_file[1563]) );
  DFFPOSX1 reg_file_reg_12__28_ ( .D(n23564), .CLK(clk), .Q(reg_file[1564]) );
  DFFPOSX1 reg_file_reg_12__29_ ( .D(n23563), .CLK(clk), .Q(reg_file[1565]) );
  DFFPOSX1 reg_file_reg_12__30_ ( .D(n23562), .CLK(clk), .Q(reg_file[1566]) );
  DFFPOSX1 reg_file_reg_12__31_ ( .D(n23561), .CLK(clk), .Q(reg_file[1567]) );
  DFFPOSX1 reg_file_reg_12__32_ ( .D(n23560), .CLK(clk), .Q(reg_file[1568]) );
  DFFPOSX1 reg_file_reg_12__33_ ( .D(n23559), .CLK(clk), .Q(reg_file[1569]) );
  DFFPOSX1 reg_file_reg_12__34_ ( .D(n23558), .CLK(clk), .Q(reg_file[1570]) );
  DFFPOSX1 reg_file_reg_12__35_ ( .D(n23557), .CLK(clk), .Q(reg_file[1571]) );
  DFFPOSX1 reg_file_reg_12__36_ ( .D(n23556), .CLK(clk), .Q(reg_file[1572]) );
  DFFPOSX1 reg_file_reg_12__37_ ( .D(n23555), .CLK(clk), .Q(reg_file[1573]) );
  DFFPOSX1 reg_file_reg_12__38_ ( .D(n23554), .CLK(clk), .Q(reg_file[1574]) );
  DFFPOSX1 reg_file_reg_12__39_ ( .D(n23553), .CLK(clk), .Q(reg_file[1575]) );
  DFFPOSX1 reg_file_reg_12__40_ ( .D(n23552), .CLK(clk), .Q(reg_file[1576]) );
  DFFPOSX1 reg_file_reg_12__41_ ( .D(n23551), .CLK(clk), .Q(reg_file[1577]) );
  DFFPOSX1 reg_file_reg_12__42_ ( .D(n23550), .CLK(clk), .Q(reg_file[1578]) );
  DFFPOSX1 reg_file_reg_12__43_ ( .D(n23549), .CLK(clk), .Q(reg_file[1579]) );
  DFFPOSX1 reg_file_reg_12__44_ ( .D(n23548), .CLK(clk), .Q(reg_file[1580]) );
  DFFPOSX1 reg_file_reg_12__45_ ( .D(n23547), .CLK(clk), .Q(reg_file[1581]) );
  DFFPOSX1 reg_file_reg_12__46_ ( .D(n23546), .CLK(clk), .Q(reg_file[1582]) );
  DFFPOSX1 reg_file_reg_12__47_ ( .D(n23545), .CLK(clk), .Q(reg_file[1583]) );
  DFFPOSX1 reg_file_reg_12__48_ ( .D(n23544), .CLK(clk), .Q(reg_file[1584]) );
  DFFPOSX1 reg_file_reg_12__49_ ( .D(n23543), .CLK(clk), .Q(reg_file[1585]) );
  DFFPOSX1 reg_file_reg_12__50_ ( .D(n23542), .CLK(clk), .Q(reg_file[1586]) );
  DFFPOSX1 reg_file_reg_12__51_ ( .D(n23541), .CLK(clk), .Q(reg_file[1587]) );
  DFFPOSX1 reg_file_reg_12__52_ ( .D(n23540), .CLK(clk), .Q(reg_file[1588]) );
  DFFPOSX1 reg_file_reg_12__53_ ( .D(n23539), .CLK(clk), .Q(reg_file[1589]) );
  DFFPOSX1 reg_file_reg_12__54_ ( .D(n23538), .CLK(clk), .Q(reg_file[1590]) );
  DFFPOSX1 reg_file_reg_12__55_ ( .D(n23537), .CLK(clk), .Q(reg_file[1591]) );
  DFFPOSX1 reg_file_reg_12__56_ ( .D(n23536), .CLK(clk), .Q(reg_file[1592]) );
  DFFPOSX1 reg_file_reg_12__57_ ( .D(n23535), .CLK(clk), .Q(reg_file[1593]) );
  DFFPOSX1 reg_file_reg_12__58_ ( .D(n23534), .CLK(clk), .Q(reg_file[1594]) );
  DFFPOSX1 reg_file_reg_12__59_ ( .D(n23533), .CLK(clk), .Q(reg_file[1595]) );
  DFFPOSX1 reg_file_reg_12__60_ ( .D(n23532), .CLK(clk), .Q(reg_file[1596]) );
  DFFPOSX1 reg_file_reg_12__61_ ( .D(n23531), .CLK(clk), .Q(reg_file[1597]) );
  DFFPOSX1 reg_file_reg_12__62_ ( .D(n23530), .CLK(clk), .Q(reg_file[1598]) );
  DFFPOSX1 reg_file_reg_12__63_ ( .D(n23529), .CLK(clk), .Q(reg_file[1599]) );
  DFFPOSX1 reg_file_reg_12__64_ ( .D(n23528), .CLK(clk), .Q(reg_file[1600]) );
  DFFPOSX1 reg_file_reg_12__65_ ( .D(n23527), .CLK(clk), .Q(reg_file[1601]) );
  DFFPOSX1 reg_file_reg_12__66_ ( .D(n23526), .CLK(clk), .Q(reg_file[1602]) );
  DFFPOSX1 reg_file_reg_12__67_ ( .D(n23525), .CLK(clk), .Q(reg_file[1603]) );
  DFFPOSX1 reg_file_reg_12__68_ ( .D(n23524), .CLK(clk), .Q(reg_file[1604]) );
  DFFPOSX1 reg_file_reg_12__69_ ( .D(n23523), .CLK(clk), .Q(reg_file[1605]) );
  DFFPOSX1 reg_file_reg_12__70_ ( .D(n23522), .CLK(clk), .Q(reg_file[1606]) );
  DFFPOSX1 reg_file_reg_12__71_ ( .D(n23521), .CLK(clk), .Q(reg_file[1607]) );
  DFFPOSX1 reg_file_reg_12__72_ ( .D(n23520), .CLK(clk), .Q(reg_file[1608]) );
  DFFPOSX1 reg_file_reg_12__73_ ( .D(n23519), .CLK(clk), .Q(reg_file[1609]) );
  DFFPOSX1 reg_file_reg_12__74_ ( .D(n23518), .CLK(clk), .Q(reg_file[1610]) );
  DFFPOSX1 reg_file_reg_12__75_ ( .D(n23517), .CLK(clk), .Q(reg_file[1611]) );
  DFFPOSX1 reg_file_reg_12__76_ ( .D(n23516), .CLK(clk), .Q(reg_file[1612]) );
  DFFPOSX1 reg_file_reg_12__77_ ( .D(n23515), .CLK(clk), .Q(reg_file[1613]) );
  DFFPOSX1 reg_file_reg_12__78_ ( .D(n23514), .CLK(clk), .Q(reg_file[1614]) );
  DFFPOSX1 reg_file_reg_12__79_ ( .D(n23513), .CLK(clk), .Q(reg_file[1615]) );
  DFFPOSX1 reg_file_reg_12__80_ ( .D(n23512), .CLK(clk), .Q(reg_file[1616]) );
  DFFPOSX1 reg_file_reg_12__81_ ( .D(n23511), .CLK(clk), .Q(reg_file[1617]) );
  DFFPOSX1 reg_file_reg_12__82_ ( .D(n23510), .CLK(clk), .Q(reg_file[1618]) );
  DFFPOSX1 reg_file_reg_12__83_ ( .D(n23509), .CLK(clk), .Q(reg_file[1619]) );
  DFFPOSX1 reg_file_reg_12__84_ ( .D(n23508), .CLK(clk), .Q(reg_file[1620]) );
  DFFPOSX1 reg_file_reg_12__85_ ( .D(n23507), .CLK(clk), .Q(reg_file[1621]) );
  DFFPOSX1 reg_file_reg_12__86_ ( .D(n23506), .CLK(clk), .Q(reg_file[1622]) );
  DFFPOSX1 reg_file_reg_12__87_ ( .D(n23505), .CLK(clk), .Q(reg_file[1623]) );
  DFFPOSX1 reg_file_reg_12__88_ ( .D(n23504), .CLK(clk), .Q(reg_file[1624]) );
  DFFPOSX1 reg_file_reg_12__89_ ( .D(n23503), .CLK(clk), .Q(reg_file[1625]) );
  DFFPOSX1 reg_file_reg_12__90_ ( .D(n23502), .CLK(clk), .Q(reg_file[1626]) );
  DFFPOSX1 reg_file_reg_12__91_ ( .D(n23501), .CLK(clk), .Q(reg_file[1627]) );
  DFFPOSX1 reg_file_reg_12__92_ ( .D(n23500), .CLK(clk), .Q(reg_file[1628]) );
  DFFPOSX1 reg_file_reg_12__93_ ( .D(n23499), .CLK(clk), .Q(reg_file[1629]) );
  DFFPOSX1 reg_file_reg_12__94_ ( .D(n23498), .CLK(clk), .Q(reg_file[1630]) );
  DFFPOSX1 reg_file_reg_12__95_ ( .D(n23497), .CLK(clk), .Q(reg_file[1631]) );
  DFFPOSX1 reg_file_reg_12__96_ ( .D(n23496), .CLK(clk), .Q(reg_file[1632]) );
  DFFPOSX1 reg_file_reg_12__97_ ( .D(n23495), .CLK(clk), .Q(reg_file[1633]) );
  DFFPOSX1 reg_file_reg_12__98_ ( .D(n23494), .CLK(clk), .Q(reg_file[1634]) );
  DFFPOSX1 reg_file_reg_12__99_ ( .D(n23493), .CLK(clk), .Q(reg_file[1635]) );
  DFFPOSX1 reg_file_reg_12__100_ ( .D(n23492), .CLK(clk), .Q(reg_file[1636])
         );
  DFFPOSX1 reg_file_reg_12__101_ ( .D(n23491), .CLK(clk), .Q(reg_file[1637])
         );
  DFFPOSX1 reg_file_reg_12__102_ ( .D(n23490), .CLK(clk), .Q(reg_file[1638])
         );
  DFFPOSX1 reg_file_reg_12__103_ ( .D(n23489), .CLK(clk), .Q(reg_file[1639])
         );
  DFFPOSX1 reg_file_reg_12__104_ ( .D(n23488), .CLK(clk), .Q(reg_file[1640])
         );
  DFFPOSX1 reg_file_reg_12__105_ ( .D(n23487), .CLK(clk), .Q(reg_file[1641])
         );
  DFFPOSX1 reg_file_reg_12__106_ ( .D(n23486), .CLK(clk), .Q(reg_file[1642])
         );
  DFFPOSX1 reg_file_reg_12__107_ ( .D(n23485), .CLK(clk), .Q(reg_file[1643])
         );
  DFFPOSX1 reg_file_reg_12__108_ ( .D(n23484), .CLK(clk), .Q(reg_file[1644])
         );
  DFFPOSX1 reg_file_reg_12__109_ ( .D(n23483), .CLK(clk), .Q(reg_file[1645])
         );
  DFFPOSX1 reg_file_reg_12__110_ ( .D(n23482), .CLK(clk), .Q(reg_file[1646])
         );
  DFFPOSX1 reg_file_reg_12__111_ ( .D(n23481), .CLK(clk), .Q(reg_file[1647])
         );
  DFFPOSX1 reg_file_reg_12__112_ ( .D(n23480), .CLK(clk), .Q(reg_file[1648])
         );
  DFFPOSX1 reg_file_reg_12__113_ ( .D(n23479), .CLK(clk), .Q(reg_file[1649])
         );
  DFFPOSX1 reg_file_reg_12__114_ ( .D(n23478), .CLK(clk), .Q(reg_file[1650])
         );
  DFFPOSX1 reg_file_reg_12__115_ ( .D(n23477), .CLK(clk), .Q(reg_file[1651])
         );
  DFFPOSX1 reg_file_reg_12__116_ ( .D(n23476), .CLK(clk), .Q(reg_file[1652])
         );
  DFFPOSX1 reg_file_reg_12__117_ ( .D(n23475), .CLK(clk), .Q(reg_file[1653])
         );
  DFFPOSX1 reg_file_reg_12__118_ ( .D(n23474), .CLK(clk), .Q(reg_file[1654])
         );
  DFFPOSX1 reg_file_reg_12__119_ ( .D(n23473), .CLK(clk), .Q(reg_file[1655])
         );
  DFFPOSX1 reg_file_reg_12__120_ ( .D(n23472), .CLK(clk), .Q(reg_file[1656])
         );
  DFFPOSX1 reg_file_reg_12__121_ ( .D(n23471), .CLK(clk), .Q(reg_file[1657])
         );
  DFFPOSX1 reg_file_reg_12__122_ ( .D(n23470), .CLK(clk), .Q(reg_file[1658])
         );
  DFFPOSX1 reg_file_reg_12__123_ ( .D(n23469), .CLK(clk), .Q(reg_file[1659])
         );
  DFFPOSX1 reg_file_reg_12__124_ ( .D(n23468), .CLK(clk), .Q(reg_file[1660])
         );
  DFFPOSX1 reg_file_reg_12__125_ ( .D(n23467), .CLK(clk), .Q(reg_file[1661])
         );
  DFFPOSX1 reg_file_reg_12__126_ ( .D(n23466), .CLK(clk), .Q(reg_file[1662])
         );
  DFFPOSX1 reg_file_reg_12__127_ ( .D(n23465), .CLK(clk), .Q(reg_file[1663])
         );
  DFFPOSX1 reg_file_reg_13__0_ ( .D(n23464), .CLK(clk), .Q(reg_file[1664]) );
  DFFPOSX1 reg_file_reg_13__1_ ( .D(n23463), .CLK(clk), .Q(reg_file[1665]) );
  DFFPOSX1 reg_file_reg_13__2_ ( .D(n23462), .CLK(clk), .Q(reg_file[1666]) );
  DFFPOSX1 reg_file_reg_13__3_ ( .D(n23461), .CLK(clk), .Q(reg_file[1667]) );
  DFFPOSX1 reg_file_reg_13__4_ ( .D(n23460), .CLK(clk), .Q(reg_file[1668]) );
  DFFPOSX1 reg_file_reg_13__5_ ( .D(n23459), .CLK(clk), .Q(reg_file[1669]) );
  DFFPOSX1 reg_file_reg_13__6_ ( .D(n23458), .CLK(clk), .Q(reg_file[1670]) );
  DFFPOSX1 reg_file_reg_13__7_ ( .D(n23457), .CLK(clk), .Q(reg_file[1671]) );
  DFFPOSX1 reg_file_reg_13__8_ ( .D(n23456), .CLK(clk), .Q(reg_file[1672]) );
  DFFPOSX1 reg_file_reg_13__9_ ( .D(n23455), .CLK(clk), .Q(reg_file[1673]) );
  DFFPOSX1 reg_file_reg_13__10_ ( .D(n23454), .CLK(clk), .Q(reg_file[1674]) );
  DFFPOSX1 reg_file_reg_13__11_ ( .D(n23453), .CLK(clk), .Q(reg_file[1675]) );
  DFFPOSX1 reg_file_reg_13__12_ ( .D(n23452), .CLK(clk), .Q(reg_file[1676]) );
  DFFPOSX1 reg_file_reg_13__13_ ( .D(n23451), .CLK(clk), .Q(reg_file[1677]) );
  DFFPOSX1 reg_file_reg_13__14_ ( .D(n23450), .CLK(clk), .Q(reg_file[1678]) );
  DFFPOSX1 reg_file_reg_13__15_ ( .D(n23449), .CLK(clk), .Q(reg_file[1679]) );
  DFFPOSX1 reg_file_reg_13__16_ ( .D(n23448), .CLK(clk), .Q(reg_file[1680]) );
  DFFPOSX1 reg_file_reg_13__17_ ( .D(n23447), .CLK(clk), .Q(reg_file[1681]) );
  DFFPOSX1 reg_file_reg_13__18_ ( .D(n23446), .CLK(clk), .Q(reg_file[1682]) );
  DFFPOSX1 reg_file_reg_13__19_ ( .D(n23445), .CLK(clk), .Q(reg_file[1683]) );
  DFFPOSX1 reg_file_reg_13__20_ ( .D(n23444), .CLK(clk), .Q(reg_file[1684]) );
  DFFPOSX1 reg_file_reg_13__21_ ( .D(n23443), .CLK(clk), .Q(reg_file[1685]) );
  DFFPOSX1 reg_file_reg_13__22_ ( .D(n23442), .CLK(clk), .Q(reg_file[1686]) );
  DFFPOSX1 reg_file_reg_13__23_ ( .D(n23441), .CLK(clk), .Q(reg_file[1687]) );
  DFFPOSX1 reg_file_reg_13__24_ ( .D(n23440), .CLK(clk), .Q(reg_file[1688]) );
  DFFPOSX1 reg_file_reg_13__25_ ( .D(n23439), .CLK(clk), .Q(reg_file[1689]) );
  DFFPOSX1 reg_file_reg_13__26_ ( .D(n23438), .CLK(clk), .Q(reg_file[1690]) );
  DFFPOSX1 reg_file_reg_13__27_ ( .D(n23437), .CLK(clk), .Q(reg_file[1691]) );
  DFFPOSX1 reg_file_reg_13__28_ ( .D(n23436), .CLK(clk), .Q(reg_file[1692]) );
  DFFPOSX1 reg_file_reg_13__29_ ( .D(n23435), .CLK(clk), .Q(reg_file[1693]) );
  DFFPOSX1 reg_file_reg_13__30_ ( .D(n23434), .CLK(clk), .Q(reg_file[1694]) );
  DFFPOSX1 reg_file_reg_13__31_ ( .D(n23433), .CLK(clk), .Q(reg_file[1695]) );
  DFFPOSX1 reg_file_reg_13__32_ ( .D(n23432), .CLK(clk), .Q(reg_file[1696]) );
  DFFPOSX1 reg_file_reg_13__33_ ( .D(n23431), .CLK(clk), .Q(reg_file[1697]) );
  DFFPOSX1 reg_file_reg_13__34_ ( .D(n23430), .CLK(clk), .Q(reg_file[1698]) );
  DFFPOSX1 reg_file_reg_13__35_ ( .D(n23429), .CLK(clk), .Q(reg_file[1699]) );
  DFFPOSX1 reg_file_reg_13__36_ ( .D(n23428), .CLK(clk), .Q(reg_file[1700]) );
  DFFPOSX1 reg_file_reg_13__37_ ( .D(n23427), .CLK(clk), .Q(reg_file[1701]) );
  DFFPOSX1 reg_file_reg_13__38_ ( .D(n23426), .CLK(clk), .Q(reg_file[1702]) );
  DFFPOSX1 reg_file_reg_13__39_ ( .D(n23425), .CLK(clk), .Q(reg_file[1703]) );
  DFFPOSX1 reg_file_reg_13__40_ ( .D(n23424), .CLK(clk), .Q(reg_file[1704]) );
  DFFPOSX1 reg_file_reg_13__41_ ( .D(n23423), .CLK(clk), .Q(reg_file[1705]) );
  DFFPOSX1 reg_file_reg_13__42_ ( .D(n23422), .CLK(clk), .Q(reg_file[1706]) );
  DFFPOSX1 reg_file_reg_13__43_ ( .D(n23421), .CLK(clk), .Q(reg_file[1707]) );
  DFFPOSX1 reg_file_reg_13__44_ ( .D(n23420), .CLK(clk), .Q(reg_file[1708]) );
  DFFPOSX1 reg_file_reg_13__45_ ( .D(n23419), .CLK(clk), .Q(reg_file[1709]) );
  DFFPOSX1 reg_file_reg_13__46_ ( .D(n23418), .CLK(clk), .Q(reg_file[1710]) );
  DFFPOSX1 reg_file_reg_13__47_ ( .D(n23417), .CLK(clk), .Q(reg_file[1711]) );
  DFFPOSX1 reg_file_reg_13__48_ ( .D(n23416), .CLK(clk), .Q(reg_file[1712]) );
  DFFPOSX1 reg_file_reg_13__49_ ( .D(n23415), .CLK(clk), .Q(reg_file[1713]) );
  DFFPOSX1 reg_file_reg_13__50_ ( .D(n23414), .CLK(clk), .Q(reg_file[1714]) );
  DFFPOSX1 reg_file_reg_13__51_ ( .D(n23413), .CLK(clk), .Q(reg_file[1715]) );
  DFFPOSX1 reg_file_reg_13__52_ ( .D(n23412), .CLK(clk), .Q(reg_file[1716]) );
  DFFPOSX1 reg_file_reg_13__53_ ( .D(n23411), .CLK(clk), .Q(reg_file[1717]) );
  DFFPOSX1 reg_file_reg_13__54_ ( .D(n23410), .CLK(clk), .Q(reg_file[1718]) );
  DFFPOSX1 reg_file_reg_13__55_ ( .D(n23409), .CLK(clk), .Q(reg_file[1719]) );
  DFFPOSX1 reg_file_reg_13__56_ ( .D(n23408), .CLK(clk), .Q(reg_file[1720]) );
  DFFPOSX1 reg_file_reg_13__57_ ( .D(n23407), .CLK(clk), .Q(reg_file[1721]) );
  DFFPOSX1 reg_file_reg_13__58_ ( .D(n23406), .CLK(clk), .Q(reg_file[1722]) );
  DFFPOSX1 reg_file_reg_13__59_ ( .D(n23405), .CLK(clk), .Q(reg_file[1723]) );
  DFFPOSX1 reg_file_reg_13__60_ ( .D(n23404), .CLK(clk), .Q(reg_file[1724]) );
  DFFPOSX1 reg_file_reg_13__61_ ( .D(n23403), .CLK(clk), .Q(reg_file[1725]) );
  DFFPOSX1 reg_file_reg_13__62_ ( .D(n23402), .CLK(clk), .Q(reg_file[1726]) );
  DFFPOSX1 reg_file_reg_13__63_ ( .D(n23401), .CLK(clk), .Q(reg_file[1727]) );
  DFFPOSX1 reg_file_reg_13__64_ ( .D(n23400), .CLK(clk), .Q(reg_file[1728]) );
  DFFPOSX1 reg_file_reg_13__65_ ( .D(n23399), .CLK(clk), .Q(reg_file[1729]) );
  DFFPOSX1 reg_file_reg_13__66_ ( .D(n23398), .CLK(clk), .Q(reg_file[1730]) );
  DFFPOSX1 reg_file_reg_13__67_ ( .D(n23397), .CLK(clk), .Q(reg_file[1731]) );
  DFFPOSX1 reg_file_reg_13__68_ ( .D(n23396), .CLK(clk), .Q(reg_file[1732]) );
  DFFPOSX1 reg_file_reg_13__69_ ( .D(n23395), .CLK(clk), .Q(reg_file[1733]) );
  DFFPOSX1 reg_file_reg_13__70_ ( .D(n23394), .CLK(clk), .Q(reg_file[1734]) );
  DFFPOSX1 reg_file_reg_13__71_ ( .D(n23393), .CLK(clk), .Q(reg_file[1735]) );
  DFFPOSX1 reg_file_reg_13__72_ ( .D(n23392), .CLK(clk), .Q(reg_file[1736]) );
  DFFPOSX1 reg_file_reg_13__73_ ( .D(n23391), .CLK(clk), .Q(reg_file[1737]) );
  DFFPOSX1 reg_file_reg_13__74_ ( .D(n23390), .CLK(clk), .Q(reg_file[1738]) );
  DFFPOSX1 reg_file_reg_13__75_ ( .D(n23389), .CLK(clk), .Q(reg_file[1739]) );
  DFFPOSX1 reg_file_reg_13__76_ ( .D(n23388), .CLK(clk), .Q(reg_file[1740]) );
  DFFPOSX1 reg_file_reg_13__77_ ( .D(n23387), .CLK(clk), .Q(reg_file[1741]) );
  DFFPOSX1 reg_file_reg_13__78_ ( .D(n23386), .CLK(clk), .Q(reg_file[1742]) );
  DFFPOSX1 reg_file_reg_13__79_ ( .D(n23385), .CLK(clk), .Q(reg_file[1743]) );
  DFFPOSX1 reg_file_reg_13__80_ ( .D(n23384), .CLK(clk), .Q(reg_file[1744]) );
  DFFPOSX1 reg_file_reg_13__81_ ( .D(n23383), .CLK(clk), .Q(reg_file[1745]) );
  DFFPOSX1 reg_file_reg_13__82_ ( .D(n23382), .CLK(clk), .Q(reg_file[1746]) );
  DFFPOSX1 reg_file_reg_13__83_ ( .D(n23381), .CLK(clk), .Q(reg_file[1747]) );
  DFFPOSX1 reg_file_reg_13__84_ ( .D(n23380), .CLK(clk), .Q(reg_file[1748]) );
  DFFPOSX1 reg_file_reg_13__85_ ( .D(n23379), .CLK(clk), .Q(reg_file[1749]) );
  DFFPOSX1 reg_file_reg_13__86_ ( .D(n23378), .CLK(clk), .Q(reg_file[1750]) );
  DFFPOSX1 reg_file_reg_13__87_ ( .D(n23377), .CLK(clk), .Q(reg_file[1751]) );
  DFFPOSX1 reg_file_reg_13__88_ ( .D(n23376), .CLK(clk), .Q(reg_file[1752]) );
  DFFPOSX1 reg_file_reg_13__89_ ( .D(n23375), .CLK(clk), .Q(reg_file[1753]) );
  DFFPOSX1 reg_file_reg_13__90_ ( .D(n23374), .CLK(clk), .Q(reg_file[1754]) );
  DFFPOSX1 reg_file_reg_13__91_ ( .D(n23373), .CLK(clk), .Q(reg_file[1755]) );
  DFFPOSX1 reg_file_reg_13__92_ ( .D(n23372), .CLK(clk), .Q(reg_file[1756]) );
  DFFPOSX1 reg_file_reg_13__93_ ( .D(n23371), .CLK(clk), .Q(reg_file[1757]) );
  DFFPOSX1 reg_file_reg_13__94_ ( .D(n23370), .CLK(clk), .Q(reg_file[1758]) );
  DFFPOSX1 reg_file_reg_13__95_ ( .D(n23369), .CLK(clk), .Q(reg_file[1759]) );
  DFFPOSX1 reg_file_reg_13__96_ ( .D(n23368), .CLK(clk), .Q(reg_file[1760]) );
  DFFPOSX1 reg_file_reg_13__97_ ( .D(n23367), .CLK(clk), .Q(reg_file[1761]) );
  DFFPOSX1 reg_file_reg_13__98_ ( .D(n23366), .CLK(clk), .Q(reg_file[1762]) );
  DFFPOSX1 reg_file_reg_13__99_ ( .D(n23365), .CLK(clk), .Q(reg_file[1763]) );
  DFFPOSX1 reg_file_reg_13__100_ ( .D(n23364), .CLK(clk), .Q(reg_file[1764])
         );
  DFFPOSX1 reg_file_reg_13__101_ ( .D(n23363), .CLK(clk), .Q(reg_file[1765])
         );
  DFFPOSX1 reg_file_reg_13__102_ ( .D(n23362), .CLK(clk), .Q(reg_file[1766])
         );
  DFFPOSX1 reg_file_reg_13__103_ ( .D(n23361), .CLK(clk), .Q(reg_file[1767])
         );
  DFFPOSX1 reg_file_reg_13__104_ ( .D(n23360), .CLK(clk), .Q(reg_file[1768])
         );
  DFFPOSX1 reg_file_reg_13__105_ ( .D(n23359), .CLK(clk), .Q(reg_file[1769])
         );
  DFFPOSX1 reg_file_reg_13__106_ ( .D(n23358), .CLK(clk), .Q(reg_file[1770])
         );
  DFFPOSX1 reg_file_reg_13__107_ ( .D(n23357), .CLK(clk), .Q(reg_file[1771])
         );
  DFFPOSX1 reg_file_reg_13__108_ ( .D(n23356), .CLK(clk), .Q(reg_file[1772])
         );
  DFFPOSX1 reg_file_reg_13__109_ ( .D(n23355), .CLK(clk), .Q(reg_file[1773])
         );
  DFFPOSX1 reg_file_reg_13__110_ ( .D(n23354), .CLK(clk), .Q(reg_file[1774])
         );
  DFFPOSX1 reg_file_reg_13__111_ ( .D(n23353), .CLK(clk), .Q(reg_file[1775])
         );
  DFFPOSX1 reg_file_reg_13__112_ ( .D(n23352), .CLK(clk), .Q(reg_file[1776])
         );
  DFFPOSX1 reg_file_reg_13__113_ ( .D(n23351), .CLK(clk), .Q(reg_file[1777])
         );
  DFFPOSX1 reg_file_reg_13__114_ ( .D(n23350), .CLK(clk), .Q(reg_file[1778])
         );
  DFFPOSX1 reg_file_reg_13__115_ ( .D(n23349), .CLK(clk), .Q(reg_file[1779])
         );
  DFFPOSX1 reg_file_reg_13__116_ ( .D(n23348), .CLK(clk), .Q(reg_file[1780])
         );
  DFFPOSX1 reg_file_reg_13__117_ ( .D(n23347), .CLK(clk), .Q(reg_file[1781])
         );
  DFFPOSX1 reg_file_reg_13__118_ ( .D(n23346), .CLK(clk), .Q(reg_file[1782])
         );
  DFFPOSX1 reg_file_reg_13__119_ ( .D(n23345), .CLK(clk), .Q(reg_file[1783])
         );
  DFFPOSX1 reg_file_reg_13__120_ ( .D(n23344), .CLK(clk), .Q(reg_file[1784])
         );
  DFFPOSX1 reg_file_reg_13__121_ ( .D(n23343), .CLK(clk), .Q(reg_file[1785])
         );
  DFFPOSX1 reg_file_reg_13__122_ ( .D(n23342), .CLK(clk), .Q(reg_file[1786])
         );
  DFFPOSX1 reg_file_reg_13__123_ ( .D(n23341), .CLK(clk), .Q(reg_file[1787])
         );
  DFFPOSX1 reg_file_reg_13__124_ ( .D(n23340), .CLK(clk), .Q(reg_file[1788])
         );
  DFFPOSX1 reg_file_reg_13__125_ ( .D(n23339), .CLK(clk), .Q(reg_file[1789])
         );
  DFFPOSX1 reg_file_reg_13__126_ ( .D(n23338), .CLK(clk), .Q(reg_file[1790])
         );
  DFFPOSX1 reg_file_reg_13__127_ ( .D(n23337), .CLK(clk), .Q(reg_file[1791])
         );
  DFFPOSX1 reg_file_reg_14__0_ ( .D(n23336), .CLK(clk), .Q(reg_file[1792]) );
  DFFPOSX1 reg_file_reg_14__1_ ( .D(n23335), .CLK(clk), .Q(reg_file[1793]) );
  DFFPOSX1 reg_file_reg_14__2_ ( .D(n23334), .CLK(clk), .Q(reg_file[1794]) );
  DFFPOSX1 reg_file_reg_14__3_ ( .D(n23333), .CLK(clk), .Q(reg_file[1795]) );
  DFFPOSX1 reg_file_reg_14__4_ ( .D(n23332), .CLK(clk), .Q(reg_file[1796]) );
  DFFPOSX1 reg_file_reg_14__5_ ( .D(n23331), .CLK(clk), .Q(reg_file[1797]) );
  DFFPOSX1 reg_file_reg_14__6_ ( .D(n23330), .CLK(clk), .Q(reg_file[1798]) );
  DFFPOSX1 reg_file_reg_14__7_ ( .D(n23329), .CLK(clk), .Q(reg_file[1799]) );
  DFFPOSX1 reg_file_reg_14__8_ ( .D(n23328), .CLK(clk), .Q(reg_file[1800]) );
  DFFPOSX1 reg_file_reg_14__9_ ( .D(n23327), .CLK(clk), .Q(reg_file[1801]) );
  DFFPOSX1 reg_file_reg_14__10_ ( .D(n23326), .CLK(clk), .Q(reg_file[1802]) );
  DFFPOSX1 reg_file_reg_14__11_ ( .D(n23325), .CLK(clk), .Q(reg_file[1803]) );
  DFFPOSX1 reg_file_reg_14__12_ ( .D(n23324), .CLK(clk), .Q(reg_file[1804]) );
  DFFPOSX1 reg_file_reg_14__13_ ( .D(n23323), .CLK(clk), .Q(reg_file[1805]) );
  DFFPOSX1 reg_file_reg_14__14_ ( .D(n23322), .CLK(clk), .Q(reg_file[1806]) );
  DFFPOSX1 reg_file_reg_14__15_ ( .D(n23321), .CLK(clk), .Q(reg_file[1807]) );
  DFFPOSX1 reg_file_reg_14__16_ ( .D(n23320), .CLK(clk), .Q(reg_file[1808]) );
  DFFPOSX1 reg_file_reg_14__17_ ( .D(n23319), .CLK(clk), .Q(reg_file[1809]) );
  DFFPOSX1 reg_file_reg_14__18_ ( .D(n23318), .CLK(clk), .Q(reg_file[1810]) );
  DFFPOSX1 reg_file_reg_14__19_ ( .D(n23317), .CLK(clk), .Q(reg_file[1811]) );
  DFFPOSX1 reg_file_reg_14__20_ ( .D(n23316), .CLK(clk), .Q(reg_file[1812]) );
  DFFPOSX1 reg_file_reg_14__21_ ( .D(n23315), .CLK(clk), .Q(reg_file[1813]) );
  DFFPOSX1 reg_file_reg_14__22_ ( .D(n23314), .CLK(clk), .Q(reg_file[1814]) );
  DFFPOSX1 reg_file_reg_14__23_ ( .D(n23313), .CLK(clk), .Q(reg_file[1815]) );
  DFFPOSX1 reg_file_reg_14__24_ ( .D(n23312), .CLK(clk), .Q(reg_file[1816]) );
  DFFPOSX1 reg_file_reg_14__25_ ( .D(n23311), .CLK(clk), .Q(reg_file[1817]) );
  DFFPOSX1 reg_file_reg_14__26_ ( .D(n23310), .CLK(clk), .Q(reg_file[1818]) );
  DFFPOSX1 reg_file_reg_14__27_ ( .D(n23309), .CLK(clk), .Q(reg_file[1819]) );
  DFFPOSX1 reg_file_reg_14__28_ ( .D(n23308), .CLK(clk), .Q(reg_file[1820]) );
  DFFPOSX1 reg_file_reg_14__29_ ( .D(n23307), .CLK(clk), .Q(reg_file[1821]) );
  DFFPOSX1 reg_file_reg_14__30_ ( .D(n23306), .CLK(clk), .Q(reg_file[1822]) );
  DFFPOSX1 reg_file_reg_14__31_ ( .D(n23305), .CLK(clk), .Q(reg_file[1823]) );
  DFFPOSX1 reg_file_reg_14__32_ ( .D(n23304), .CLK(clk), .Q(reg_file[1824]) );
  DFFPOSX1 reg_file_reg_14__33_ ( .D(n23303), .CLK(clk), .Q(reg_file[1825]) );
  DFFPOSX1 reg_file_reg_14__34_ ( .D(n23302), .CLK(clk), .Q(reg_file[1826]) );
  DFFPOSX1 reg_file_reg_14__35_ ( .D(n23301), .CLK(clk), .Q(reg_file[1827]) );
  DFFPOSX1 reg_file_reg_14__36_ ( .D(n23300), .CLK(clk), .Q(reg_file[1828]) );
  DFFPOSX1 reg_file_reg_14__37_ ( .D(n23299), .CLK(clk), .Q(reg_file[1829]) );
  DFFPOSX1 reg_file_reg_14__38_ ( .D(n23298), .CLK(clk), .Q(reg_file[1830]) );
  DFFPOSX1 reg_file_reg_14__39_ ( .D(n23297), .CLK(clk), .Q(reg_file[1831]) );
  DFFPOSX1 reg_file_reg_14__40_ ( .D(n23296), .CLK(clk), .Q(reg_file[1832]) );
  DFFPOSX1 reg_file_reg_14__41_ ( .D(n23295), .CLK(clk), .Q(reg_file[1833]) );
  DFFPOSX1 reg_file_reg_14__42_ ( .D(n23294), .CLK(clk), .Q(reg_file[1834]) );
  DFFPOSX1 reg_file_reg_14__43_ ( .D(n23293), .CLK(clk), .Q(reg_file[1835]) );
  DFFPOSX1 reg_file_reg_14__44_ ( .D(n23292), .CLK(clk), .Q(reg_file[1836]) );
  DFFPOSX1 reg_file_reg_14__45_ ( .D(n23291), .CLK(clk), .Q(reg_file[1837]) );
  DFFPOSX1 reg_file_reg_14__46_ ( .D(n23290), .CLK(clk), .Q(reg_file[1838]) );
  DFFPOSX1 reg_file_reg_14__47_ ( .D(n23289), .CLK(clk), .Q(reg_file[1839]) );
  DFFPOSX1 reg_file_reg_14__48_ ( .D(n23288), .CLK(clk), .Q(reg_file[1840]) );
  DFFPOSX1 reg_file_reg_14__49_ ( .D(n23287), .CLK(clk), .Q(reg_file[1841]) );
  DFFPOSX1 reg_file_reg_14__50_ ( .D(n23286), .CLK(clk), .Q(reg_file[1842]) );
  DFFPOSX1 reg_file_reg_14__51_ ( .D(n23285), .CLK(clk), .Q(reg_file[1843]) );
  DFFPOSX1 reg_file_reg_14__52_ ( .D(n23284), .CLK(clk), .Q(reg_file[1844]) );
  DFFPOSX1 reg_file_reg_14__53_ ( .D(n23283), .CLK(clk), .Q(reg_file[1845]) );
  DFFPOSX1 reg_file_reg_14__54_ ( .D(n23282), .CLK(clk), .Q(reg_file[1846]) );
  DFFPOSX1 reg_file_reg_14__55_ ( .D(n23281), .CLK(clk), .Q(reg_file[1847]) );
  DFFPOSX1 reg_file_reg_14__56_ ( .D(n23280), .CLK(clk), .Q(reg_file[1848]) );
  DFFPOSX1 reg_file_reg_14__57_ ( .D(n23279), .CLK(clk), .Q(reg_file[1849]) );
  DFFPOSX1 reg_file_reg_14__58_ ( .D(n23278), .CLK(clk), .Q(reg_file[1850]) );
  DFFPOSX1 reg_file_reg_14__59_ ( .D(n23277), .CLK(clk), .Q(reg_file[1851]) );
  DFFPOSX1 reg_file_reg_14__60_ ( .D(n23276), .CLK(clk), .Q(reg_file[1852]) );
  DFFPOSX1 reg_file_reg_14__61_ ( .D(n23275), .CLK(clk), .Q(reg_file[1853]) );
  DFFPOSX1 reg_file_reg_14__62_ ( .D(n23274), .CLK(clk), .Q(reg_file[1854]) );
  DFFPOSX1 reg_file_reg_14__63_ ( .D(n23273), .CLK(clk), .Q(reg_file[1855]) );
  DFFPOSX1 reg_file_reg_14__64_ ( .D(n23272), .CLK(clk), .Q(reg_file[1856]) );
  DFFPOSX1 reg_file_reg_14__65_ ( .D(n23271), .CLK(clk), .Q(reg_file[1857]) );
  DFFPOSX1 reg_file_reg_14__66_ ( .D(n23270), .CLK(clk), .Q(reg_file[1858]) );
  DFFPOSX1 reg_file_reg_14__67_ ( .D(n23269), .CLK(clk), .Q(reg_file[1859]) );
  DFFPOSX1 reg_file_reg_14__68_ ( .D(n23268), .CLK(clk), .Q(reg_file[1860]) );
  DFFPOSX1 reg_file_reg_14__69_ ( .D(n23267), .CLK(clk), .Q(reg_file[1861]) );
  DFFPOSX1 reg_file_reg_14__70_ ( .D(n23266), .CLK(clk), .Q(reg_file[1862]) );
  DFFPOSX1 reg_file_reg_14__71_ ( .D(n23265), .CLK(clk), .Q(reg_file[1863]) );
  DFFPOSX1 reg_file_reg_14__72_ ( .D(n23264), .CLK(clk), .Q(reg_file[1864]) );
  DFFPOSX1 reg_file_reg_14__73_ ( .D(n23263), .CLK(clk), .Q(reg_file[1865]) );
  DFFPOSX1 reg_file_reg_14__74_ ( .D(n23262), .CLK(clk), .Q(reg_file[1866]) );
  DFFPOSX1 reg_file_reg_14__75_ ( .D(n23261), .CLK(clk), .Q(reg_file[1867]) );
  DFFPOSX1 reg_file_reg_14__76_ ( .D(n23260), .CLK(clk), .Q(reg_file[1868]) );
  DFFPOSX1 reg_file_reg_14__77_ ( .D(n23259), .CLK(clk), .Q(reg_file[1869]) );
  DFFPOSX1 reg_file_reg_14__78_ ( .D(n23258), .CLK(clk), .Q(reg_file[1870]) );
  DFFPOSX1 reg_file_reg_14__79_ ( .D(n23257), .CLK(clk), .Q(reg_file[1871]) );
  DFFPOSX1 reg_file_reg_14__80_ ( .D(n23256), .CLK(clk), .Q(reg_file[1872]) );
  DFFPOSX1 reg_file_reg_14__81_ ( .D(n23255), .CLK(clk), .Q(reg_file[1873]) );
  DFFPOSX1 reg_file_reg_14__82_ ( .D(n23254), .CLK(clk), .Q(reg_file[1874]) );
  DFFPOSX1 reg_file_reg_14__83_ ( .D(n23253), .CLK(clk), .Q(reg_file[1875]) );
  DFFPOSX1 reg_file_reg_14__84_ ( .D(n23252), .CLK(clk), .Q(reg_file[1876]) );
  DFFPOSX1 reg_file_reg_14__85_ ( .D(n23251), .CLK(clk), .Q(reg_file[1877]) );
  DFFPOSX1 reg_file_reg_14__86_ ( .D(n23250), .CLK(clk), .Q(reg_file[1878]) );
  DFFPOSX1 reg_file_reg_14__87_ ( .D(n23249), .CLK(clk), .Q(reg_file[1879]) );
  DFFPOSX1 reg_file_reg_14__88_ ( .D(n23248), .CLK(clk), .Q(reg_file[1880]) );
  DFFPOSX1 reg_file_reg_14__89_ ( .D(n23247), .CLK(clk), .Q(reg_file[1881]) );
  DFFPOSX1 reg_file_reg_14__90_ ( .D(n23246), .CLK(clk), .Q(reg_file[1882]) );
  DFFPOSX1 reg_file_reg_14__91_ ( .D(n23245), .CLK(clk), .Q(reg_file[1883]) );
  DFFPOSX1 reg_file_reg_14__92_ ( .D(n23244), .CLK(clk), .Q(reg_file[1884]) );
  DFFPOSX1 reg_file_reg_14__93_ ( .D(n23243), .CLK(clk), .Q(reg_file[1885]) );
  DFFPOSX1 reg_file_reg_14__94_ ( .D(n23242), .CLK(clk), .Q(reg_file[1886]) );
  DFFPOSX1 reg_file_reg_14__95_ ( .D(n23241), .CLK(clk), .Q(reg_file[1887]) );
  DFFPOSX1 reg_file_reg_14__96_ ( .D(n23240), .CLK(clk), .Q(reg_file[1888]) );
  DFFPOSX1 reg_file_reg_14__97_ ( .D(n23239), .CLK(clk), .Q(reg_file[1889]) );
  DFFPOSX1 reg_file_reg_14__98_ ( .D(n23238), .CLK(clk), .Q(reg_file[1890]) );
  DFFPOSX1 reg_file_reg_14__99_ ( .D(n23237), .CLK(clk), .Q(reg_file[1891]) );
  DFFPOSX1 reg_file_reg_14__100_ ( .D(n23236), .CLK(clk), .Q(reg_file[1892])
         );
  DFFPOSX1 reg_file_reg_14__101_ ( .D(n23235), .CLK(clk), .Q(reg_file[1893])
         );
  DFFPOSX1 reg_file_reg_14__102_ ( .D(n23234), .CLK(clk), .Q(reg_file[1894])
         );
  DFFPOSX1 reg_file_reg_14__103_ ( .D(n23233), .CLK(clk), .Q(reg_file[1895])
         );
  DFFPOSX1 reg_file_reg_14__104_ ( .D(n23232), .CLK(clk), .Q(reg_file[1896])
         );
  DFFPOSX1 reg_file_reg_14__105_ ( .D(n23231), .CLK(clk), .Q(reg_file[1897])
         );
  DFFPOSX1 reg_file_reg_14__106_ ( .D(n23230), .CLK(clk), .Q(reg_file[1898])
         );
  DFFPOSX1 reg_file_reg_14__107_ ( .D(n23229), .CLK(clk), .Q(reg_file[1899])
         );
  DFFPOSX1 reg_file_reg_14__108_ ( .D(n23228), .CLK(clk), .Q(reg_file[1900])
         );
  DFFPOSX1 reg_file_reg_14__109_ ( .D(n23227), .CLK(clk), .Q(reg_file[1901])
         );
  DFFPOSX1 reg_file_reg_14__110_ ( .D(n23226), .CLK(clk), .Q(reg_file[1902])
         );
  DFFPOSX1 reg_file_reg_14__111_ ( .D(n23225), .CLK(clk), .Q(reg_file[1903])
         );
  DFFPOSX1 reg_file_reg_14__112_ ( .D(n23224), .CLK(clk), .Q(reg_file[1904])
         );
  DFFPOSX1 reg_file_reg_14__113_ ( .D(n23223), .CLK(clk), .Q(reg_file[1905])
         );
  DFFPOSX1 reg_file_reg_14__114_ ( .D(n23222), .CLK(clk), .Q(reg_file[1906])
         );
  DFFPOSX1 reg_file_reg_14__115_ ( .D(n23221), .CLK(clk), .Q(reg_file[1907])
         );
  DFFPOSX1 reg_file_reg_14__116_ ( .D(n23220), .CLK(clk), .Q(reg_file[1908])
         );
  DFFPOSX1 reg_file_reg_14__117_ ( .D(n23219), .CLK(clk), .Q(reg_file[1909])
         );
  DFFPOSX1 reg_file_reg_14__118_ ( .D(n23218), .CLK(clk), .Q(reg_file[1910])
         );
  DFFPOSX1 reg_file_reg_14__119_ ( .D(n23217), .CLK(clk), .Q(reg_file[1911])
         );
  DFFPOSX1 reg_file_reg_14__120_ ( .D(n23216), .CLK(clk), .Q(reg_file[1912])
         );
  DFFPOSX1 reg_file_reg_14__121_ ( .D(n23215), .CLK(clk), .Q(reg_file[1913])
         );
  DFFPOSX1 reg_file_reg_14__122_ ( .D(n23214), .CLK(clk), .Q(reg_file[1914])
         );
  DFFPOSX1 reg_file_reg_14__123_ ( .D(n23213), .CLK(clk), .Q(reg_file[1915])
         );
  DFFPOSX1 reg_file_reg_14__124_ ( .D(n23212), .CLK(clk), .Q(reg_file[1916])
         );
  DFFPOSX1 reg_file_reg_14__125_ ( .D(n23211), .CLK(clk), .Q(reg_file[1917])
         );
  DFFPOSX1 reg_file_reg_14__126_ ( .D(n23210), .CLK(clk), .Q(reg_file[1918])
         );
  DFFPOSX1 reg_file_reg_14__127_ ( .D(n23209), .CLK(clk), .Q(reg_file[1919])
         );
  DFFPOSX1 reg_file_reg_15__0_ ( .D(n23208), .CLK(clk), .Q(reg_file[1920]) );
  DFFPOSX1 reg_file_reg_15__1_ ( .D(n23207), .CLK(clk), .Q(reg_file[1921]) );
  DFFPOSX1 reg_file_reg_15__2_ ( .D(n23206), .CLK(clk), .Q(reg_file[1922]) );
  DFFPOSX1 reg_file_reg_15__3_ ( .D(n23205), .CLK(clk), .Q(reg_file[1923]) );
  DFFPOSX1 reg_file_reg_15__4_ ( .D(n23204), .CLK(clk), .Q(reg_file[1924]) );
  DFFPOSX1 reg_file_reg_15__5_ ( .D(n23203), .CLK(clk), .Q(reg_file[1925]) );
  DFFPOSX1 reg_file_reg_15__6_ ( .D(n23202), .CLK(clk), .Q(reg_file[1926]) );
  DFFPOSX1 reg_file_reg_15__7_ ( .D(n23201), .CLK(clk), .Q(reg_file[1927]) );
  DFFPOSX1 reg_file_reg_15__8_ ( .D(n23200), .CLK(clk), .Q(reg_file[1928]) );
  DFFPOSX1 reg_file_reg_15__9_ ( .D(n23199), .CLK(clk), .Q(reg_file[1929]) );
  DFFPOSX1 reg_file_reg_15__10_ ( .D(n23198), .CLK(clk), .Q(reg_file[1930]) );
  DFFPOSX1 reg_file_reg_15__11_ ( .D(n23197), .CLK(clk), .Q(reg_file[1931]) );
  DFFPOSX1 reg_file_reg_15__12_ ( .D(n23196), .CLK(clk), .Q(reg_file[1932]) );
  DFFPOSX1 reg_file_reg_15__13_ ( .D(n23195), .CLK(clk), .Q(reg_file[1933]) );
  DFFPOSX1 reg_file_reg_15__14_ ( .D(n23194), .CLK(clk), .Q(reg_file[1934]) );
  DFFPOSX1 reg_file_reg_15__15_ ( .D(n23193), .CLK(clk), .Q(reg_file[1935]) );
  DFFPOSX1 reg_file_reg_15__16_ ( .D(n23192), .CLK(clk), .Q(reg_file[1936]) );
  DFFPOSX1 reg_file_reg_15__17_ ( .D(n23191), .CLK(clk), .Q(reg_file[1937]) );
  DFFPOSX1 reg_file_reg_15__18_ ( .D(n23190), .CLK(clk), .Q(reg_file[1938]) );
  DFFPOSX1 reg_file_reg_15__19_ ( .D(n23189), .CLK(clk), .Q(reg_file[1939]) );
  DFFPOSX1 reg_file_reg_15__20_ ( .D(n23188), .CLK(clk), .Q(reg_file[1940]) );
  DFFPOSX1 reg_file_reg_15__21_ ( .D(n23187), .CLK(clk), .Q(reg_file[1941]) );
  DFFPOSX1 reg_file_reg_15__22_ ( .D(n23186), .CLK(clk), .Q(reg_file[1942]) );
  DFFPOSX1 reg_file_reg_15__23_ ( .D(n23185), .CLK(clk), .Q(reg_file[1943]) );
  DFFPOSX1 reg_file_reg_15__24_ ( .D(n23184), .CLK(clk), .Q(reg_file[1944]) );
  DFFPOSX1 reg_file_reg_15__25_ ( .D(n23183), .CLK(clk), .Q(reg_file[1945]) );
  DFFPOSX1 reg_file_reg_15__26_ ( .D(n23182), .CLK(clk), .Q(reg_file[1946]) );
  DFFPOSX1 reg_file_reg_15__27_ ( .D(n23181), .CLK(clk), .Q(reg_file[1947]) );
  DFFPOSX1 reg_file_reg_15__28_ ( .D(n23180), .CLK(clk), .Q(reg_file[1948]) );
  DFFPOSX1 reg_file_reg_15__29_ ( .D(n23179), .CLK(clk), .Q(reg_file[1949]) );
  DFFPOSX1 reg_file_reg_15__30_ ( .D(n23178), .CLK(clk), .Q(reg_file[1950]) );
  DFFPOSX1 reg_file_reg_15__31_ ( .D(n23177), .CLK(clk), .Q(reg_file[1951]) );
  DFFPOSX1 reg_file_reg_15__32_ ( .D(n23176), .CLK(clk), .Q(reg_file[1952]) );
  DFFPOSX1 reg_file_reg_15__33_ ( .D(n23175), .CLK(clk), .Q(reg_file[1953]) );
  DFFPOSX1 reg_file_reg_15__34_ ( .D(n23174), .CLK(clk), .Q(reg_file[1954]) );
  DFFPOSX1 reg_file_reg_15__35_ ( .D(n23173), .CLK(clk), .Q(reg_file[1955]) );
  DFFPOSX1 reg_file_reg_15__36_ ( .D(n23172), .CLK(clk), .Q(reg_file[1956]) );
  DFFPOSX1 reg_file_reg_15__37_ ( .D(n23171), .CLK(clk), .Q(reg_file[1957]) );
  DFFPOSX1 reg_file_reg_15__38_ ( .D(n23170), .CLK(clk), .Q(reg_file[1958]) );
  DFFPOSX1 reg_file_reg_15__39_ ( .D(n23169), .CLK(clk), .Q(reg_file[1959]) );
  DFFPOSX1 reg_file_reg_15__40_ ( .D(n23168), .CLK(clk), .Q(reg_file[1960]) );
  DFFPOSX1 reg_file_reg_15__41_ ( .D(n23167), .CLK(clk), .Q(reg_file[1961]) );
  DFFPOSX1 reg_file_reg_15__42_ ( .D(n23166), .CLK(clk), .Q(reg_file[1962]) );
  DFFPOSX1 reg_file_reg_15__43_ ( .D(n23165), .CLK(clk), .Q(reg_file[1963]) );
  DFFPOSX1 reg_file_reg_15__44_ ( .D(n23164), .CLK(clk), .Q(reg_file[1964]) );
  DFFPOSX1 reg_file_reg_15__45_ ( .D(n23163), .CLK(clk), .Q(reg_file[1965]) );
  DFFPOSX1 reg_file_reg_15__46_ ( .D(n23162), .CLK(clk), .Q(reg_file[1966]) );
  DFFPOSX1 reg_file_reg_15__47_ ( .D(n23161), .CLK(clk), .Q(reg_file[1967]) );
  DFFPOSX1 reg_file_reg_15__48_ ( .D(n23160), .CLK(clk), .Q(reg_file[1968]) );
  DFFPOSX1 reg_file_reg_15__49_ ( .D(n23159), .CLK(clk), .Q(reg_file[1969]) );
  DFFPOSX1 reg_file_reg_15__50_ ( .D(n23158), .CLK(clk), .Q(reg_file[1970]) );
  DFFPOSX1 reg_file_reg_15__51_ ( .D(n23157), .CLK(clk), .Q(reg_file[1971]) );
  DFFPOSX1 reg_file_reg_15__52_ ( .D(n23156), .CLK(clk), .Q(reg_file[1972]) );
  DFFPOSX1 reg_file_reg_15__53_ ( .D(n23155), .CLK(clk), .Q(reg_file[1973]) );
  DFFPOSX1 reg_file_reg_15__54_ ( .D(n23154), .CLK(clk), .Q(reg_file[1974]) );
  DFFPOSX1 reg_file_reg_15__55_ ( .D(n23153), .CLK(clk), .Q(reg_file[1975]) );
  DFFPOSX1 reg_file_reg_15__56_ ( .D(n23152), .CLK(clk), .Q(reg_file[1976]) );
  DFFPOSX1 reg_file_reg_15__57_ ( .D(n23151), .CLK(clk), .Q(reg_file[1977]) );
  DFFPOSX1 reg_file_reg_15__58_ ( .D(n23150), .CLK(clk), .Q(reg_file[1978]) );
  DFFPOSX1 reg_file_reg_15__59_ ( .D(n23149), .CLK(clk), .Q(reg_file[1979]) );
  DFFPOSX1 reg_file_reg_15__60_ ( .D(n23148), .CLK(clk), .Q(reg_file[1980]) );
  DFFPOSX1 reg_file_reg_15__61_ ( .D(n23147), .CLK(clk), .Q(reg_file[1981]) );
  DFFPOSX1 reg_file_reg_15__62_ ( .D(n23146), .CLK(clk), .Q(reg_file[1982]) );
  DFFPOSX1 reg_file_reg_15__63_ ( .D(n23145), .CLK(clk), .Q(reg_file[1983]) );
  DFFPOSX1 reg_file_reg_15__64_ ( .D(n23144), .CLK(clk), .Q(reg_file[1984]) );
  DFFPOSX1 reg_file_reg_15__65_ ( .D(n23143), .CLK(clk), .Q(reg_file[1985]) );
  DFFPOSX1 reg_file_reg_15__66_ ( .D(n23142), .CLK(clk), .Q(reg_file[1986]) );
  DFFPOSX1 reg_file_reg_15__67_ ( .D(n23141), .CLK(clk), .Q(reg_file[1987]) );
  DFFPOSX1 reg_file_reg_15__68_ ( .D(n23140), .CLK(clk), .Q(reg_file[1988]) );
  DFFPOSX1 reg_file_reg_15__69_ ( .D(n23139), .CLK(clk), .Q(reg_file[1989]) );
  DFFPOSX1 reg_file_reg_15__70_ ( .D(n23138), .CLK(clk), .Q(reg_file[1990]) );
  DFFPOSX1 reg_file_reg_15__71_ ( .D(n23137), .CLK(clk), .Q(reg_file[1991]) );
  DFFPOSX1 reg_file_reg_15__72_ ( .D(n23136), .CLK(clk), .Q(reg_file[1992]) );
  DFFPOSX1 reg_file_reg_15__73_ ( .D(n23135), .CLK(clk), .Q(reg_file[1993]) );
  DFFPOSX1 reg_file_reg_15__74_ ( .D(n23134), .CLK(clk), .Q(reg_file[1994]) );
  DFFPOSX1 reg_file_reg_15__75_ ( .D(n23133), .CLK(clk), .Q(reg_file[1995]) );
  DFFPOSX1 reg_file_reg_15__76_ ( .D(n23132), .CLK(clk), .Q(reg_file[1996]) );
  DFFPOSX1 reg_file_reg_15__77_ ( .D(n23131), .CLK(clk), .Q(reg_file[1997]) );
  DFFPOSX1 reg_file_reg_15__78_ ( .D(n23130), .CLK(clk), .Q(reg_file[1998]) );
  DFFPOSX1 reg_file_reg_15__79_ ( .D(n23129), .CLK(clk), .Q(reg_file[1999]) );
  DFFPOSX1 reg_file_reg_15__80_ ( .D(n23128), .CLK(clk), .Q(reg_file[2000]) );
  DFFPOSX1 reg_file_reg_15__81_ ( .D(n23127), .CLK(clk), .Q(reg_file[2001]) );
  DFFPOSX1 reg_file_reg_15__82_ ( .D(n23126), .CLK(clk), .Q(reg_file[2002]) );
  DFFPOSX1 reg_file_reg_15__83_ ( .D(n23125), .CLK(clk), .Q(reg_file[2003]) );
  DFFPOSX1 reg_file_reg_15__84_ ( .D(n23124), .CLK(clk), .Q(reg_file[2004]) );
  DFFPOSX1 reg_file_reg_15__85_ ( .D(n23123), .CLK(clk), .Q(reg_file[2005]) );
  DFFPOSX1 reg_file_reg_15__86_ ( .D(n23122), .CLK(clk), .Q(reg_file[2006]) );
  DFFPOSX1 reg_file_reg_15__87_ ( .D(n23121), .CLK(clk), .Q(reg_file[2007]) );
  DFFPOSX1 reg_file_reg_15__88_ ( .D(n23120), .CLK(clk), .Q(reg_file[2008]) );
  DFFPOSX1 reg_file_reg_15__89_ ( .D(n23119), .CLK(clk), .Q(reg_file[2009]) );
  DFFPOSX1 reg_file_reg_15__90_ ( .D(n23118), .CLK(clk), .Q(reg_file[2010]) );
  DFFPOSX1 reg_file_reg_15__91_ ( .D(n23117), .CLK(clk), .Q(reg_file[2011]) );
  DFFPOSX1 reg_file_reg_15__92_ ( .D(n23116), .CLK(clk), .Q(reg_file[2012]) );
  DFFPOSX1 reg_file_reg_15__93_ ( .D(n23115), .CLK(clk), .Q(reg_file[2013]) );
  DFFPOSX1 reg_file_reg_15__94_ ( .D(n23114), .CLK(clk), .Q(reg_file[2014]) );
  DFFPOSX1 reg_file_reg_15__95_ ( .D(n23113), .CLK(clk), .Q(reg_file[2015]) );
  DFFPOSX1 reg_file_reg_15__96_ ( .D(n23112), .CLK(clk), .Q(reg_file[2016]) );
  DFFPOSX1 reg_file_reg_15__97_ ( .D(n23111), .CLK(clk), .Q(reg_file[2017]) );
  DFFPOSX1 reg_file_reg_15__98_ ( .D(n23110), .CLK(clk), .Q(reg_file[2018]) );
  DFFPOSX1 reg_file_reg_15__99_ ( .D(n23109), .CLK(clk), .Q(reg_file[2019]) );
  DFFPOSX1 reg_file_reg_15__100_ ( .D(n23108), .CLK(clk), .Q(reg_file[2020])
         );
  DFFPOSX1 reg_file_reg_15__101_ ( .D(n23107), .CLK(clk), .Q(reg_file[2021])
         );
  DFFPOSX1 reg_file_reg_15__102_ ( .D(n23106), .CLK(clk), .Q(reg_file[2022])
         );
  DFFPOSX1 reg_file_reg_15__103_ ( .D(n23105), .CLK(clk), .Q(reg_file[2023])
         );
  DFFPOSX1 reg_file_reg_15__104_ ( .D(n23104), .CLK(clk), .Q(reg_file[2024])
         );
  DFFPOSX1 reg_file_reg_15__105_ ( .D(n23103), .CLK(clk), .Q(reg_file[2025])
         );
  DFFPOSX1 reg_file_reg_15__106_ ( .D(n23102), .CLK(clk), .Q(reg_file[2026])
         );
  DFFPOSX1 reg_file_reg_15__107_ ( .D(n23101), .CLK(clk), .Q(reg_file[2027])
         );
  DFFPOSX1 reg_file_reg_15__108_ ( .D(n23100), .CLK(clk), .Q(reg_file[2028])
         );
  DFFPOSX1 reg_file_reg_15__109_ ( .D(n23099), .CLK(clk), .Q(reg_file[2029])
         );
  DFFPOSX1 reg_file_reg_15__110_ ( .D(n23098), .CLK(clk), .Q(reg_file[2030])
         );
  DFFPOSX1 reg_file_reg_15__111_ ( .D(n23097), .CLK(clk), .Q(reg_file[2031])
         );
  DFFPOSX1 reg_file_reg_15__112_ ( .D(n23096), .CLK(clk), .Q(reg_file[2032])
         );
  DFFPOSX1 reg_file_reg_15__113_ ( .D(n23095), .CLK(clk), .Q(reg_file[2033])
         );
  DFFPOSX1 reg_file_reg_15__114_ ( .D(n23094), .CLK(clk), .Q(reg_file[2034])
         );
  DFFPOSX1 reg_file_reg_15__115_ ( .D(n23093), .CLK(clk), .Q(reg_file[2035])
         );
  DFFPOSX1 reg_file_reg_15__116_ ( .D(n23092), .CLK(clk), .Q(reg_file[2036])
         );
  DFFPOSX1 reg_file_reg_15__117_ ( .D(n23091), .CLK(clk), .Q(reg_file[2037])
         );
  DFFPOSX1 reg_file_reg_15__118_ ( .D(n23090), .CLK(clk), .Q(reg_file[2038])
         );
  DFFPOSX1 reg_file_reg_15__119_ ( .D(n23089), .CLK(clk), .Q(reg_file[2039])
         );
  DFFPOSX1 reg_file_reg_15__120_ ( .D(n23088), .CLK(clk), .Q(reg_file[2040])
         );
  DFFPOSX1 reg_file_reg_15__121_ ( .D(n23087), .CLK(clk), .Q(reg_file[2041])
         );
  DFFPOSX1 reg_file_reg_15__122_ ( .D(n23086), .CLK(clk), .Q(reg_file[2042])
         );
  DFFPOSX1 reg_file_reg_15__123_ ( .D(n23085), .CLK(clk), .Q(reg_file[2043])
         );
  DFFPOSX1 reg_file_reg_15__124_ ( .D(n23084), .CLK(clk), .Q(reg_file[2044])
         );
  DFFPOSX1 reg_file_reg_15__125_ ( .D(n23083), .CLK(clk), .Q(reg_file[2045])
         );
  DFFPOSX1 reg_file_reg_15__126_ ( .D(n23082), .CLK(clk), .Q(reg_file[2046])
         );
  DFFPOSX1 reg_file_reg_15__127_ ( .D(n23081), .CLK(clk), .Q(reg_file[2047])
         );
  DFFPOSX1 reg_file_reg_16__0_ ( .D(n23080), .CLK(clk), .Q(reg_file[2048]) );
  DFFPOSX1 reg_file_reg_16__1_ ( .D(n23079), .CLK(clk), .Q(reg_file[2049]) );
  DFFPOSX1 reg_file_reg_16__2_ ( .D(n23078), .CLK(clk), .Q(reg_file[2050]) );
  DFFPOSX1 reg_file_reg_16__3_ ( .D(n23077), .CLK(clk), .Q(reg_file[2051]) );
  DFFPOSX1 reg_file_reg_16__4_ ( .D(n23076), .CLK(clk), .Q(reg_file[2052]) );
  DFFPOSX1 reg_file_reg_16__5_ ( .D(n23075), .CLK(clk), .Q(reg_file[2053]) );
  DFFPOSX1 reg_file_reg_16__6_ ( .D(n23074), .CLK(clk), .Q(reg_file[2054]) );
  DFFPOSX1 reg_file_reg_16__7_ ( .D(n23073), .CLK(clk), .Q(reg_file[2055]) );
  DFFPOSX1 reg_file_reg_16__8_ ( .D(n23072), .CLK(clk), .Q(reg_file[2056]) );
  DFFPOSX1 reg_file_reg_16__9_ ( .D(n23071), .CLK(clk), .Q(reg_file[2057]) );
  DFFPOSX1 reg_file_reg_16__10_ ( .D(n23070), .CLK(clk), .Q(reg_file[2058]) );
  DFFPOSX1 reg_file_reg_16__11_ ( .D(n23069), .CLK(clk), .Q(reg_file[2059]) );
  DFFPOSX1 reg_file_reg_16__12_ ( .D(n23068), .CLK(clk), .Q(reg_file[2060]) );
  DFFPOSX1 reg_file_reg_16__13_ ( .D(n23067), .CLK(clk), .Q(reg_file[2061]) );
  DFFPOSX1 reg_file_reg_16__14_ ( .D(n23066), .CLK(clk), .Q(reg_file[2062]) );
  DFFPOSX1 reg_file_reg_16__15_ ( .D(n23065), .CLK(clk), .Q(reg_file[2063]) );
  DFFPOSX1 reg_file_reg_16__16_ ( .D(n23064), .CLK(clk), .Q(reg_file[2064]) );
  DFFPOSX1 reg_file_reg_16__17_ ( .D(n23063), .CLK(clk), .Q(reg_file[2065]) );
  DFFPOSX1 reg_file_reg_16__18_ ( .D(n23062), .CLK(clk), .Q(reg_file[2066]) );
  DFFPOSX1 reg_file_reg_16__19_ ( .D(n23061), .CLK(clk), .Q(reg_file[2067]) );
  DFFPOSX1 reg_file_reg_16__20_ ( .D(n23060), .CLK(clk), .Q(reg_file[2068]) );
  DFFPOSX1 reg_file_reg_16__21_ ( .D(n23059), .CLK(clk), .Q(reg_file[2069]) );
  DFFPOSX1 reg_file_reg_16__22_ ( .D(n23058), .CLK(clk), .Q(reg_file[2070]) );
  DFFPOSX1 reg_file_reg_16__23_ ( .D(n23057), .CLK(clk), .Q(reg_file[2071]) );
  DFFPOSX1 reg_file_reg_16__24_ ( .D(n23056), .CLK(clk), .Q(reg_file[2072]) );
  DFFPOSX1 reg_file_reg_16__25_ ( .D(n23055), .CLK(clk), .Q(reg_file[2073]) );
  DFFPOSX1 reg_file_reg_16__26_ ( .D(n23054), .CLK(clk), .Q(reg_file[2074]) );
  DFFPOSX1 reg_file_reg_16__27_ ( .D(n23053), .CLK(clk), .Q(reg_file[2075]) );
  DFFPOSX1 reg_file_reg_16__28_ ( .D(n23052), .CLK(clk), .Q(reg_file[2076]) );
  DFFPOSX1 reg_file_reg_16__29_ ( .D(n23051), .CLK(clk), .Q(reg_file[2077]) );
  DFFPOSX1 reg_file_reg_16__30_ ( .D(n23050), .CLK(clk), .Q(reg_file[2078]) );
  DFFPOSX1 reg_file_reg_16__31_ ( .D(n23049), .CLK(clk), .Q(reg_file[2079]) );
  DFFPOSX1 reg_file_reg_16__32_ ( .D(n23048), .CLK(clk), .Q(reg_file[2080]) );
  DFFPOSX1 reg_file_reg_16__33_ ( .D(n23047), .CLK(clk), .Q(reg_file[2081]) );
  DFFPOSX1 reg_file_reg_16__34_ ( .D(n23046), .CLK(clk), .Q(reg_file[2082]) );
  DFFPOSX1 reg_file_reg_16__35_ ( .D(n23045), .CLK(clk), .Q(reg_file[2083]) );
  DFFPOSX1 reg_file_reg_16__36_ ( .D(n23044), .CLK(clk), .Q(reg_file[2084]) );
  DFFPOSX1 reg_file_reg_16__37_ ( .D(n23043), .CLK(clk), .Q(reg_file[2085]) );
  DFFPOSX1 reg_file_reg_16__38_ ( .D(n23042), .CLK(clk), .Q(reg_file[2086]) );
  DFFPOSX1 reg_file_reg_16__39_ ( .D(n23041), .CLK(clk), .Q(reg_file[2087]) );
  DFFPOSX1 reg_file_reg_16__40_ ( .D(n23040), .CLK(clk), .Q(reg_file[2088]) );
  DFFPOSX1 reg_file_reg_16__41_ ( .D(n23039), .CLK(clk), .Q(reg_file[2089]) );
  DFFPOSX1 reg_file_reg_16__42_ ( .D(n23038), .CLK(clk), .Q(reg_file[2090]) );
  DFFPOSX1 reg_file_reg_16__43_ ( .D(n23037), .CLK(clk), .Q(reg_file[2091]) );
  DFFPOSX1 reg_file_reg_16__44_ ( .D(n23036), .CLK(clk), .Q(reg_file[2092]) );
  DFFPOSX1 reg_file_reg_16__45_ ( .D(n23035), .CLK(clk), .Q(reg_file[2093]) );
  DFFPOSX1 reg_file_reg_16__46_ ( .D(n23034), .CLK(clk), .Q(reg_file[2094]) );
  DFFPOSX1 reg_file_reg_16__47_ ( .D(n23033), .CLK(clk), .Q(reg_file[2095]) );
  DFFPOSX1 reg_file_reg_16__48_ ( .D(n23032), .CLK(clk), .Q(reg_file[2096]) );
  DFFPOSX1 reg_file_reg_16__49_ ( .D(n23031), .CLK(clk), .Q(reg_file[2097]) );
  DFFPOSX1 reg_file_reg_16__50_ ( .D(n23030), .CLK(clk), .Q(reg_file[2098]) );
  DFFPOSX1 reg_file_reg_16__51_ ( .D(n23029), .CLK(clk), .Q(reg_file[2099]) );
  DFFPOSX1 reg_file_reg_16__52_ ( .D(n23028), .CLK(clk), .Q(reg_file[2100]) );
  DFFPOSX1 reg_file_reg_16__53_ ( .D(n23027), .CLK(clk), .Q(reg_file[2101]) );
  DFFPOSX1 reg_file_reg_16__54_ ( .D(n23026), .CLK(clk), .Q(reg_file[2102]) );
  DFFPOSX1 reg_file_reg_16__55_ ( .D(n23025), .CLK(clk), .Q(reg_file[2103]) );
  DFFPOSX1 reg_file_reg_16__56_ ( .D(n23024), .CLK(clk), .Q(reg_file[2104]) );
  DFFPOSX1 reg_file_reg_16__57_ ( .D(n23023), .CLK(clk), .Q(reg_file[2105]) );
  DFFPOSX1 reg_file_reg_16__58_ ( .D(n23022), .CLK(clk), .Q(reg_file[2106]) );
  DFFPOSX1 reg_file_reg_16__59_ ( .D(n23021), .CLK(clk), .Q(reg_file[2107]) );
  DFFPOSX1 reg_file_reg_16__60_ ( .D(n23020), .CLK(clk), .Q(reg_file[2108]) );
  DFFPOSX1 reg_file_reg_16__61_ ( .D(n23019), .CLK(clk), .Q(reg_file[2109]) );
  DFFPOSX1 reg_file_reg_16__62_ ( .D(n23018), .CLK(clk), .Q(reg_file[2110]) );
  DFFPOSX1 reg_file_reg_16__63_ ( .D(n23017), .CLK(clk), .Q(reg_file[2111]) );
  DFFPOSX1 reg_file_reg_16__64_ ( .D(n23016), .CLK(clk), .Q(reg_file[2112]) );
  DFFPOSX1 reg_file_reg_16__65_ ( .D(n23015), .CLK(clk), .Q(reg_file[2113]) );
  DFFPOSX1 reg_file_reg_16__66_ ( .D(n23014), .CLK(clk), .Q(reg_file[2114]) );
  DFFPOSX1 reg_file_reg_16__67_ ( .D(n23013), .CLK(clk), .Q(reg_file[2115]) );
  DFFPOSX1 reg_file_reg_16__68_ ( .D(n23012), .CLK(clk), .Q(reg_file[2116]) );
  DFFPOSX1 reg_file_reg_16__69_ ( .D(n23011), .CLK(clk), .Q(reg_file[2117]) );
  DFFPOSX1 reg_file_reg_16__70_ ( .D(n23010), .CLK(clk), .Q(reg_file[2118]) );
  DFFPOSX1 reg_file_reg_16__71_ ( .D(n23009), .CLK(clk), .Q(reg_file[2119]) );
  DFFPOSX1 reg_file_reg_16__72_ ( .D(n23008), .CLK(clk), .Q(reg_file[2120]) );
  DFFPOSX1 reg_file_reg_16__73_ ( .D(n23007), .CLK(clk), .Q(reg_file[2121]) );
  DFFPOSX1 reg_file_reg_16__74_ ( .D(n23006), .CLK(clk), .Q(reg_file[2122]) );
  DFFPOSX1 reg_file_reg_16__75_ ( .D(n23005), .CLK(clk), .Q(reg_file[2123]) );
  DFFPOSX1 reg_file_reg_16__76_ ( .D(n23004), .CLK(clk), .Q(reg_file[2124]) );
  DFFPOSX1 reg_file_reg_16__77_ ( .D(n23003), .CLK(clk), .Q(reg_file[2125]) );
  DFFPOSX1 reg_file_reg_16__78_ ( .D(n23002), .CLK(clk), .Q(reg_file[2126]) );
  DFFPOSX1 reg_file_reg_16__79_ ( .D(n23001), .CLK(clk), .Q(reg_file[2127]) );
  DFFPOSX1 reg_file_reg_16__80_ ( .D(n23000), .CLK(clk), .Q(reg_file[2128]) );
  DFFPOSX1 reg_file_reg_16__81_ ( .D(n22999), .CLK(clk), .Q(reg_file[2129]) );
  DFFPOSX1 reg_file_reg_16__82_ ( .D(n22998), .CLK(clk), .Q(reg_file[2130]) );
  DFFPOSX1 reg_file_reg_16__83_ ( .D(n22997), .CLK(clk), .Q(reg_file[2131]) );
  DFFPOSX1 reg_file_reg_16__84_ ( .D(n22996), .CLK(clk), .Q(reg_file[2132]) );
  DFFPOSX1 reg_file_reg_16__85_ ( .D(n22995), .CLK(clk), .Q(reg_file[2133]) );
  DFFPOSX1 reg_file_reg_16__86_ ( .D(n22994), .CLK(clk), .Q(reg_file[2134]) );
  DFFPOSX1 reg_file_reg_16__87_ ( .D(n22993), .CLK(clk), .Q(reg_file[2135]) );
  DFFPOSX1 reg_file_reg_16__88_ ( .D(n22992), .CLK(clk), .Q(reg_file[2136]) );
  DFFPOSX1 reg_file_reg_16__89_ ( .D(n22991), .CLK(clk), .Q(reg_file[2137]) );
  DFFPOSX1 reg_file_reg_16__90_ ( .D(n22990), .CLK(clk), .Q(reg_file[2138]) );
  DFFPOSX1 reg_file_reg_16__91_ ( .D(n22989), .CLK(clk), .Q(reg_file[2139]) );
  DFFPOSX1 reg_file_reg_16__92_ ( .D(n22988), .CLK(clk), .Q(reg_file[2140]) );
  DFFPOSX1 reg_file_reg_16__93_ ( .D(n22987), .CLK(clk), .Q(reg_file[2141]) );
  DFFPOSX1 reg_file_reg_16__94_ ( .D(n22986), .CLK(clk), .Q(reg_file[2142]) );
  DFFPOSX1 reg_file_reg_16__95_ ( .D(n22985), .CLK(clk), .Q(reg_file[2143]) );
  DFFPOSX1 reg_file_reg_16__96_ ( .D(n22984), .CLK(clk), .Q(reg_file[2144]) );
  DFFPOSX1 reg_file_reg_16__97_ ( .D(n22983), .CLK(clk), .Q(reg_file[2145]) );
  DFFPOSX1 reg_file_reg_16__98_ ( .D(n22982), .CLK(clk), .Q(reg_file[2146]) );
  DFFPOSX1 reg_file_reg_16__99_ ( .D(n22981), .CLK(clk), .Q(reg_file[2147]) );
  DFFPOSX1 reg_file_reg_16__100_ ( .D(n22980), .CLK(clk), .Q(reg_file[2148])
         );
  DFFPOSX1 reg_file_reg_16__101_ ( .D(n22979), .CLK(clk), .Q(reg_file[2149])
         );
  DFFPOSX1 reg_file_reg_16__102_ ( .D(n22978), .CLK(clk), .Q(reg_file[2150])
         );
  DFFPOSX1 reg_file_reg_16__103_ ( .D(n22977), .CLK(clk), .Q(reg_file[2151])
         );
  DFFPOSX1 reg_file_reg_16__104_ ( .D(n22976), .CLK(clk), .Q(reg_file[2152])
         );
  DFFPOSX1 reg_file_reg_16__105_ ( .D(n22975), .CLK(clk), .Q(reg_file[2153])
         );
  DFFPOSX1 reg_file_reg_16__106_ ( .D(n22974), .CLK(clk), .Q(reg_file[2154])
         );
  DFFPOSX1 reg_file_reg_16__107_ ( .D(n22973), .CLK(clk), .Q(reg_file[2155])
         );
  DFFPOSX1 reg_file_reg_16__108_ ( .D(n22972), .CLK(clk), .Q(reg_file[2156])
         );
  DFFPOSX1 reg_file_reg_16__109_ ( .D(n22971), .CLK(clk), .Q(reg_file[2157])
         );
  DFFPOSX1 reg_file_reg_16__110_ ( .D(n22970), .CLK(clk), .Q(reg_file[2158])
         );
  DFFPOSX1 reg_file_reg_16__111_ ( .D(n22969), .CLK(clk), .Q(reg_file[2159])
         );
  DFFPOSX1 reg_file_reg_16__112_ ( .D(n22968), .CLK(clk), .Q(reg_file[2160])
         );
  DFFPOSX1 reg_file_reg_16__113_ ( .D(n22967), .CLK(clk), .Q(reg_file[2161])
         );
  DFFPOSX1 reg_file_reg_16__114_ ( .D(n22966), .CLK(clk), .Q(reg_file[2162])
         );
  DFFPOSX1 reg_file_reg_16__115_ ( .D(n22965), .CLK(clk), .Q(reg_file[2163])
         );
  DFFPOSX1 reg_file_reg_16__116_ ( .D(n22964), .CLK(clk), .Q(reg_file[2164])
         );
  DFFPOSX1 reg_file_reg_16__117_ ( .D(n22963), .CLK(clk), .Q(reg_file[2165])
         );
  DFFPOSX1 reg_file_reg_16__118_ ( .D(n22962), .CLK(clk), .Q(reg_file[2166])
         );
  DFFPOSX1 reg_file_reg_16__119_ ( .D(n22961), .CLK(clk), .Q(reg_file[2167])
         );
  DFFPOSX1 reg_file_reg_16__120_ ( .D(n22960), .CLK(clk), .Q(reg_file[2168])
         );
  DFFPOSX1 reg_file_reg_16__121_ ( .D(n22959), .CLK(clk), .Q(reg_file[2169])
         );
  DFFPOSX1 reg_file_reg_16__122_ ( .D(n22958), .CLK(clk), .Q(reg_file[2170])
         );
  DFFPOSX1 reg_file_reg_16__123_ ( .D(n22957), .CLK(clk), .Q(reg_file[2171])
         );
  DFFPOSX1 reg_file_reg_16__124_ ( .D(n22956), .CLK(clk), .Q(reg_file[2172])
         );
  DFFPOSX1 reg_file_reg_16__125_ ( .D(n22955), .CLK(clk), .Q(reg_file[2173])
         );
  DFFPOSX1 reg_file_reg_16__126_ ( .D(n22954), .CLK(clk), .Q(reg_file[2174])
         );
  DFFPOSX1 reg_file_reg_16__127_ ( .D(n22953), .CLK(clk), .Q(reg_file[2175])
         );
  DFFPOSX1 reg_file_reg_17__0_ ( .D(n22952), .CLK(clk), .Q(reg_file[2176]) );
  DFFPOSX1 reg_file_reg_17__1_ ( .D(n22951), .CLK(clk), .Q(reg_file[2177]) );
  DFFPOSX1 reg_file_reg_17__2_ ( .D(n22950), .CLK(clk), .Q(reg_file[2178]) );
  DFFPOSX1 reg_file_reg_17__3_ ( .D(n22949), .CLK(clk), .Q(reg_file[2179]) );
  DFFPOSX1 reg_file_reg_17__4_ ( .D(n22948), .CLK(clk), .Q(reg_file[2180]) );
  DFFPOSX1 reg_file_reg_17__5_ ( .D(n22947), .CLK(clk), .Q(reg_file[2181]) );
  DFFPOSX1 reg_file_reg_17__6_ ( .D(n22946), .CLK(clk), .Q(reg_file[2182]) );
  DFFPOSX1 reg_file_reg_17__7_ ( .D(n22945), .CLK(clk), .Q(reg_file[2183]) );
  DFFPOSX1 reg_file_reg_17__8_ ( .D(n22944), .CLK(clk), .Q(reg_file[2184]) );
  DFFPOSX1 reg_file_reg_17__9_ ( .D(n22943), .CLK(clk), .Q(reg_file[2185]) );
  DFFPOSX1 reg_file_reg_17__10_ ( .D(n22942), .CLK(clk), .Q(reg_file[2186]) );
  DFFPOSX1 reg_file_reg_17__11_ ( .D(n22941), .CLK(clk), .Q(reg_file[2187]) );
  DFFPOSX1 reg_file_reg_17__12_ ( .D(n22940), .CLK(clk), .Q(reg_file[2188]) );
  DFFPOSX1 reg_file_reg_17__13_ ( .D(n22939), .CLK(clk), .Q(reg_file[2189]) );
  DFFPOSX1 reg_file_reg_17__14_ ( .D(n22938), .CLK(clk), .Q(reg_file[2190]) );
  DFFPOSX1 reg_file_reg_17__15_ ( .D(n22937), .CLK(clk), .Q(reg_file[2191]) );
  DFFPOSX1 reg_file_reg_17__16_ ( .D(n22936), .CLK(clk), .Q(reg_file[2192]) );
  DFFPOSX1 reg_file_reg_17__17_ ( .D(n22935), .CLK(clk), .Q(reg_file[2193]) );
  DFFPOSX1 reg_file_reg_17__18_ ( .D(n22934), .CLK(clk), .Q(reg_file[2194]) );
  DFFPOSX1 reg_file_reg_17__19_ ( .D(n22933), .CLK(clk), .Q(reg_file[2195]) );
  DFFPOSX1 reg_file_reg_17__20_ ( .D(n22932), .CLK(clk), .Q(reg_file[2196]) );
  DFFPOSX1 reg_file_reg_17__21_ ( .D(n22931), .CLK(clk), .Q(reg_file[2197]) );
  DFFPOSX1 reg_file_reg_17__22_ ( .D(n22930), .CLK(clk), .Q(reg_file[2198]) );
  DFFPOSX1 reg_file_reg_17__23_ ( .D(n22929), .CLK(clk), .Q(reg_file[2199]) );
  DFFPOSX1 reg_file_reg_17__24_ ( .D(n22928), .CLK(clk), .Q(reg_file[2200]) );
  DFFPOSX1 reg_file_reg_17__25_ ( .D(n22927), .CLK(clk), .Q(reg_file[2201]) );
  DFFPOSX1 reg_file_reg_17__26_ ( .D(n22926), .CLK(clk), .Q(reg_file[2202]) );
  DFFPOSX1 reg_file_reg_17__27_ ( .D(n22925), .CLK(clk), .Q(reg_file[2203]) );
  DFFPOSX1 reg_file_reg_17__28_ ( .D(n22924), .CLK(clk), .Q(reg_file[2204]) );
  DFFPOSX1 reg_file_reg_17__29_ ( .D(n22923), .CLK(clk), .Q(reg_file[2205]) );
  DFFPOSX1 reg_file_reg_17__30_ ( .D(n22922), .CLK(clk), .Q(reg_file[2206]) );
  DFFPOSX1 reg_file_reg_17__31_ ( .D(n22921), .CLK(clk), .Q(reg_file[2207]) );
  DFFPOSX1 reg_file_reg_17__32_ ( .D(n22920), .CLK(clk), .Q(reg_file[2208]) );
  DFFPOSX1 reg_file_reg_17__33_ ( .D(n22919), .CLK(clk), .Q(reg_file[2209]) );
  DFFPOSX1 reg_file_reg_17__34_ ( .D(n22918), .CLK(clk), .Q(reg_file[2210]) );
  DFFPOSX1 reg_file_reg_17__35_ ( .D(n22917), .CLK(clk), .Q(reg_file[2211]) );
  DFFPOSX1 reg_file_reg_17__36_ ( .D(n22916), .CLK(clk), .Q(reg_file[2212]) );
  DFFPOSX1 reg_file_reg_17__37_ ( .D(n22915), .CLK(clk), .Q(reg_file[2213]) );
  DFFPOSX1 reg_file_reg_17__38_ ( .D(n22914), .CLK(clk), .Q(reg_file[2214]) );
  DFFPOSX1 reg_file_reg_17__39_ ( .D(n22913), .CLK(clk), .Q(reg_file[2215]) );
  DFFPOSX1 reg_file_reg_17__40_ ( .D(n22912), .CLK(clk), .Q(reg_file[2216]) );
  DFFPOSX1 reg_file_reg_17__41_ ( .D(n22911), .CLK(clk), .Q(reg_file[2217]) );
  DFFPOSX1 reg_file_reg_17__42_ ( .D(n22910), .CLK(clk), .Q(reg_file[2218]) );
  DFFPOSX1 reg_file_reg_17__43_ ( .D(n22909), .CLK(clk), .Q(reg_file[2219]) );
  DFFPOSX1 reg_file_reg_17__44_ ( .D(n22908), .CLK(clk), .Q(reg_file[2220]) );
  DFFPOSX1 reg_file_reg_17__45_ ( .D(n22907), .CLK(clk), .Q(reg_file[2221]) );
  DFFPOSX1 reg_file_reg_17__46_ ( .D(n22906), .CLK(clk), .Q(reg_file[2222]) );
  DFFPOSX1 reg_file_reg_17__47_ ( .D(n22905), .CLK(clk), .Q(reg_file[2223]) );
  DFFPOSX1 reg_file_reg_17__48_ ( .D(n22904), .CLK(clk), .Q(reg_file[2224]) );
  DFFPOSX1 reg_file_reg_17__49_ ( .D(n22903), .CLK(clk), .Q(reg_file[2225]) );
  DFFPOSX1 reg_file_reg_17__50_ ( .D(n22902), .CLK(clk), .Q(reg_file[2226]) );
  DFFPOSX1 reg_file_reg_17__51_ ( .D(n22901), .CLK(clk), .Q(reg_file[2227]) );
  DFFPOSX1 reg_file_reg_17__52_ ( .D(n22900), .CLK(clk), .Q(reg_file[2228]) );
  DFFPOSX1 reg_file_reg_17__53_ ( .D(n22899), .CLK(clk), .Q(reg_file[2229]) );
  DFFPOSX1 reg_file_reg_17__54_ ( .D(n22898), .CLK(clk), .Q(reg_file[2230]) );
  DFFPOSX1 reg_file_reg_17__55_ ( .D(n22897), .CLK(clk), .Q(reg_file[2231]) );
  DFFPOSX1 reg_file_reg_17__56_ ( .D(n22896), .CLK(clk), .Q(reg_file[2232]) );
  DFFPOSX1 reg_file_reg_17__57_ ( .D(n22895), .CLK(clk), .Q(reg_file[2233]) );
  DFFPOSX1 reg_file_reg_17__58_ ( .D(n22894), .CLK(clk), .Q(reg_file[2234]) );
  DFFPOSX1 reg_file_reg_17__59_ ( .D(n22893), .CLK(clk), .Q(reg_file[2235]) );
  DFFPOSX1 reg_file_reg_17__60_ ( .D(n22892), .CLK(clk), .Q(reg_file[2236]) );
  DFFPOSX1 reg_file_reg_17__61_ ( .D(n22891), .CLK(clk), .Q(reg_file[2237]) );
  DFFPOSX1 reg_file_reg_17__62_ ( .D(n22890), .CLK(clk), .Q(reg_file[2238]) );
  DFFPOSX1 reg_file_reg_17__63_ ( .D(n22889), .CLK(clk), .Q(reg_file[2239]) );
  DFFPOSX1 reg_file_reg_17__64_ ( .D(n22888), .CLK(clk), .Q(reg_file[2240]) );
  DFFPOSX1 reg_file_reg_17__65_ ( .D(n22887), .CLK(clk), .Q(reg_file[2241]) );
  DFFPOSX1 reg_file_reg_17__66_ ( .D(n22886), .CLK(clk), .Q(reg_file[2242]) );
  DFFPOSX1 reg_file_reg_17__67_ ( .D(n22885), .CLK(clk), .Q(reg_file[2243]) );
  DFFPOSX1 reg_file_reg_17__68_ ( .D(n22884), .CLK(clk), .Q(reg_file[2244]) );
  DFFPOSX1 reg_file_reg_17__69_ ( .D(n22883), .CLK(clk), .Q(reg_file[2245]) );
  DFFPOSX1 reg_file_reg_17__70_ ( .D(n22882), .CLK(clk), .Q(reg_file[2246]) );
  DFFPOSX1 reg_file_reg_17__71_ ( .D(n22881), .CLK(clk), .Q(reg_file[2247]) );
  DFFPOSX1 reg_file_reg_17__72_ ( .D(n22880), .CLK(clk), .Q(reg_file[2248]) );
  DFFPOSX1 reg_file_reg_17__73_ ( .D(n22879), .CLK(clk), .Q(reg_file[2249]) );
  DFFPOSX1 reg_file_reg_17__74_ ( .D(n22878), .CLK(clk), .Q(reg_file[2250]) );
  DFFPOSX1 reg_file_reg_17__75_ ( .D(n22877), .CLK(clk), .Q(reg_file[2251]) );
  DFFPOSX1 reg_file_reg_17__76_ ( .D(n22876), .CLK(clk), .Q(reg_file[2252]) );
  DFFPOSX1 reg_file_reg_17__77_ ( .D(n22875), .CLK(clk), .Q(reg_file[2253]) );
  DFFPOSX1 reg_file_reg_17__78_ ( .D(n22874), .CLK(clk), .Q(reg_file[2254]) );
  DFFPOSX1 reg_file_reg_17__79_ ( .D(n22873), .CLK(clk), .Q(reg_file[2255]) );
  DFFPOSX1 reg_file_reg_17__80_ ( .D(n22872), .CLK(clk), .Q(reg_file[2256]) );
  DFFPOSX1 reg_file_reg_17__81_ ( .D(n22871), .CLK(clk), .Q(reg_file[2257]) );
  DFFPOSX1 reg_file_reg_17__82_ ( .D(n22870), .CLK(clk), .Q(reg_file[2258]) );
  DFFPOSX1 reg_file_reg_17__83_ ( .D(n22869), .CLK(clk), .Q(reg_file[2259]) );
  DFFPOSX1 reg_file_reg_17__84_ ( .D(n22868), .CLK(clk), .Q(reg_file[2260]) );
  DFFPOSX1 reg_file_reg_17__85_ ( .D(n22867), .CLK(clk), .Q(reg_file[2261]) );
  DFFPOSX1 reg_file_reg_17__86_ ( .D(n22866), .CLK(clk), .Q(reg_file[2262]) );
  DFFPOSX1 reg_file_reg_17__87_ ( .D(n22865), .CLK(clk), .Q(reg_file[2263]) );
  DFFPOSX1 reg_file_reg_17__88_ ( .D(n22864), .CLK(clk), .Q(reg_file[2264]) );
  DFFPOSX1 reg_file_reg_17__89_ ( .D(n22863), .CLK(clk), .Q(reg_file[2265]) );
  DFFPOSX1 reg_file_reg_17__90_ ( .D(n22862), .CLK(clk), .Q(reg_file[2266]) );
  DFFPOSX1 reg_file_reg_17__91_ ( .D(n22861), .CLK(clk), .Q(reg_file[2267]) );
  DFFPOSX1 reg_file_reg_17__92_ ( .D(n22860), .CLK(clk), .Q(reg_file[2268]) );
  DFFPOSX1 reg_file_reg_17__93_ ( .D(n22859), .CLK(clk), .Q(reg_file[2269]) );
  DFFPOSX1 reg_file_reg_17__94_ ( .D(n22858), .CLK(clk), .Q(reg_file[2270]) );
  DFFPOSX1 reg_file_reg_17__95_ ( .D(n22857), .CLK(clk), .Q(reg_file[2271]) );
  DFFPOSX1 reg_file_reg_17__96_ ( .D(n22856), .CLK(clk), .Q(reg_file[2272]) );
  DFFPOSX1 reg_file_reg_17__97_ ( .D(n22855), .CLK(clk), .Q(reg_file[2273]) );
  DFFPOSX1 reg_file_reg_17__98_ ( .D(n22854), .CLK(clk), .Q(reg_file[2274]) );
  DFFPOSX1 reg_file_reg_17__99_ ( .D(n22853), .CLK(clk), .Q(reg_file[2275]) );
  DFFPOSX1 reg_file_reg_17__100_ ( .D(n22852), .CLK(clk), .Q(reg_file[2276])
         );
  DFFPOSX1 reg_file_reg_17__101_ ( .D(n22851), .CLK(clk), .Q(reg_file[2277])
         );
  DFFPOSX1 reg_file_reg_17__102_ ( .D(n22850), .CLK(clk), .Q(reg_file[2278])
         );
  DFFPOSX1 reg_file_reg_17__103_ ( .D(n22849), .CLK(clk), .Q(reg_file[2279])
         );
  DFFPOSX1 reg_file_reg_17__104_ ( .D(n22848), .CLK(clk), .Q(reg_file[2280])
         );
  DFFPOSX1 reg_file_reg_17__105_ ( .D(n22847), .CLK(clk), .Q(reg_file[2281])
         );
  DFFPOSX1 reg_file_reg_17__106_ ( .D(n22846), .CLK(clk), .Q(reg_file[2282])
         );
  DFFPOSX1 reg_file_reg_17__107_ ( .D(n22845), .CLK(clk), .Q(reg_file[2283])
         );
  DFFPOSX1 reg_file_reg_17__108_ ( .D(n22844), .CLK(clk), .Q(reg_file[2284])
         );
  DFFPOSX1 reg_file_reg_17__109_ ( .D(n22843), .CLK(clk), .Q(reg_file[2285])
         );
  DFFPOSX1 reg_file_reg_17__110_ ( .D(n22842), .CLK(clk), .Q(reg_file[2286])
         );
  DFFPOSX1 reg_file_reg_17__111_ ( .D(n22841), .CLK(clk), .Q(reg_file[2287])
         );
  DFFPOSX1 reg_file_reg_17__112_ ( .D(n22840), .CLK(clk), .Q(reg_file[2288])
         );
  DFFPOSX1 reg_file_reg_17__113_ ( .D(n22839), .CLK(clk), .Q(reg_file[2289])
         );
  DFFPOSX1 reg_file_reg_17__114_ ( .D(n22838), .CLK(clk), .Q(reg_file[2290])
         );
  DFFPOSX1 reg_file_reg_17__115_ ( .D(n22837), .CLK(clk), .Q(reg_file[2291])
         );
  DFFPOSX1 reg_file_reg_17__116_ ( .D(n22836), .CLK(clk), .Q(reg_file[2292])
         );
  DFFPOSX1 reg_file_reg_17__117_ ( .D(n22835), .CLK(clk), .Q(reg_file[2293])
         );
  DFFPOSX1 reg_file_reg_17__118_ ( .D(n22834), .CLK(clk), .Q(reg_file[2294])
         );
  DFFPOSX1 reg_file_reg_17__119_ ( .D(n22833), .CLK(clk), .Q(reg_file[2295])
         );
  DFFPOSX1 reg_file_reg_17__120_ ( .D(n22832), .CLK(clk), .Q(reg_file[2296])
         );
  DFFPOSX1 reg_file_reg_17__121_ ( .D(n22831), .CLK(clk), .Q(reg_file[2297])
         );
  DFFPOSX1 reg_file_reg_17__122_ ( .D(n22830), .CLK(clk), .Q(reg_file[2298])
         );
  DFFPOSX1 reg_file_reg_17__123_ ( .D(n22829), .CLK(clk), .Q(reg_file[2299])
         );
  DFFPOSX1 reg_file_reg_17__124_ ( .D(n22828), .CLK(clk), .Q(reg_file[2300])
         );
  DFFPOSX1 reg_file_reg_17__125_ ( .D(n22827), .CLK(clk), .Q(reg_file[2301])
         );
  DFFPOSX1 reg_file_reg_17__126_ ( .D(n22826), .CLK(clk), .Q(reg_file[2302])
         );
  DFFPOSX1 reg_file_reg_17__127_ ( .D(n22825), .CLK(clk), .Q(reg_file[2303])
         );
  DFFPOSX1 reg_file_reg_18__0_ ( .D(n22824), .CLK(clk), .Q(reg_file[2304]) );
  DFFPOSX1 reg_file_reg_18__1_ ( .D(n22823), .CLK(clk), .Q(reg_file[2305]) );
  DFFPOSX1 reg_file_reg_18__2_ ( .D(n22822), .CLK(clk), .Q(reg_file[2306]) );
  DFFPOSX1 reg_file_reg_18__3_ ( .D(n22821), .CLK(clk), .Q(reg_file[2307]) );
  DFFPOSX1 reg_file_reg_18__4_ ( .D(n22820), .CLK(clk), .Q(reg_file[2308]) );
  DFFPOSX1 reg_file_reg_18__5_ ( .D(n22819), .CLK(clk), .Q(reg_file[2309]) );
  DFFPOSX1 reg_file_reg_18__6_ ( .D(n22818), .CLK(clk), .Q(reg_file[2310]) );
  DFFPOSX1 reg_file_reg_18__7_ ( .D(n22817), .CLK(clk), .Q(reg_file[2311]) );
  DFFPOSX1 reg_file_reg_18__8_ ( .D(n22816), .CLK(clk), .Q(reg_file[2312]) );
  DFFPOSX1 reg_file_reg_18__9_ ( .D(n22815), .CLK(clk), .Q(reg_file[2313]) );
  DFFPOSX1 reg_file_reg_18__10_ ( .D(n22814), .CLK(clk), .Q(reg_file[2314]) );
  DFFPOSX1 reg_file_reg_18__11_ ( .D(n22813), .CLK(clk), .Q(reg_file[2315]) );
  DFFPOSX1 reg_file_reg_18__12_ ( .D(n22812), .CLK(clk), .Q(reg_file[2316]) );
  DFFPOSX1 reg_file_reg_18__13_ ( .D(n22811), .CLK(clk), .Q(reg_file[2317]) );
  DFFPOSX1 reg_file_reg_18__14_ ( .D(n22810), .CLK(clk), .Q(reg_file[2318]) );
  DFFPOSX1 reg_file_reg_18__15_ ( .D(n22809), .CLK(clk), .Q(reg_file[2319]) );
  DFFPOSX1 reg_file_reg_18__16_ ( .D(n22808), .CLK(clk), .Q(reg_file[2320]) );
  DFFPOSX1 reg_file_reg_18__17_ ( .D(n22807), .CLK(clk), .Q(reg_file[2321]) );
  DFFPOSX1 reg_file_reg_18__18_ ( .D(n22806), .CLK(clk), .Q(reg_file[2322]) );
  DFFPOSX1 reg_file_reg_18__19_ ( .D(n22805), .CLK(clk), .Q(reg_file[2323]) );
  DFFPOSX1 reg_file_reg_18__20_ ( .D(n22804), .CLK(clk), .Q(reg_file[2324]) );
  DFFPOSX1 reg_file_reg_18__21_ ( .D(n22803), .CLK(clk), .Q(reg_file[2325]) );
  DFFPOSX1 reg_file_reg_18__22_ ( .D(n22802), .CLK(clk), .Q(reg_file[2326]) );
  DFFPOSX1 reg_file_reg_18__23_ ( .D(n22801), .CLK(clk), .Q(reg_file[2327]) );
  DFFPOSX1 reg_file_reg_18__24_ ( .D(n22800), .CLK(clk), .Q(reg_file[2328]) );
  DFFPOSX1 reg_file_reg_18__25_ ( .D(n22799), .CLK(clk), .Q(reg_file[2329]) );
  DFFPOSX1 reg_file_reg_18__26_ ( .D(n22798), .CLK(clk), .Q(reg_file[2330]) );
  DFFPOSX1 reg_file_reg_18__27_ ( .D(n22797), .CLK(clk), .Q(reg_file[2331]) );
  DFFPOSX1 reg_file_reg_18__28_ ( .D(n22796), .CLK(clk), .Q(reg_file[2332]) );
  DFFPOSX1 reg_file_reg_18__29_ ( .D(n22795), .CLK(clk), .Q(reg_file[2333]) );
  DFFPOSX1 reg_file_reg_18__30_ ( .D(n22794), .CLK(clk), .Q(reg_file[2334]) );
  DFFPOSX1 reg_file_reg_18__31_ ( .D(n22793), .CLK(clk), .Q(reg_file[2335]) );
  DFFPOSX1 reg_file_reg_18__32_ ( .D(n22792), .CLK(clk), .Q(reg_file[2336]) );
  DFFPOSX1 reg_file_reg_18__33_ ( .D(n22791), .CLK(clk), .Q(reg_file[2337]) );
  DFFPOSX1 reg_file_reg_18__34_ ( .D(n22790), .CLK(clk), .Q(reg_file[2338]) );
  DFFPOSX1 reg_file_reg_18__35_ ( .D(n22789), .CLK(clk), .Q(reg_file[2339]) );
  DFFPOSX1 reg_file_reg_18__36_ ( .D(n22788), .CLK(clk), .Q(reg_file[2340]) );
  DFFPOSX1 reg_file_reg_18__37_ ( .D(n22787), .CLK(clk), .Q(reg_file[2341]) );
  DFFPOSX1 reg_file_reg_18__38_ ( .D(n22786), .CLK(clk), .Q(reg_file[2342]) );
  DFFPOSX1 reg_file_reg_18__39_ ( .D(n22785), .CLK(clk), .Q(reg_file[2343]) );
  DFFPOSX1 reg_file_reg_18__40_ ( .D(n22784), .CLK(clk), .Q(reg_file[2344]) );
  DFFPOSX1 reg_file_reg_18__41_ ( .D(n22783), .CLK(clk), .Q(reg_file[2345]) );
  DFFPOSX1 reg_file_reg_18__42_ ( .D(n22782), .CLK(clk), .Q(reg_file[2346]) );
  DFFPOSX1 reg_file_reg_18__43_ ( .D(n22781), .CLK(clk), .Q(reg_file[2347]) );
  DFFPOSX1 reg_file_reg_18__44_ ( .D(n22780), .CLK(clk), .Q(reg_file[2348]) );
  DFFPOSX1 reg_file_reg_18__45_ ( .D(n22779), .CLK(clk), .Q(reg_file[2349]) );
  DFFPOSX1 reg_file_reg_18__46_ ( .D(n22778), .CLK(clk), .Q(reg_file[2350]) );
  DFFPOSX1 reg_file_reg_18__47_ ( .D(n22777), .CLK(clk), .Q(reg_file[2351]) );
  DFFPOSX1 reg_file_reg_18__48_ ( .D(n22776), .CLK(clk), .Q(reg_file[2352]) );
  DFFPOSX1 reg_file_reg_18__49_ ( .D(n22775), .CLK(clk), .Q(reg_file[2353]) );
  DFFPOSX1 reg_file_reg_18__50_ ( .D(n22774), .CLK(clk), .Q(reg_file[2354]) );
  DFFPOSX1 reg_file_reg_18__51_ ( .D(n22773), .CLK(clk), .Q(reg_file[2355]) );
  DFFPOSX1 reg_file_reg_18__52_ ( .D(n22772), .CLK(clk), .Q(reg_file[2356]) );
  DFFPOSX1 reg_file_reg_18__53_ ( .D(n22771), .CLK(clk), .Q(reg_file[2357]) );
  DFFPOSX1 reg_file_reg_18__54_ ( .D(n22770), .CLK(clk), .Q(reg_file[2358]) );
  DFFPOSX1 reg_file_reg_18__55_ ( .D(n22769), .CLK(clk), .Q(reg_file[2359]) );
  DFFPOSX1 reg_file_reg_18__56_ ( .D(n22768), .CLK(clk), .Q(reg_file[2360]) );
  DFFPOSX1 reg_file_reg_18__57_ ( .D(n22767), .CLK(clk), .Q(reg_file[2361]) );
  DFFPOSX1 reg_file_reg_18__58_ ( .D(n22766), .CLK(clk), .Q(reg_file[2362]) );
  DFFPOSX1 reg_file_reg_18__59_ ( .D(n22765), .CLK(clk), .Q(reg_file[2363]) );
  DFFPOSX1 reg_file_reg_18__60_ ( .D(n22764), .CLK(clk), .Q(reg_file[2364]) );
  DFFPOSX1 reg_file_reg_18__61_ ( .D(n22763), .CLK(clk), .Q(reg_file[2365]) );
  DFFPOSX1 reg_file_reg_18__62_ ( .D(n22762), .CLK(clk), .Q(reg_file[2366]) );
  DFFPOSX1 reg_file_reg_18__63_ ( .D(n22761), .CLK(clk), .Q(reg_file[2367]) );
  DFFPOSX1 reg_file_reg_18__64_ ( .D(n22760), .CLK(clk), .Q(reg_file[2368]) );
  DFFPOSX1 reg_file_reg_18__65_ ( .D(n22759), .CLK(clk), .Q(reg_file[2369]) );
  DFFPOSX1 reg_file_reg_18__66_ ( .D(n22758), .CLK(clk), .Q(reg_file[2370]) );
  DFFPOSX1 reg_file_reg_18__67_ ( .D(n22757), .CLK(clk), .Q(reg_file[2371]) );
  DFFPOSX1 reg_file_reg_18__68_ ( .D(n22756), .CLK(clk), .Q(reg_file[2372]) );
  DFFPOSX1 reg_file_reg_18__69_ ( .D(n22755), .CLK(clk), .Q(reg_file[2373]) );
  DFFPOSX1 reg_file_reg_18__70_ ( .D(n22754), .CLK(clk), .Q(reg_file[2374]) );
  DFFPOSX1 reg_file_reg_18__71_ ( .D(n22753), .CLK(clk), .Q(reg_file[2375]) );
  DFFPOSX1 reg_file_reg_18__72_ ( .D(n22752), .CLK(clk), .Q(reg_file[2376]) );
  DFFPOSX1 reg_file_reg_18__73_ ( .D(n22751), .CLK(clk), .Q(reg_file[2377]) );
  DFFPOSX1 reg_file_reg_18__74_ ( .D(n22750), .CLK(clk), .Q(reg_file[2378]) );
  DFFPOSX1 reg_file_reg_18__75_ ( .D(n22749), .CLK(clk), .Q(reg_file[2379]) );
  DFFPOSX1 reg_file_reg_18__76_ ( .D(n22748), .CLK(clk), .Q(reg_file[2380]) );
  DFFPOSX1 reg_file_reg_18__77_ ( .D(n22747), .CLK(clk), .Q(reg_file[2381]) );
  DFFPOSX1 reg_file_reg_18__78_ ( .D(n22746), .CLK(clk), .Q(reg_file[2382]) );
  DFFPOSX1 reg_file_reg_18__79_ ( .D(n22745), .CLK(clk), .Q(reg_file[2383]) );
  DFFPOSX1 reg_file_reg_18__80_ ( .D(n22744), .CLK(clk), .Q(reg_file[2384]) );
  DFFPOSX1 reg_file_reg_18__81_ ( .D(n22743), .CLK(clk), .Q(reg_file[2385]) );
  DFFPOSX1 reg_file_reg_18__82_ ( .D(n22742), .CLK(clk), .Q(reg_file[2386]) );
  DFFPOSX1 reg_file_reg_18__83_ ( .D(n22741), .CLK(clk), .Q(reg_file[2387]) );
  DFFPOSX1 reg_file_reg_18__84_ ( .D(n22740), .CLK(clk), .Q(reg_file[2388]) );
  DFFPOSX1 reg_file_reg_18__85_ ( .D(n22739), .CLK(clk), .Q(reg_file[2389]) );
  DFFPOSX1 reg_file_reg_18__86_ ( .D(n22738), .CLK(clk), .Q(reg_file[2390]) );
  DFFPOSX1 reg_file_reg_18__87_ ( .D(n22737), .CLK(clk), .Q(reg_file[2391]) );
  DFFPOSX1 reg_file_reg_18__88_ ( .D(n22736), .CLK(clk), .Q(reg_file[2392]) );
  DFFPOSX1 reg_file_reg_18__89_ ( .D(n22735), .CLK(clk), .Q(reg_file[2393]) );
  DFFPOSX1 reg_file_reg_18__90_ ( .D(n22734), .CLK(clk), .Q(reg_file[2394]) );
  DFFPOSX1 reg_file_reg_18__91_ ( .D(n22733), .CLK(clk), .Q(reg_file[2395]) );
  DFFPOSX1 reg_file_reg_18__92_ ( .D(n22732), .CLK(clk), .Q(reg_file[2396]) );
  DFFPOSX1 reg_file_reg_18__93_ ( .D(n22731), .CLK(clk), .Q(reg_file[2397]) );
  DFFPOSX1 reg_file_reg_18__94_ ( .D(n22730), .CLK(clk), .Q(reg_file[2398]) );
  DFFPOSX1 reg_file_reg_18__95_ ( .D(n22729), .CLK(clk), .Q(reg_file[2399]) );
  DFFPOSX1 reg_file_reg_18__96_ ( .D(n22728), .CLK(clk), .Q(reg_file[2400]) );
  DFFPOSX1 reg_file_reg_18__97_ ( .D(n22727), .CLK(clk), .Q(reg_file[2401]) );
  DFFPOSX1 reg_file_reg_18__98_ ( .D(n22726), .CLK(clk), .Q(reg_file[2402]) );
  DFFPOSX1 reg_file_reg_18__99_ ( .D(n22725), .CLK(clk), .Q(reg_file[2403]) );
  DFFPOSX1 reg_file_reg_18__100_ ( .D(n22724), .CLK(clk), .Q(reg_file[2404])
         );
  DFFPOSX1 reg_file_reg_18__101_ ( .D(n22723), .CLK(clk), .Q(reg_file[2405])
         );
  DFFPOSX1 reg_file_reg_18__102_ ( .D(n22722), .CLK(clk), .Q(reg_file[2406])
         );
  DFFPOSX1 reg_file_reg_18__103_ ( .D(n22721), .CLK(clk), .Q(reg_file[2407])
         );
  DFFPOSX1 reg_file_reg_18__104_ ( .D(n22720), .CLK(clk), .Q(reg_file[2408])
         );
  DFFPOSX1 reg_file_reg_18__105_ ( .D(n22719), .CLK(clk), .Q(reg_file[2409])
         );
  DFFPOSX1 reg_file_reg_18__106_ ( .D(n22718), .CLK(clk), .Q(reg_file[2410])
         );
  DFFPOSX1 reg_file_reg_18__107_ ( .D(n22717), .CLK(clk), .Q(reg_file[2411])
         );
  DFFPOSX1 reg_file_reg_18__108_ ( .D(n22716), .CLK(clk), .Q(reg_file[2412])
         );
  DFFPOSX1 reg_file_reg_18__109_ ( .D(n22715), .CLK(clk), .Q(reg_file[2413])
         );
  DFFPOSX1 reg_file_reg_18__110_ ( .D(n22714), .CLK(clk), .Q(reg_file[2414])
         );
  DFFPOSX1 reg_file_reg_18__111_ ( .D(n22713), .CLK(clk), .Q(reg_file[2415])
         );
  DFFPOSX1 reg_file_reg_18__112_ ( .D(n22712), .CLK(clk), .Q(reg_file[2416])
         );
  DFFPOSX1 reg_file_reg_18__113_ ( .D(n22711), .CLK(clk), .Q(reg_file[2417])
         );
  DFFPOSX1 reg_file_reg_18__114_ ( .D(n22710), .CLK(clk), .Q(reg_file[2418])
         );
  DFFPOSX1 reg_file_reg_18__115_ ( .D(n22709), .CLK(clk), .Q(reg_file[2419])
         );
  DFFPOSX1 reg_file_reg_18__116_ ( .D(n22708), .CLK(clk), .Q(reg_file[2420])
         );
  DFFPOSX1 reg_file_reg_18__117_ ( .D(n22707), .CLK(clk), .Q(reg_file[2421])
         );
  DFFPOSX1 reg_file_reg_18__118_ ( .D(n22706), .CLK(clk), .Q(reg_file[2422])
         );
  DFFPOSX1 reg_file_reg_18__119_ ( .D(n22705), .CLK(clk), .Q(reg_file[2423])
         );
  DFFPOSX1 reg_file_reg_18__120_ ( .D(n22704), .CLK(clk), .Q(reg_file[2424])
         );
  DFFPOSX1 reg_file_reg_18__121_ ( .D(n22703), .CLK(clk), .Q(reg_file[2425])
         );
  DFFPOSX1 reg_file_reg_18__122_ ( .D(n22702), .CLK(clk), .Q(reg_file[2426])
         );
  DFFPOSX1 reg_file_reg_18__123_ ( .D(n22701), .CLK(clk), .Q(reg_file[2427])
         );
  DFFPOSX1 reg_file_reg_18__124_ ( .D(n22700), .CLK(clk), .Q(reg_file[2428])
         );
  DFFPOSX1 reg_file_reg_18__125_ ( .D(n22699), .CLK(clk), .Q(reg_file[2429])
         );
  DFFPOSX1 reg_file_reg_18__126_ ( .D(n22698), .CLK(clk), .Q(reg_file[2430])
         );
  DFFPOSX1 reg_file_reg_18__127_ ( .D(n22697), .CLK(clk), .Q(reg_file[2431])
         );
  DFFPOSX1 reg_file_reg_19__0_ ( .D(n22696), .CLK(clk), .Q(reg_file[2432]) );
  DFFPOSX1 reg_file_reg_19__1_ ( .D(n22695), .CLK(clk), .Q(reg_file[2433]) );
  DFFPOSX1 reg_file_reg_19__2_ ( .D(n22694), .CLK(clk), .Q(reg_file[2434]) );
  DFFPOSX1 reg_file_reg_19__3_ ( .D(n22693), .CLK(clk), .Q(reg_file[2435]) );
  DFFPOSX1 reg_file_reg_19__4_ ( .D(n22692), .CLK(clk), .Q(reg_file[2436]) );
  DFFPOSX1 reg_file_reg_19__5_ ( .D(n22691), .CLK(clk), .Q(reg_file[2437]) );
  DFFPOSX1 reg_file_reg_19__6_ ( .D(n22690), .CLK(clk), .Q(reg_file[2438]) );
  DFFPOSX1 reg_file_reg_19__7_ ( .D(n22689), .CLK(clk), .Q(reg_file[2439]) );
  DFFPOSX1 reg_file_reg_19__8_ ( .D(n22688), .CLK(clk), .Q(reg_file[2440]) );
  DFFPOSX1 reg_file_reg_19__9_ ( .D(n22687), .CLK(clk), .Q(reg_file[2441]) );
  DFFPOSX1 reg_file_reg_19__10_ ( .D(n22686), .CLK(clk), .Q(reg_file[2442]) );
  DFFPOSX1 reg_file_reg_19__11_ ( .D(n22685), .CLK(clk), .Q(reg_file[2443]) );
  DFFPOSX1 reg_file_reg_19__12_ ( .D(n22684), .CLK(clk), .Q(reg_file[2444]) );
  DFFPOSX1 reg_file_reg_19__13_ ( .D(n22683), .CLK(clk), .Q(reg_file[2445]) );
  DFFPOSX1 reg_file_reg_19__14_ ( .D(n22682), .CLK(clk), .Q(reg_file[2446]) );
  DFFPOSX1 reg_file_reg_19__15_ ( .D(n22681), .CLK(clk), .Q(reg_file[2447]) );
  DFFPOSX1 reg_file_reg_19__16_ ( .D(n22680), .CLK(clk), .Q(reg_file[2448]) );
  DFFPOSX1 reg_file_reg_19__17_ ( .D(n22679), .CLK(clk), .Q(reg_file[2449]) );
  DFFPOSX1 reg_file_reg_19__18_ ( .D(n22678), .CLK(clk), .Q(reg_file[2450]) );
  DFFPOSX1 reg_file_reg_19__19_ ( .D(n22677), .CLK(clk), .Q(reg_file[2451]) );
  DFFPOSX1 reg_file_reg_19__20_ ( .D(n22676), .CLK(clk), .Q(reg_file[2452]) );
  DFFPOSX1 reg_file_reg_19__21_ ( .D(n22675), .CLK(clk), .Q(reg_file[2453]) );
  DFFPOSX1 reg_file_reg_19__22_ ( .D(n22674), .CLK(clk), .Q(reg_file[2454]) );
  DFFPOSX1 reg_file_reg_19__23_ ( .D(n22673), .CLK(clk), .Q(reg_file[2455]) );
  DFFPOSX1 reg_file_reg_19__24_ ( .D(n22672), .CLK(clk), .Q(reg_file[2456]) );
  DFFPOSX1 reg_file_reg_19__25_ ( .D(n22671), .CLK(clk), .Q(reg_file[2457]) );
  DFFPOSX1 reg_file_reg_19__26_ ( .D(n22670), .CLK(clk), .Q(reg_file[2458]) );
  DFFPOSX1 reg_file_reg_19__27_ ( .D(n22669), .CLK(clk), .Q(reg_file[2459]) );
  DFFPOSX1 reg_file_reg_19__28_ ( .D(n22668), .CLK(clk), .Q(reg_file[2460]) );
  DFFPOSX1 reg_file_reg_19__29_ ( .D(n22667), .CLK(clk), .Q(reg_file[2461]) );
  DFFPOSX1 reg_file_reg_19__30_ ( .D(n22666), .CLK(clk), .Q(reg_file[2462]) );
  DFFPOSX1 reg_file_reg_19__31_ ( .D(n22665), .CLK(clk), .Q(reg_file[2463]) );
  DFFPOSX1 reg_file_reg_19__32_ ( .D(n22664), .CLK(clk), .Q(reg_file[2464]) );
  DFFPOSX1 reg_file_reg_19__33_ ( .D(n22663), .CLK(clk), .Q(reg_file[2465]) );
  DFFPOSX1 reg_file_reg_19__34_ ( .D(n22662), .CLK(clk), .Q(reg_file[2466]) );
  DFFPOSX1 reg_file_reg_19__35_ ( .D(n22661), .CLK(clk), .Q(reg_file[2467]) );
  DFFPOSX1 reg_file_reg_19__36_ ( .D(n22660), .CLK(clk), .Q(reg_file[2468]) );
  DFFPOSX1 reg_file_reg_19__37_ ( .D(n22659), .CLK(clk), .Q(reg_file[2469]) );
  DFFPOSX1 reg_file_reg_19__38_ ( .D(n22658), .CLK(clk), .Q(reg_file[2470]) );
  DFFPOSX1 reg_file_reg_19__39_ ( .D(n22657), .CLK(clk), .Q(reg_file[2471]) );
  DFFPOSX1 reg_file_reg_19__40_ ( .D(n22656), .CLK(clk), .Q(reg_file[2472]) );
  DFFPOSX1 reg_file_reg_19__41_ ( .D(n22655), .CLK(clk), .Q(reg_file[2473]) );
  DFFPOSX1 reg_file_reg_19__42_ ( .D(n22654), .CLK(clk), .Q(reg_file[2474]) );
  DFFPOSX1 reg_file_reg_19__43_ ( .D(n22653), .CLK(clk), .Q(reg_file[2475]) );
  DFFPOSX1 reg_file_reg_19__44_ ( .D(n22652), .CLK(clk), .Q(reg_file[2476]) );
  DFFPOSX1 reg_file_reg_19__45_ ( .D(n22651), .CLK(clk), .Q(reg_file[2477]) );
  DFFPOSX1 reg_file_reg_19__46_ ( .D(n22650), .CLK(clk), .Q(reg_file[2478]) );
  DFFPOSX1 reg_file_reg_19__47_ ( .D(n22649), .CLK(clk), .Q(reg_file[2479]) );
  DFFPOSX1 reg_file_reg_19__48_ ( .D(n22648), .CLK(clk), .Q(reg_file[2480]) );
  DFFPOSX1 reg_file_reg_19__49_ ( .D(n22647), .CLK(clk), .Q(reg_file[2481]) );
  DFFPOSX1 reg_file_reg_19__50_ ( .D(n22646), .CLK(clk), .Q(reg_file[2482]) );
  DFFPOSX1 reg_file_reg_19__51_ ( .D(n22645), .CLK(clk), .Q(reg_file[2483]) );
  DFFPOSX1 reg_file_reg_19__52_ ( .D(n22644), .CLK(clk), .Q(reg_file[2484]) );
  DFFPOSX1 reg_file_reg_19__53_ ( .D(n22643), .CLK(clk), .Q(reg_file[2485]) );
  DFFPOSX1 reg_file_reg_19__54_ ( .D(n22642), .CLK(clk), .Q(reg_file[2486]) );
  DFFPOSX1 reg_file_reg_19__55_ ( .D(n22641), .CLK(clk), .Q(reg_file[2487]) );
  DFFPOSX1 reg_file_reg_19__56_ ( .D(n22640), .CLK(clk), .Q(reg_file[2488]) );
  DFFPOSX1 reg_file_reg_19__57_ ( .D(n22639), .CLK(clk), .Q(reg_file[2489]) );
  DFFPOSX1 reg_file_reg_19__58_ ( .D(n22638), .CLK(clk), .Q(reg_file[2490]) );
  DFFPOSX1 reg_file_reg_19__59_ ( .D(n22637), .CLK(clk), .Q(reg_file[2491]) );
  DFFPOSX1 reg_file_reg_19__60_ ( .D(n22636), .CLK(clk), .Q(reg_file[2492]) );
  DFFPOSX1 reg_file_reg_19__61_ ( .D(n22635), .CLK(clk), .Q(reg_file[2493]) );
  DFFPOSX1 reg_file_reg_19__62_ ( .D(n22634), .CLK(clk), .Q(reg_file[2494]) );
  DFFPOSX1 reg_file_reg_19__63_ ( .D(n22633), .CLK(clk), .Q(reg_file[2495]) );
  DFFPOSX1 reg_file_reg_19__64_ ( .D(n22632), .CLK(clk), .Q(reg_file[2496]) );
  DFFPOSX1 reg_file_reg_19__65_ ( .D(n22631), .CLK(clk), .Q(reg_file[2497]) );
  DFFPOSX1 reg_file_reg_19__66_ ( .D(n22630), .CLK(clk), .Q(reg_file[2498]) );
  DFFPOSX1 reg_file_reg_19__67_ ( .D(n22629), .CLK(clk), .Q(reg_file[2499]) );
  DFFPOSX1 reg_file_reg_19__68_ ( .D(n22628), .CLK(clk), .Q(reg_file[2500]) );
  DFFPOSX1 reg_file_reg_19__69_ ( .D(n22627), .CLK(clk), .Q(reg_file[2501]) );
  DFFPOSX1 reg_file_reg_19__70_ ( .D(n22626), .CLK(clk), .Q(reg_file[2502]) );
  DFFPOSX1 reg_file_reg_19__71_ ( .D(n22625), .CLK(clk), .Q(reg_file[2503]) );
  DFFPOSX1 reg_file_reg_19__72_ ( .D(n22624), .CLK(clk), .Q(reg_file[2504]) );
  DFFPOSX1 reg_file_reg_19__73_ ( .D(n22623), .CLK(clk), .Q(reg_file[2505]) );
  DFFPOSX1 reg_file_reg_19__74_ ( .D(n22622), .CLK(clk), .Q(reg_file[2506]) );
  DFFPOSX1 reg_file_reg_19__75_ ( .D(n22621), .CLK(clk), .Q(reg_file[2507]) );
  DFFPOSX1 reg_file_reg_19__76_ ( .D(n22620), .CLK(clk), .Q(reg_file[2508]) );
  DFFPOSX1 reg_file_reg_19__77_ ( .D(n22619), .CLK(clk), .Q(reg_file[2509]) );
  DFFPOSX1 reg_file_reg_19__78_ ( .D(n22618), .CLK(clk), .Q(reg_file[2510]) );
  DFFPOSX1 reg_file_reg_19__79_ ( .D(n22617), .CLK(clk), .Q(reg_file[2511]) );
  DFFPOSX1 reg_file_reg_19__80_ ( .D(n22616), .CLK(clk), .Q(reg_file[2512]) );
  DFFPOSX1 reg_file_reg_19__81_ ( .D(n22615), .CLK(clk), .Q(reg_file[2513]) );
  DFFPOSX1 reg_file_reg_19__82_ ( .D(n22614), .CLK(clk), .Q(reg_file[2514]) );
  DFFPOSX1 reg_file_reg_19__83_ ( .D(n22613), .CLK(clk), .Q(reg_file[2515]) );
  DFFPOSX1 reg_file_reg_19__84_ ( .D(n22612), .CLK(clk), .Q(reg_file[2516]) );
  DFFPOSX1 reg_file_reg_19__85_ ( .D(n22611), .CLK(clk), .Q(reg_file[2517]) );
  DFFPOSX1 reg_file_reg_19__86_ ( .D(n22610), .CLK(clk), .Q(reg_file[2518]) );
  DFFPOSX1 reg_file_reg_19__87_ ( .D(n22609), .CLK(clk), .Q(reg_file[2519]) );
  DFFPOSX1 reg_file_reg_19__88_ ( .D(n22608), .CLK(clk), .Q(reg_file[2520]) );
  DFFPOSX1 reg_file_reg_19__89_ ( .D(n22607), .CLK(clk), .Q(reg_file[2521]) );
  DFFPOSX1 reg_file_reg_19__90_ ( .D(n22606), .CLK(clk), .Q(reg_file[2522]) );
  DFFPOSX1 reg_file_reg_19__91_ ( .D(n22605), .CLK(clk), .Q(reg_file[2523]) );
  DFFPOSX1 reg_file_reg_19__92_ ( .D(n22604), .CLK(clk), .Q(reg_file[2524]) );
  DFFPOSX1 reg_file_reg_19__93_ ( .D(n22603), .CLK(clk), .Q(reg_file[2525]) );
  DFFPOSX1 reg_file_reg_19__94_ ( .D(n22602), .CLK(clk), .Q(reg_file[2526]) );
  DFFPOSX1 reg_file_reg_19__95_ ( .D(n22601), .CLK(clk), .Q(reg_file[2527]) );
  DFFPOSX1 reg_file_reg_19__96_ ( .D(n22600), .CLK(clk), .Q(reg_file[2528]) );
  DFFPOSX1 reg_file_reg_19__97_ ( .D(n22599), .CLK(clk), .Q(reg_file[2529]) );
  DFFPOSX1 reg_file_reg_19__98_ ( .D(n22598), .CLK(clk), .Q(reg_file[2530]) );
  DFFPOSX1 reg_file_reg_19__99_ ( .D(n22597), .CLK(clk), .Q(reg_file[2531]) );
  DFFPOSX1 reg_file_reg_19__100_ ( .D(n22596), .CLK(clk), .Q(reg_file[2532])
         );
  DFFPOSX1 reg_file_reg_19__101_ ( .D(n22595), .CLK(clk), .Q(reg_file[2533])
         );
  DFFPOSX1 reg_file_reg_19__102_ ( .D(n22594), .CLK(clk), .Q(reg_file[2534])
         );
  DFFPOSX1 reg_file_reg_19__103_ ( .D(n22593), .CLK(clk), .Q(reg_file[2535])
         );
  DFFPOSX1 reg_file_reg_19__104_ ( .D(n22592), .CLK(clk), .Q(reg_file[2536])
         );
  DFFPOSX1 reg_file_reg_19__105_ ( .D(n22591), .CLK(clk), .Q(reg_file[2537])
         );
  DFFPOSX1 reg_file_reg_19__106_ ( .D(n22590), .CLK(clk), .Q(reg_file[2538])
         );
  DFFPOSX1 reg_file_reg_19__107_ ( .D(n22589), .CLK(clk), .Q(reg_file[2539])
         );
  DFFPOSX1 reg_file_reg_19__108_ ( .D(n22588), .CLK(clk), .Q(reg_file[2540])
         );
  DFFPOSX1 reg_file_reg_19__109_ ( .D(n22587), .CLK(clk), .Q(reg_file[2541])
         );
  DFFPOSX1 reg_file_reg_19__110_ ( .D(n22586), .CLK(clk), .Q(reg_file[2542])
         );
  DFFPOSX1 reg_file_reg_19__111_ ( .D(n22585), .CLK(clk), .Q(reg_file[2543])
         );
  DFFPOSX1 reg_file_reg_19__112_ ( .D(n22584), .CLK(clk), .Q(reg_file[2544])
         );
  DFFPOSX1 reg_file_reg_19__113_ ( .D(n22583), .CLK(clk), .Q(reg_file[2545])
         );
  DFFPOSX1 reg_file_reg_19__114_ ( .D(n22582), .CLK(clk), .Q(reg_file[2546])
         );
  DFFPOSX1 reg_file_reg_19__115_ ( .D(n22581), .CLK(clk), .Q(reg_file[2547])
         );
  DFFPOSX1 reg_file_reg_19__116_ ( .D(n22580), .CLK(clk), .Q(reg_file[2548])
         );
  DFFPOSX1 reg_file_reg_19__117_ ( .D(n22579), .CLK(clk), .Q(reg_file[2549])
         );
  DFFPOSX1 reg_file_reg_19__118_ ( .D(n22578), .CLK(clk), .Q(reg_file[2550])
         );
  DFFPOSX1 reg_file_reg_19__119_ ( .D(n22577), .CLK(clk), .Q(reg_file[2551])
         );
  DFFPOSX1 reg_file_reg_19__120_ ( .D(n22576), .CLK(clk), .Q(reg_file[2552])
         );
  DFFPOSX1 reg_file_reg_19__121_ ( .D(n22575), .CLK(clk), .Q(reg_file[2553])
         );
  DFFPOSX1 reg_file_reg_19__122_ ( .D(n22574), .CLK(clk), .Q(reg_file[2554])
         );
  DFFPOSX1 reg_file_reg_19__123_ ( .D(n22573), .CLK(clk), .Q(reg_file[2555])
         );
  DFFPOSX1 reg_file_reg_19__124_ ( .D(n22572), .CLK(clk), .Q(reg_file[2556])
         );
  DFFPOSX1 reg_file_reg_19__125_ ( .D(n22571), .CLK(clk), .Q(reg_file[2557])
         );
  DFFPOSX1 reg_file_reg_19__126_ ( .D(n22570), .CLK(clk), .Q(reg_file[2558])
         );
  DFFPOSX1 reg_file_reg_19__127_ ( .D(n22569), .CLK(clk), .Q(reg_file[2559])
         );
  DFFPOSX1 reg_file_reg_20__0_ ( .D(n22568), .CLK(clk), .Q(reg_file[2560]) );
  DFFPOSX1 reg_file_reg_20__1_ ( .D(n22567), .CLK(clk), .Q(reg_file[2561]) );
  DFFPOSX1 reg_file_reg_20__2_ ( .D(n22566), .CLK(clk), .Q(reg_file[2562]) );
  DFFPOSX1 reg_file_reg_20__3_ ( .D(n22565), .CLK(clk), .Q(reg_file[2563]) );
  DFFPOSX1 reg_file_reg_20__4_ ( .D(n22564), .CLK(clk), .Q(reg_file[2564]) );
  DFFPOSX1 reg_file_reg_20__5_ ( .D(n22563), .CLK(clk), .Q(reg_file[2565]) );
  DFFPOSX1 reg_file_reg_20__6_ ( .D(n22562), .CLK(clk), .Q(reg_file[2566]) );
  DFFPOSX1 reg_file_reg_20__7_ ( .D(n22561), .CLK(clk), .Q(reg_file[2567]) );
  DFFPOSX1 reg_file_reg_20__8_ ( .D(n22560), .CLK(clk), .Q(reg_file[2568]) );
  DFFPOSX1 reg_file_reg_20__9_ ( .D(n22559), .CLK(clk), .Q(reg_file[2569]) );
  DFFPOSX1 reg_file_reg_20__10_ ( .D(n22558), .CLK(clk), .Q(reg_file[2570]) );
  DFFPOSX1 reg_file_reg_20__11_ ( .D(n22557), .CLK(clk), .Q(reg_file[2571]) );
  DFFPOSX1 reg_file_reg_20__12_ ( .D(n22556), .CLK(clk), .Q(reg_file[2572]) );
  DFFPOSX1 reg_file_reg_20__13_ ( .D(n22555), .CLK(clk), .Q(reg_file[2573]) );
  DFFPOSX1 reg_file_reg_20__14_ ( .D(n22554), .CLK(clk), .Q(reg_file[2574]) );
  DFFPOSX1 reg_file_reg_20__15_ ( .D(n22553), .CLK(clk), .Q(reg_file[2575]) );
  DFFPOSX1 reg_file_reg_20__16_ ( .D(n22552), .CLK(clk), .Q(reg_file[2576]) );
  DFFPOSX1 reg_file_reg_20__17_ ( .D(n22551), .CLK(clk), .Q(reg_file[2577]) );
  DFFPOSX1 reg_file_reg_20__18_ ( .D(n22550), .CLK(clk), .Q(reg_file[2578]) );
  DFFPOSX1 reg_file_reg_20__19_ ( .D(n22549), .CLK(clk), .Q(reg_file[2579]) );
  DFFPOSX1 reg_file_reg_20__20_ ( .D(n22548), .CLK(clk), .Q(reg_file[2580]) );
  DFFPOSX1 reg_file_reg_20__21_ ( .D(n22547), .CLK(clk), .Q(reg_file[2581]) );
  DFFPOSX1 reg_file_reg_20__22_ ( .D(n22546), .CLK(clk), .Q(reg_file[2582]) );
  DFFPOSX1 reg_file_reg_20__23_ ( .D(n22545), .CLK(clk), .Q(reg_file[2583]) );
  DFFPOSX1 reg_file_reg_20__24_ ( .D(n22544), .CLK(clk), .Q(reg_file[2584]) );
  DFFPOSX1 reg_file_reg_20__25_ ( .D(n22543), .CLK(clk), .Q(reg_file[2585]) );
  DFFPOSX1 reg_file_reg_20__26_ ( .D(n22542), .CLK(clk), .Q(reg_file[2586]) );
  DFFPOSX1 reg_file_reg_20__27_ ( .D(n22541), .CLK(clk), .Q(reg_file[2587]) );
  DFFPOSX1 reg_file_reg_20__28_ ( .D(n22540), .CLK(clk), .Q(reg_file[2588]) );
  DFFPOSX1 reg_file_reg_20__29_ ( .D(n22539), .CLK(clk), .Q(reg_file[2589]) );
  DFFPOSX1 reg_file_reg_20__30_ ( .D(n22538), .CLK(clk), .Q(reg_file[2590]) );
  DFFPOSX1 reg_file_reg_20__31_ ( .D(n22537), .CLK(clk), .Q(reg_file[2591]) );
  DFFPOSX1 reg_file_reg_20__32_ ( .D(n22536), .CLK(clk), .Q(reg_file[2592]) );
  DFFPOSX1 reg_file_reg_20__33_ ( .D(n22535), .CLK(clk), .Q(reg_file[2593]) );
  DFFPOSX1 reg_file_reg_20__34_ ( .D(n22534), .CLK(clk), .Q(reg_file[2594]) );
  DFFPOSX1 reg_file_reg_20__35_ ( .D(n22533), .CLK(clk), .Q(reg_file[2595]) );
  DFFPOSX1 reg_file_reg_20__36_ ( .D(n22532), .CLK(clk), .Q(reg_file[2596]) );
  DFFPOSX1 reg_file_reg_20__37_ ( .D(n22531), .CLK(clk), .Q(reg_file[2597]) );
  DFFPOSX1 reg_file_reg_20__38_ ( .D(n22530), .CLK(clk), .Q(reg_file[2598]) );
  DFFPOSX1 reg_file_reg_20__39_ ( .D(n22529), .CLK(clk), .Q(reg_file[2599]) );
  DFFPOSX1 reg_file_reg_20__40_ ( .D(n22528), .CLK(clk), .Q(reg_file[2600]) );
  DFFPOSX1 reg_file_reg_20__41_ ( .D(n22527), .CLK(clk), .Q(reg_file[2601]) );
  DFFPOSX1 reg_file_reg_20__42_ ( .D(n22526), .CLK(clk), .Q(reg_file[2602]) );
  DFFPOSX1 reg_file_reg_20__43_ ( .D(n22525), .CLK(clk), .Q(reg_file[2603]) );
  DFFPOSX1 reg_file_reg_20__44_ ( .D(n22524), .CLK(clk), .Q(reg_file[2604]) );
  DFFPOSX1 reg_file_reg_20__45_ ( .D(n22523), .CLK(clk), .Q(reg_file[2605]) );
  DFFPOSX1 reg_file_reg_20__46_ ( .D(n22522), .CLK(clk), .Q(reg_file[2606]) );
  DFFPOSX1 reg_file_reg_20__47_ ( .D(n22521), .CLK(clk), .Q(reg_file[2607]) );
  DFFPOSX1 reg_file_reg_20__48_ ( .D(n22520), .CLK(clk), .Q(reg_file[2608]) );
  DFFPOSX1 reg_file_reg_20__49_ ( .D(n22519), .CLK(clk), .Q(reg_file[2609]) );
  DFFPOSX1 reg_file_reg_20__50_ ( .D(n22518), .CLK(clk), .Q(reg_file[2610]) );
  DFFPOSX1 reg_file_reg_20__51_ ( .D(n22517), .CLK(clk), .Q(reg_file[2611]) );
  DFFPOSX1 reg_file_reg_20__52_ ( .D(n22516), .CLK(clk), .Q(reg_file[2612]) );
  DFFPOSX1 reg_file_reg_20__53_ ( .D(n22515), .CLK(clk), .Q(reg_file[2613]) );
  DFFPOSX1 reg_file_reg_20__54_ ( .D(n22514), .CLK(clk), .Q(reg_file[2614]) );
  DFFPOSX1 reg_file_reg_20__55_ ( .D(n22513), .CLK(clk), .Q(reg_file[2615]) );
  DFFPOSX1 reg_file_reg_20__56_ ( .D(n22512), .CLK(clk), .Q(reg_file[2616]) );
  DFFPOSX1 reg_file_reg_20__57_ ( .D(n22511), .CLK(clk), .Q(reg_file[2617]) );
  DFFPOSX1 reg_file_reg_20__58_ ( .D(n22510), .CLK(clk), .Q(reg_file[2618]) );
  DFFPOSX1 reg_file_reg_20__59_ ( .D(n22509), .CLK(clk), .Q(reg_file[2619]) );
  DFFPOSX1 reg_file_reg_20__60_ ( .D(n22508), .CLK(clk), .Q(reg_file[2620]) );
  DFFPOSX1 reg_file_reg_20__61_ ( .D(n22507), .CLK(clk), .Q(reg_file[2621]) );
  DFFPOSX1 reg_file_reg_20__62_ ( .D(n22506), .CLK(clk), .Q(reg_file[2622]) );
  DFFPOSX1 reg_file_reg_20__63_ ( .D(n22505), .CLK(clk), .Q(reg_file[2623]) );
  DFFPOSX1 reg_file_reg_20__64_ ( .D(n22504), .CLK(clk), .Q(reg_file[2624]) );
  DFFPOSX1 reg_file_reg_20__65_ ( .D(n22503), .CLK(clk), .Q(reg_file[2625]) );
  DFFPOSX1 reg_file_reg_20__66_ ( .D(n22502), .CLK(clk), .Q(reg_file[2626]) );
  DFFPOSX1 reg_file_reg_20__67_ ( .D(n22501), .CLK(clk), .Q(reg_file[2627]) );
  DFFPOSX1 reg_file_reg_20__68_ ( .D(n22500), .CLK(clk), .Q(reg_file[2628]) );
  DFFPOSX1 reg_file_reg_20__69_ ( .D(n22499), .CLK(clk), .Q(reg_file[2629]) );
  DFFPOSX1 reg_file_reg_20__70_ ( .D(n22498), .CLK(clk), .Q(reg_file[2630]) );
  DFFPOSX1 reg_file_reg_20__71_ ( .D(n22497), .CLK(clk), .Q(reg_file[2631]) );
  DFFPOSX1 reg_file_reg_20__72_ ( .D(n22496), .CLK(clk), .Q(reg_file[2632]) );
  DFFPOSX1 reg_file_reg_20__73_ ( .D(n22495), .CLK(clk), .Q(reg_file[2633]) );
  DFFPOSX1 reg_file_reg_20__74_ ( .D(n22494), .CLK(clk), .Q(reg_file[2634]) );
  DFFPOSX1 reg_file_reg_20__75_ ( .D(n22493), .CLK(clk), .Q(reg_file[2635]) );
  DFFPOSX1 reg_file_reg_20__76_ ( .D(n22492), .CLK(clk), .Q(reg_file[2636]) );
  DFFPOSX1 reg_file_reg_20__77_ ( .D(n22491), .CLK(clk), .Q(reg_file[2637]) );
  DFFPOSX1 reg_file_reg_20__78_ ( .D(n22490), .CLK(clk), .Q(reg_file[2638]) );
  DFFPOSX1 reg_file_reg_20__79_ ( .D(n22489), .CLK(clk), .Q(reg_file[2639]) );
  DFFPOSX1 reg_file_reg_20__80_ ( .D(n22488), .CLK(clk), .Q(reg_file[2640]) );
  DFFPOSX1 reg_file_reg_20__81_ ( .D(n22487), .CLK(clk), .Q(reg_file[2641]) );
  DFFPOSX1 reg_file_reg_20__82_ ( .D(n22486), .CLK(clk), .Q(reg_file[2642]) );
  DFFPOSX1 reg_file_reg_20__83_ ( .D(n22485), .CLK(clk), .Q(reg_file[2643]) );
  DFFPOSX1 reg_file_reg_20__84_ ( .D(n22484), .CLK(clk), .Q(reg_file[2644]) );
  DFFPOSX1 reg_file_reg_20__85_ ( .D(n22483), .CLK(clk), .Q(reg_file[2645]) );
  DFFPOSX1 reg_file_reg_20__86_ ( .D(n22482), .CLK(clk), .Q(reg_file[2646]) );
  DFFPOSX1 reg_file_reg_20__87_ ( .D(n22481), .CLK(clk), .Q(reg_file[2647]) );
  DFFPOSX1 reg_file_reg_20__88_ ( .D(n22480), .CLK(clk), .Q(reg_file[2648]) );
  DFFPOSX1 reg_file_reg_20__89_ ( .D(n22479), .CLK(clk), .Q(reg_file[2649]) );
  DFFPOSX1 reg_file_reg_20__90_ ( .D(n22478), .CLK(clk), .Q(reg_file[2650]) );
  DFFPOSX1 reg_file_reg_20__91_ ( .D(n22477), .CLK(clk), .Q(reg_file[2651]) );
  DFFPOSX1 reg_file_reg_20__92_ ( .D(n22476), .CLK(clk), .Q(reg_file[2652]) );
  DFFPOSX1 reg_file_reg_20__93_ ( .D(n22475), .CLK(clk), .Q(reg_file[2653]) );
  DFFPOSX1 reg_file_reg_20__94_ ( .D(n22474), .CLK(clk), .Q(reg_file[2654]) );
  DFFPOSX1 reg_file_reg_20__95_ ( .D(n22473), .CLK(clk), .Q(reg_file[2655]) );
  DFFPOSX1 reg_file_reg_20__96_ ( .D(n22472), .CLK(clk), .Q(reg_file[2656]) );
  DFFPOSX1 reg_file_reg_20__97_ ( .D(n22471), .CLK(clk), .Q(reg_file[2657]) );
  DFFPOSX1 reg_file_reg_20__98_ ( .D(n22470), .CLK(clk), .Q(reg_file[2658]) );
  DFFPOSX1 reg_file_reg_20__99_ ( .D(n22469), .CLK(clk), .Q(reg_file[2659]) );
  DFFPOSX1 reg_file_reg_20__100_ ( .D(n22468), .CLK(clk), .Q(reg_file[2660])
         );
  DFFPOSX1 reg_file_reg_20__101_ ( .D(n22467), .CLK(clk), .Q(reg_file[2661])
         );
  DFFPOSX1 reg_file_reg_20__102_ ( .D(n22466), .CLK(clk), .Q(reg_file[2662])
         );
  DFFPOSX1 reg_file_reg_20__103_ ( .D(n22465), .CLK(clk), .Q(reg_file[2663])
         );
  DFFPOSX1 reg_file_reg_20__104_ ( .D(n22464), .CLK(clk), .Q(reg_file[2664])
         );
  DFFPOSX1 reg_file_reg_20__105_ ( .D(n22463), .CLK(clk), .Q(reg_file[2665])
         );
  DFFPOSX1 reg_file_reg_20__106_ ( .D(n22462), .CLK(clk), .Q(reg_file[2666])
         );
  DFFPOSX1 reg_file_reg_20__107_ ( .D(n22461), .CLK(clk), .Q(reg_file[2667])
         );
  DFFPOSX1 reg_file_reg_20__108_ ( .D(n22460), .CLK(clk), .Q(reg_file[2668])
         );
  DFFPOSX1 reg_file_reg_20__109_ ( .D(n22459), .CLK(clk), .Q(reg_file[2669])
         );
  DFFPOSX1 reg_file_reg_20__110_ ( .D(n22458), .CLK(clk), .Q(reg_file[2670])
         );
  DFFPOSX1 reg_file_reg_20__111_ ( .D(n22457), .CLK(clk), .Q(reg_file[2671])
         );
  DFFPOSX1 reg_file_reg_20__112_ ( .D(n22456), .CLK(clk), .Q(reg_file[2672])
         );
  DFFPOSX1 reg_file_reg_20__113_ ( .D(n22455), .CLK(clk), .Q(reg_file[2673])
         );
  DFFPOSX1 reg_file_reg_20__114_ ( .D(n22454), .CLK(clk), .Q(reg_file[2674])
         );
  DFFPOSX1 reg_file_reg_20__115_ ( .D(n22453), .CLK(clk), .Q(reg_file[2675])
         );
  DFFPOSX1 reg_file_reg_20__116_ ( .D(n22452), .CLK(clk), .Q(reg_file[2676])
         );
  DFFPOSX1 reg_file_reg_20__117_ ( .D(n22451), .CLK(clk), .Q(reg_file[2677])
         );
  DFFPOSX1 reg_file_reg_20__118_ ( .D(n22450), .CLK(clk), .Q(reg_file[2678])
         );
  DFFPOSX1 reg_file_reg_20__119_ ( .D(n22449), .CLK(clk), .Q(reg_file[2679])
         );
  DFFPOSX1 reg_file_reg_20__120_ ( .D(n22448), .CLK(clk), .Q(reg_file[2680])
         );
  DFFPOSX1 reg_file_reg_20__121_ ( .D(n22447), .CLK(clk), .Q(reg_file[2681])
         );
  DFFPOSX1 reg_file_reg_20__122_ ( .D(n22446), .CLK(clk), .Q(reg_file[2682])
         );
  DFFPOSX1 reg_file_reg_20__123_ ( .D(n22445), .CLK(clk), .Q(reg_file[2683])
         );
  DFFPOSX1 reg_file_reg_20__124_ ( .D(n22444), .CLK(clk), .Q(reg_file[2684])
         );
  DFFPOSX1 reg_file_reg_20__125_ ( .D(n22443), .CLK(clk), .Q(reg_file[2685])
         );
  DFFPOSX1 reg_file_reg_20__126_ ( .D(n22442), .CLK(clk), .Q(reg_file[2686])
         );
  DFFPOSX1 reg_file_reg_20__127_ ( .D(n22441), .CLK(clk), .Q(reg_file[2687])
         );
  DFFPOSX1 reg_file_reg_21__0_ ( .D(n22440), .CLK(clk), .Q(reg_file[2688]) );
  DFFPOSX1 reg_file_reg_21__1_ ( .D(n22439), .CLK(clk), .Q(reg_file[2689]) );
  DFFPOSX1 reg_file_reg_21__2_ ( .D(n22438), .CLK(clk), .Q(reg_file[2690]) );
  DFFPOSX1 reg_file_reg_21__3_ ( .D(n22437), .CLK(clk), .Q(reg_file[2691]) );
  DFFPOSX1 reg_file_reg_21__4_ ( .D(n22436), .CLK(clk), .Q(reg_file[2692]) );
  DFFPOSX1 reg_file_reg_21__5_ ( .D(n22435), .CLK(clk), .Q(reg_file[2693]) );
  DFFPOSX1 reg_file_reg_21__6_ ( .D(n22434), .CLK(clk), .Q(reg_file[2694]) );
  DFFPOSX1 reg_file_reg_21__7_ ( .D(n22433), .CLK(clk), .Q(reg_file[2695]) );
  DFFPOSX1 reg_file_reg_21__8_ ( .D(n22432), .CLK(clk), .Q(reg_file[2696]) );
  DFFPOSX1 reg_file_reg_21__9_ ( .D(n22431), .CLK(clk), .Q(reg_file[2697]) );
  DFFPOSX1 reg_file_reg_21__10_ ( .D(n22430), .CLK(clk), .Q(reg_file[2698]) );
  DFFPOSX1 reg_file_reg_21__11_ ( .D(n22429), .CLK(clk), .Q(reg_file[2699]) );
  DFFPOSX1 reg_file_reg_21__12_ ( .D(n22428), .CLK(clk), .Q(reg_file[2700]) );
  DFFPOSX1 reg_file_reg_21__13_ ( .D(n22427), .CLK(clk), .Q(reg_file[2701]) );
  DFFPOSX1 reg_file_reg_21__14_ ( .D(n22426), .CLK(clk), .Q(reg_file[2702]) );
  DFFPOSX1 reg_file_reg_21__15_ ( .D(n22425), .CLK(clk), .Q(reg_file[2703]) );
  DFFPOSX1 reg_file_reg_21__16_ ( .D(n22424), .CLK(clk), .Q(reg_file[2704]) );
  DFFPOSX1 reg_file_reg_21__17_ ( .D(n22423), .CLK(clk), .Q(reg_file[2705]) );
  DFFPOSX1 reg_file_reg_21__18_ ( .D(n22422), .CLK(clk), .Q(reg_file[2706]) );
  DFFPOSX1 reg_file_reg_21__19_ ( .D(n22421), .CLK(clk), .Q(reg_file[2707]) );
  DFFPOSX1 reg_file_reg_21__20_ ( .D(n22420), .CLK(clk), .Q(reg_file[2708]) );
  DFFPOSX1 reg_file_reg_21__21_ ( .D(n22419), .CLK(clk), .Q(reg_file[2709]) );
  DFFPOSX1 reg_file_reg_21__22_ ( .D(n22418), .CLK(clk), .Q(reg_file[2710]) );
  DFFPOSX1 reg_file_reg_21__23_ ( .D(n22417), .CLK(clk), .Q(reg_file[2711]) );
  DFFPOSX1 reg_file_reg_21__24_ ( .D(n22416), .CLK(clk), .Q(reg_file[2712]) );
  DFFPOSX1 reg_file_reg_21__25_ ( .D(n22415), .CLK(clk), .Q(reg_file[2713]) );
  DFFPOSX1 reg_file_reg_21__26_ ( .D(n22414), .CLK(clk), .Q(reg_file[2714]) );
  DFFPOSX1 reg_file_reg_21__27_ ( .D(n22413), .CLK(clk), .Q(reg_file[2715]) );
  DFFPOSX1 reg_file_reg_21__28_ ( .D(n22412), .CLK(clk), .Q(reg_file[2716]) );
  DFFPOSX1 reg_file_reg_21__29_ ( .D(n22411), .CLK(clk), .Q(reg_file[2717]) );
  DFFPOSX1 reg_file_reg_21__30_ ( .D(n22410), .CLK(clk), .Q(reg_file[2718]) );
  DFFPOSX1 reg_file_reg_21__31_ ( .D(n22409), .CLK(clk), .Q(reg_file[2719]) );
  DFFPOSX1 reg_file_reg_21__32_ ( .D(n22408), .CLK(clk), .Q(reg_file[2720]) );
  DFFPOSX1 reg_file_reg_21__33_ ( .D(n22407), .CLK(clk), .Q(reg_file[2721]) );
  DFFPOSX1 reg_file_reg_21__34_ ( .D(n22406), .CLK(clk), .Q(reg_file[2722]) );
  DFFPOSX1 reg_file_reg_21__35_ ( .D(n22405), .CLK(clk), .Q(reg_file[2723]) );
  DFFPOSX1 reg_file_reg_21__36_ ( .D(n22404), .CLK(clk), .Q(reg_file[2724]) );
  DFFPOSX1 reg_file_reg_21__37_ ( .D(n22403), .CLK(clk), .Q(reg_file[2725]) );
  DFFPOSX1 reg_file_reg_21__38_ ( .D(n22402), .CLK(clk), .Q(reg_file[2726]) );
  DFFPOSX1 reg_file_reg_21__39_ ( .D(n22401), .CLK(clk), .Q(reg_file[2727]) );
  DFFPOSX1 reg_file_reg_21__40_ ( .D(n22400), .CLK(clk), .Q(reg_file[2728]) );
  DFFPOSX1 reg_file_reg_21__41_ ( .D(n22399), .CLK(clk), .Q(reg_file[2729]) );
  DFFPOSX1 reg_file_reg_21__42_ ( .D(n22398), .CLK(clk), .Q(reg_file[2730]) );
  DFFPOSX1 reg_file_reg_21__43_ ( .D(n22397), .CLK(clk), .Q(reg_file[2731]) );
  DFFPOSX1 reg_file_reg_21__44_ ( .D(n22396), .CLK(clk), .Q(reg_file[2732]) );
  DFFPOSX1 reg_file_reg_21__45_ ( .D(n22395), .CLK(clk), .Q(reg_file[2733]) );
  DFFPOSX1 reg_file_reg_21__46_ ( .D(n22394), .CLK(clk), .Q(reg_file[2734]) );
  DFFPOSX1 reg_file_reg_21__47_ ( .D(n22393), .CLK(clk), .Q(reg_file[2735]) );
  DFFPOSX1 reg_file_reg_21__48_ ( .D(n22392), .CLK(clk), .Q(reg_file[2736]) );
  DFFPOSX1 reg_file_reg_21__49_ ( .D(n22391), .CLK(clk), .Q(reg_file[2737]) );
  DFFPOSX1 reg_file_reg_21__50_ ( .D(n22390), .CLK(clk), .Q(reg_file[2738]) );
  DFFPOSX1 reg_file_reg_21__51_ ( .D(n22389), .CLK(clk), .Q(reg_file[2739]) );
  DFFPOSX1 reg_file_reg_21__52_ ( .D(n22388), .CLK(clk), .Q(reg_file[2740]) );
  DFFPOSX1 reg_file_reg_21__53_ ( .D(n22387), .CLK(clk), .Q(reg_file[2741]) );
  DFFPOSX1 reg_file_reg_21__54_ ( .D(n22386), .CLK(clk), .Q(reg_file[2742]) );
  DFFPOSX1 reg_file_reg_21__55_ ( .D(n22385), .CLK(clk), .Q(reg_file[2743]) );
  DFFPOSX1 reg_file_reg_21__56_ ( .D(n22384), .CLK(clk), .Q(reg_file[2744]) );
  DFFPOSX1 reg_file_reg_21__57_ ( .D(n22383), .CLK(clk), .Q(reg_file[2745]) );
  DFFPOSX1 reg_file_reg_21__58_ ( .D(n22382), .CLK(clk), .Q(reg_file[2746]) );
  DFFPOSX1 reg_file_reg_21__59_ ( .D(n22381), .CLK(clk), .Q(reg_file[2747]) );
  DFFPOSX1 reg_file_reg_21__60_ ( .D(n22380), .CLK(clk), .Q(reg_file[2748]) );
  DFFPOSX1 reg_file_reg_21__61_ ( .D(n22379), .CLK(clk), .Q(reg_file[2749]) );
  DFFPOSX1 reg_file_reg_21__62_ ( .D(n22378), .CLK(clk), .Q(reg_file[2750]) );
  DFFPOSX1 reg_file_reg_21__63_ ( .D(n22377), .CLK(clk), .Q(reg_file[2751]) );
  DFFPOSX1 reg_file_reg_21__64_ ( .D(n22376), .CLK(clk), .Q(reg_file[2752]) );
  DFFPOSX1 reg_file_reg_21__65_ ( .D(n22375), .CLK(clk), .Q(reg_file[2753]) );
  DFFPOSX1 reg_file_reg_21__66_ ( .D(n22374), .CLK(clk), .Q(reg_file[2754]) );
  DFFPOSX1 reg_file_reg_21__67_ ( .D(n22373), .CLK(clk), .Q(reg_file[2755]) );
  DFFPOSX1 reg_file_reg_21__68_ ( .D(n22372), .CLK(clk), .Q(reg_file[2756]) );
  DFFPOSX1 reg_file_reg_21__69_ ( .D(n22371), .CLK(clk), .Q(reg_file[2757]) );
  DFFPOSX1 reg_file_reg_21__70_ ( .D(n22370), .CLK(clk), .Q(reg_file[2758]) );
  DFFPOSX1 reg_file_reg_21__71_ ( .D(n22369), .CLK(clk), .Q(reg_file[2759]) );
  DFFPOSX1 reg_file_reg_21__72_ ( .D(n22368), .CLK(clk), .Q(reg_file[2760]) );
  DFFPOSX1 reg_file_reg_21__73_ ( .D(n22367), .CLK(clk), .Q(reg_file[2761]) );
  DFFPOSX1 reg_file_reg_21__74_ ( .D(n22366), .CLK(clk), .Q(reg_file[2762]) );
  DFFPOSX1 reg_file_reg_21__75_ ( .D(n22365), .CLK(clk), .Q(reg_file[2763]) );
  DFFPOSX1 reg_file_reg_21__76_ ( .D(n22364), .CLK(clk), .Q(reg_file[2764]) );
  DFFPOSX1 reg_file_reg_21__77_ ( .D(n22363), .CLK(clk), .Q(reg_file[2765]) );
  DFFPOSX1 reg_file_reg_21__78_ ( .D(n22362), .CLK(clk), .Q(reg_file[2766]) );
  DFFPOSX1 reg_file_reg_21__79_ ( .D(n22361), .CLK(clk), .Q(reg_file[2767]) );
  DFFPOSX1 reg_file_reg_21__80_ ( .D(n22360), .CLK(clk), .Q(reg_file[2768]) );
  DFFPOSX1 reg_file_reg_21__81_ ( .D(n22359), .CLK(clk), .Q(reg_file[2769]) );
  DFFPOSX1 reg_file_reg_21__82_ ( .D(n22358), .CLK(clk), .Q(reg_file[2770]) );
  DFFPOSX1 reg_file_reg_21__83_ ( .D(n22357), .CLK(clk), .Q(reg_file[2771]) );
  DFFPOSX1 reg_file_reg_21__84_ ( .D(n22356), .CLK(clk), .Q(reg_file[2772]) );
  DFFPOSX1 reg_file_reg_21__85_ ( .D(n22355), .CLK(clk), .Q(reg_file[2773]) );
  DFFPOSX1 reg_file_reg_21__86_ ( .D(n22354), .CLK(clk), .Q(reg_file[2774]) );
  DFFPOSX1 reg_file_reg_21__87_ ( .D(n22353), .CLK(clk), .Q(reg_file[2775]) );
  DFFPOSX1 reg_file_reg_21__88_ ( .D(n22352), .CLK(clk), .Q(reg_file[2776]) );
  DFFPOSX1 reg_file_reg_21__89_ ( .D(n22351), .CLK(clk), .Q(reg_file[2777]) );
  DFFPOSX1 reg_file_reg_21__90_ ( .D(n22350), .CLK(clk), .Q(reg_file[2778]) );
  DFFPOSX1 reg_file_reg_21__91_ ( .D(n22349), .CLK(clk), .Q(reg_file[2779]) );
  DFFPOSX1 reg_file_reg_21__92_ ( .D(n22348), .CLK(clk), .Q(reg_file[2780]) );
  DFFPOSX1 reg_file_reg_21__93_ ( .D(n22347), .CLK(clk), .Q(reg_file[2781]) );
  DFFPOSX1 reg_file_reg_21__94_ ( .D(n22346), .CLK(clk), .Q(reg_file[2782]) );
  DFFPOSX1 reg_file_reg_21__95_ ( .D(n22345), .CLK(clk), .Q(reg_file[2783]) );
  DFFPOSX1 reg_file_reg_21__96_ ( .D(n22344), .CLK(clk), .Q(reg_file[2784]) );
  DFFPOSX1 reg_file_reg_21__97_ ( .D(n22343), .CLK(clk), .Q(reg_file[2785]) );
  DFFPOSX1 reg_file_reg_21__98_ ( .D(n22342), .CLK(clk), .Q(reg_file[2786]) );
  DFFPOSX1 reg_file_reg_21__99_ ( .D(n22341), .CLK(clk), .Q(reg_file[2787]) );
  DFFPOSX1 reg_file_reg_21__100_ ( .D(n22340), .CLK(clk), .Q(reg_file[2788])
         );
  DFFPOSX1 reg_file_reg_21__101_ ( .D(n22339), .CLK(clk), .Q(reg_file[2789])
         );
  DFFPOSX1 reg_file_reg_21__102_ ( .D(n22338), .CLK(clk), .Q(reg_file[2790])
         );
  DFFPOSX1 reg_file_reg_21__103_ ( .D(n22337), .CLK(clk), .Q(reg_file[2791])
         );
  DFFPOSX1 reg_file_reg_21__104_ ( .D(n22336), .CLK(clk), .Q(reg_file[2792])
         );
  DFFPOSX1 reg_file_reg_21__105_ ( .D(n22335), .CLK(clk), .Q(reg_file[2793])
         );
  DFFPOSX1 reg_file_reg_21__106_ ( .D(n22334), .CLK(clk), .Q(reg_file[2794])
         );
  DFFPOSX1 reg_file_reg_21__107_ ( .D(n22333), .CLK(clk), .Q(reg_file[2795])
         );
  DFFPOSX1 reg_file_reg_21__108_ ( .D(n22332), .CLK(clk), .Q(reg_file[2796])
         );
  DFFPOSX1 reg_file_reg_21__109_ ( .D(n22331), .CLK(clk), .Q(reg_file[2797])
         );
  DFFPOSX1 reg_file_reg_21__110_ ( .D(n22330), .CLK(clk), .Q(reg_file[2798])
         );
  DFFPOSX1 reg_file_reg_21__111_ ( .D(n22329), .CLK(clk), .Q(reg_file[2799])
         );
  DFFPOSX1 reg_file_reg_21__112_ ( .D(n22328), .CLK(clk), .Q(reg_file[2800])
         );
  DFFPOSX1 reg_file_reg_21__113_ ( .D(n22327), .CLK(clk), .Q(reg_file[2801])
         );
  DFFPOSX1 reg_file_reg_21__114_ ( .D(n22326), .CLK(clk), .Q(reg_file[2802])
         );
  DFFPOSX1 reg_file_reg_21__115_ ( .D(n22325), .CLK(clk), .Q(reg_file[2803])
         );
  DFFPOSX1 reg_file_reg_21__116_ ( .D(n22324), .CLK(clk), .Q(reg_file[2804])
         );
  DFFPOSX1 reg_file_reg_21__117_ ( .D(n22323), .CLK(clk), .Q(reg_file[2805])
         );
  DFFPOSX1 reg_file_reg_21__118_ ( .D(n22322), .CLK(clk), .Q(reg_file[2806])
         );
  DFFPOSX1 reg_file_reg_21__119_ ( .D(n22321), .CLK(clk), .Q(reg_file[2807])
         );
  DFFPOSX1 reg_file_reg_21__120_ ( .D(n22320), .CLK(clk), .Q(reg_file[2808])
         );
  DFFPOSX1 reg_file_reg_21__121_ ( .D(n22319), .CLK(clk), .Q(reg_file[2809])
         );
  DFFPOSX1 reg_file_reg_21__122_ ( .D(n22318), .CLK(clk), .Q(reg_file[2810])
         );
  DFFPOSX1 reg_file_reg_21__123_ ( .D(n22317), .CLK(clk), .Q(reg_file[2811])
         );
  DFFPOSX1 reg_file_reg_21__124_ ( .D(n22316), .CLK(clk), .Q(reg_file[2812])
         );
  DFFPOSX1 reg_file_reg_21__125_ ( .D(n22315), .CLK(clk), .Q(reg_file[2813])
         );
  DFFPOSX1 reg_file_reg_21__126_ ( .D(n22314), .CLK(clk), .Q(reg_file[2814])
         );
  DFFPOSX1 reg_file_reg_21__127_ ( .D(n22313), .CLK(clk), .Q(reg_file[2815])
         );
  DFFPOSX1 reg_file_reg_22__0_ ( .D(n22312), .CLK(clk), .Q(reg_file[2816]) );
  DFFPOSX1 reg_file_reg_22__1_ ( .D(n22311), .CLK(clk), .Q(reg_file[2817]) );
  DFFPOSX1 reg_file_reg_22__2_ ( .D(n22310), .CLK(clk), .Q(reg_file[2818]) );
  DFFPOSX1 reg_file_reg_22__3_ ( .D(n22309), .CLK(clk), .Q(reg_file[2819]) );
  DFFPOSX1 reg_file_reg_22__4_ ( .D(n22308), .CLK(clk), .Q(reg_file[2820]) );
  DFFPOSX1 reg_file_reg_22__5_ ( .D(n22307), .CLK(clk), .Q(reg_file[2821]) );
  DFFPOSX1 reg_file_reg_22__6_ ( .D(n22306), .CLK(clk), .Q(reg_file[2822]) );
  DFFPOSX1 reg_file_reg_22__7_ ( .D(n22305), .CLK(clk), .Q(reg_file[2823]) );
  DFFPOSX1 reg_file_reg_22__8_ ( .D(n22304), .CLK(clk), .Q(reg_file[2824]) );
  DFFPOSX1 reg_file_reg_22__9_ ( .D(n22303), .CLK(clk), .Q(reg_file[2825]) );
  DFFPOSX1 reg_file_reg_22__10_ ( .D(n22302), .CLK(clk), .Q(reg_file[2826]) );
  DFFPOSX1 reg_file_reg_22__11_ ( .D(n22301), .CLK(clk), .Q(reg_file[2827]) );
  DFFPOSX1 reg_file_reg_22__12_ ( .D(n22300), .CLK(clk), .Q(reg_file[2828]) );
  DFFPOSX1 reg_file_reg_22__13_ ( .D(n22299), .CLK(clk), .Q(reg_file[2829]) );
  DFFPOSX1 reg_file_reg_22__14_ ( .D(n22298), .CLK(clk), .Q(reg_file[2830]) );
  DFFPOSX1 reg_file_reg_22__15_ ( .D(n22297), .CLK(clk), .Q(reg_file[2831]) );
  DFFPOSX1 reg_file_reg_22__16_ ( .D(n22296), .CLK(clk), .Q(reg_file[2832]) );
  DFFPOSX1 reg_file_reg_22__17_ ( .D(n22295), .CLK(clk), .Q(reg_file[2833]) );
  DFFPOSX1 reg_file_reg_22__18_ ( .D(n22294), .CLK(clk), .Q(reg_file[2834]) );
  DFFPOSX1 reg_file_reg_22__19_ ( .D(n22293), .CLK(clk), .Q(reg_file[2835]) );
  DFFPOSX1 reg_file_reg_22__20_ ( .D(n22292), .CLK(clk), .Q(reg_file[2836]) );
  DFFPOSX1 reg_file_reg_22__21_ ( .D(n22291), .CLK(clk), .Q(reg_file[2837]) );
  DFFPOSX1 reg_file_reg_22__22_ ( .D(n22290), .CLK(clk), .Q(reg_file[2838]) );
  DFFPOSX1 reg_file_reg_22__23_ ( .D(n22289), .CLK(clk), .Q(reg_file[2839]) );
  DFFPOSX1 reg_file_reg_22__24_ ( .D(n22288), .CLK(clk), .Q(reg_file[2840]) );
  DFFPOSX1 reg_file_reg_22__25_ ( .D(n22287), .CLK(clk), .Q(reg_file[2841]) );
  DFFPOSX1 reg_file_reg_22__26_ ( .D(n22286), .CLK(clk), .Q(reg_file[2842]) );
  DFFPOSX1 reg_file_reg_22__27_ ( .D(n22285), .CLK(clk), .Q(reg_file[2843]) );
  DFFPOSX1 reg_file_reg_22__28_ ( .D(n22284), .CLK(clk), .Q(reg_file[2844]) );
  DFFPOSX1 reg_file_reg_22__29_ ( .D(n22283), .CLK(clk), .Q(reg_file[2845]) );
  DFFPOSX1 reg_file_reg_22__30_ ( .D(n22282), .CLK(clk), .Q(reg_file[2846]) );
  DFFPOSX1 reg_file_reg_22__31_ ( .D(n22281), .CLK(clk), .Q(reg_file[2847]) );
  DFFPOSX1 reg_file_reg_22__32_ ( .D(n22280), .CLK(clk), .Q(reg_file[2848]) );
  DFFPOSX1 reg_file_reg_22__33_ ( .D(n22279), .CLK(clk), .Q(reg_file[2849]) );
  DFFPOSX1 reg_file_reg_22__34_ ( .D(n22278), .CLK(clk), .Q(reg_file[2850]) );
  DFFPOSX1 reg_file_reg_22__35_ ( .D(n22277), .CLK(clk), .Q(reg_file[2851]) );
  DFFPOSX1 reg_file_reg_22__36_ ( .D(n22276), .CLK(clk), .Q(reg_file[2852]) );
  DFFPOSX1 reg_file_reg_22__37_ ( .D(n22275), .CLK(clk), .Q(reg_file[2853]) );
  DFFPOSX1 reg_file_reg_22__38_ ( .D(n22274), .CLK(clk), .Q(reg_file[2854]) );
  DFFPOSX1 reg_file_reg_22__39_ ( .D(n22273), .CLK(clk), .Q(reg_file[2855]) );
  DFFPOSX1 reg_file_reg_22__40_ ( .D(n22272), .CLK(clk), .Q(reg_file[2856]) );
  DFFPOSX1 reg_file_reg_22__41_ ( .D(n22271), .CLK(clk), .Q(reg_file[2857]) );
  DFFPOSX1 reg_file_reg_22__42_ ( .D(n22270), .CLK(clk), .Q(reg_file[2858]) );
  DFFPOSX1 reg_file_reg_22__43_ ( .D(n22269), .CLK(clk), .Q(reg_file[2859]) );
  DFFPOSX1 reg_file_reg_22__44_ ( .D(n22268), .CLK(clk), .Q(reg_file[2860]) );
  DFFPOSX1 reg_file_reg_22__45_ ( .D(n22267), .CLK(clk), .Q(reg_file[2861]) );
  DFFPOSX1 reg_file_reg_22__46_ ( .D(n22266), .CLK(clk), .Q(reg_file[2862]) );
  DFFPOSX1 reg_file_reg_22__47_ ( .D(n22265), .CLK(clk), .Q(reg_file[2863]) );
  DFFPOSX1 reg_file_reg_22__48_ ( .D(n22264), .CLK(clk), .Q(reg_file[2864]) );
  DFFPOSX1 reg_file_reg_22__49_ ( .D(n22263), .CLK(clk), .Q(reg_file[2865]) );
  DFFPOSX1 reg_file_reg_22__50_ ( .D(n22262), .CLK(clk), .Q(reg_file[2866]) );
  DFFPOSX1 reg_file_reg_22__51_ ( .D(n22261), .CLK(clk), .Q(reg_file[2867]) );
  DFFPOSX1 reg_file_reg_22__52_ ( .D(n22260), .CLK(clk), .Q(reg_file[2868]) );
  DFFPOSX1 reg_file_reg_22__53_ ( .D(n22259), .CLK(clk), .Q(reg_file[2869]) );
  DFFPOSX1 reg_file_reg_22__54_ ( .D(n22258), .CLK(clk), .Q(reg_file[2870]) );
  DFFPOSX1 reg_file_reg_22__55_ ( .D(n22257), .CLK(clk), .Q(reg_file[2871]) );
  DFFPOSX1 reg_file_reg_22__56_ ( .D(n22256), .CLK(clk), .Q(reg_file[2872]) );
  DFFPOSX1 reg_file_reg_22__57_ ( .D(n22255), .CLK(clk), .Q(reg_file[2873]) );
  DFFPOSX1 reg_file_reg_22__58_ ( .D(n22254), .CLK(clk), .Q(reg_file[2874]) );
  DFFPOSX1 reg_file_reg_22__59_ ( .D(n22253), .CLK(clk), .Q(reg_file[2875]) );
  DFFPOSX1 reg_file_reg_22__60_ ( .D(n22252), .CLK(clk), .Q(reg_file[2876]) );
  DFFPOSX1 reg_file_reg_22__61_ ( .D(n22251), .CLK(clk), .Q(reg_file[2877]) );
  DFFPOSX1 reg_file_reg_22__62_ ( .D(n22250), .CLK(clk), .Q(reg_file[2878]) );
  DFFPOSX1 reg_file_reg_22__63_ ( .D(n22249), .CLK(clk), .Q(reg_file[2879]) );
  DFFPOSX1 reg_file_reg_22__64_ ( .D(n22248), .CLK(clk), .Q(reg_file[2880]) );
  DFFPOSX1 reg_file_reg_22__65_ ( .D(n22247), .CLK(clk), .Q(reg_file[2881]) );
  DFFPOSX1 reg_file_reg_22__66_ ( .D(n22246), .CLK(clk), .Q(reg_file[2882]) );
  DFFPOSX1 reg_file_reg_22__67_ ( .D(n22245), .CLK(clk), .Q(reg_file[2883]) );
  DFFPOSX1 reg_file_reg_22__68_ ( .D(n22244), .CLK(clk), .Q(reg_file[2884]) );
  DFFPOSX1 reg_file_reg_22__69_ ( .D(n22243), .CLK(clk), .Q(reg_file[2885]) );
  DFFPOSX1 reg_file_reg_22__70_ ( .D(n22242), .CLK(clk), .Q(reg_file[2886]) );
  DFFPOSX1 reg_file_reg_22__71_ ( .D(n22241), .CLK(clk), .Q(reg_file[2887]) );
  DFFPOSX1 reg_file_reg_22__72_ ( .D(n22240), .CLK(clk), .Q(reg_file[2888]) );
  DFFPOSX1 reg_file_reg_22__73_ ( .D(n22239), .CLK(clk), .Q(reg_file[2889]) );
  DFFPOSX1 reg_file_reg_22__74_ ( .D(n22238), .CLK(clk), .Q(reg_file[2890]) );
  DFFPOSX1 reg_file_reg_22__75_ ( .D(n22237), .CLK(clk), .Q(reg_file[2891]) );
  DFFPOSX1 reg_file_reg_22__76_ ( .D(n22236), .CLK(clk), .Q(reg_file[2892]) );
  DFFPOSX1 reg_file_reg_22__77_ ( .D(n22235), .CLK(clk), .Q(reg_file[2893]) );
  DFFPOSX1 reg_file_reg_22__78_ ( .D(n22234), .CLK(clk), .Q(reg_file[2894]) );
  DFFPOSX1 reg_file_reg_22__79_ ( .D(n22233), .CLK(clk), .Q(reg_file[2895]) );
  DFFPOSX1 reg_file_reg_22__80_ ( .D(n22232), .CLK(clk), .Q(reg_file[2896]) );
  DFFPOSX1 reg_file_reg_22__81_ ( .D(n22231), .CLK(clk), .Q(reg_file[2897]) );
  DFFPOSX1 reg_file_reg_22__82_ ( .D(n22230), .CLK(clk), .Q(reg_file[2898]) );
  DFFPOSX1 reg_file_reg_22__83_ ( .D(n22229), .CLK(clk), .Q(reg_file[2899]) );
  DFFPOSX1 reg_file_reg_22__84_ ( .D(n22228), .CLK(clk), .Q(reg_file[2900]) );
  DFFPOSX1 reg_file_reg_22__85_ ( .D(n22227), .CLK(clk), .Q(reg_file[2901]) );
  DFFPOSX1 reg_file_reg_22__86_ ( .D(n22226), .CLK(clk), .Q(reg_file[2902]) );
  DFFPOSX1 reg_file_reg_22__87_ ( .D(n22225), .CLK(clk), .Q(reg_file[2903]) );
  DFFPOSX1 reg_file_reg_22__88_ ( .D(n22224), .CLK(clk), .Q(reg_file[2904]) );
  DFFPOSX1 reg_file_reg_22__89_ ( .D(n22223), .CLK(clk), .Q(reg_file[2905]) );
  DFFPOSX1 reg_file_reg_22__90_ ( .D(n22222), .CLK(clk), .Q(reg_file[2906]) );
  DFFPOSX1 reg_file_reg_22__91_ ( .D(n22221), .CLK(clk), .Q(reg_file[2907]) );
  DFFPOSX1 reg_file_reg_22__92_ ( .D(n22220), .CLK(clk), .Q(reg_file[2908]) );
  DFFPOSX1 reg_file_reg_22__93_ ( .D(n22219), .CLK(clk), .Q(reg_file[2909]) );
  DFFPOSX1 reg_file_reg_22__94_ ( .D(n22218), .CLK(clk), .Q(reg_file[2910]) );
  DFFPOSX1 reg_file_reg_22__95_ ( .D(n22217), .CLK(clk), .Q(reg_file[2911]) );
  DFFPOSX1 reg_file_reg_22__96_ ( .D(n22216), .CLK(clk), .Q(reg_file[2912]) );
  DFFPOSX1 reg_file_reg_22__97_ ( .D(n22215), .CLK(clk), .Q(reg_file[2913]) );
  DFFPOSX1 reg_file_reg_22__98_ ( .D(n22214), .CLK(clk), .Q(reg_file[2914]) );
  DFFPOSX1 reg_file_reg_22__99_ ( .D(n22213), .CLK(clk), .Q(reg_file[2915]) );
  DFFPOSX1 reg_file_reg_22__100_ ( .D(n22212), .CLK(clk), .Q(reg_file[2916])
         );
  DFFPOSX1 reg_file_reg_22__101_ ( .D(n22211), .CLK(clk), .Q(reg_file[2917])
         );
  DFFPOSX1 reg_file_reg_22__102_ ( .D(n22210), .CLK(clk), .Q(reg_file[2918])
         );
  DFFPOSX1 reg_file_reg_22__103_ ( .D(n22209), .CLK(clk), .Q(reg_file[2919])
         );
  DFFPOSX1 reg_file_reg_22__104_ ( .D(n22208), .CLK(clk), .Q(reg_file[2920])
         );
  DFFPOSX1 reg_file_reg_22__105_ ( .D(n22207), .CLK(clk), .Q(reg_file[2921])
         );
  DFFPOSX1 reg_file_reg_22__106_ ( .D(n22206), .CLK(clk), .Q(reg_file[2922])
         );
  DFFPOSX1 reg_file_reg_22__107_ ( .D(n22205), .CLK(clk), .Q(reg_file[2923])
         );
  DFFPOSX1 reg_file_reg_22__108_ ( .D(n22204), .CLK(clk), .Q(reg_file[2924])
         );
  DFFPOSX1 reg_file_reg_22__109_ ( .D(n22203), .CLK(clk), .Q(reg_file[2925])
         );
  DFFPOSX1 reg_file_reg_22__110_ ( .D(n22202), .CLK(clk), .Q(reg_file[2926])
         );
  DFFPOSX1 reg_file_reg_22__111_ ( .D(n22201), .CLK(clk), .Q(reg_file[2927])
         );
  DFFPOSX1 reg_file_reg_22__112_ ( .D(n22200), .CLK(clk), .Q(reg_file[2928])
         );
  DFFPOSX1 reg_file_reg_22__113_ ( .D(n22199), .CLK(clk), .Q(reg_file[2929])
         );
  DFFPOSX1 reg_file_reg_22__114_ ( .D(n22198), .CLK(clk), .Q(reg_file[2930])
         );
  DFFPOSX1 reg_file_reg_22__115_ ( .D(n22197), .CLK(clk), .Q(reg_file[2931])
         );
  DFFPOSX1 reg_file_reg_22__116_ ( .D(n22196), .CLK(clk), .Q(reg_file[2932])
         );
  DFFPOSX1 reg_file_reg_22__117_ ( .D(n22195), .CLK(clk), .Q(reg_file[2933])
         );
  DFFPOSX1 reg_file_reg_22__118_ ( .D(n22194), .CLK(clk), .Q(reg_file[2934])
         );
  DFFPOSX1 reg_file_reg_22__119_ ( .D(n22193), .CLK(clk), .Q(reg_file[2935])
         );
  DFFPOSX1 reg_file_reg_22__120_ ( .D(n22192), .CLK(clk), .Q(reg_file[2936])
         );
  DFFPOSX1 reg_file_reg_22__121_ ( .D(n22191), .CLK(clk), .Q(reg_file[2937])
         );
  DFFPOSX1 reg_file_reg_22__122_ ( .D(n22190), .CLK(clk), .Q(reg_file[2938])
         );
  DFFPOSX1 reg_file_reg_22__123_ ( .D(n22189), .CLK(clk), .Q(reg_file[2939])
         );
  DFFPOSX1 reg_file_reg_22__124_ ( .D(n22188), .CLK(clk), .Q(reg_file[2940])
         );
  DFFPOSX1 reg_file_reg_22__125_ ( .D(n22187), .CLK(clk), .Q(reg_file[2941])
         );
  DFFPOSX1 reg_file_reg_22__126_ ( .D(n22186), .CLK(clk), .Q(reg_file[2942])
         );
  DFFPOSX1 reg_file_reg_22__127_ ( .D(n22185), .CLK(clk), .Q(reg_file[2943])
         );
  DFFPOSX1 reg_file_reg_23__0_ ( .D(n22184), .CLK(clk), .Q(reg_file[2944]) );
  DFFPOSX1 reg_file_reg_23__1_ ( .D(n22183), .CLK(clk), .Q(reg_file[2945]) );
  DFFPOSX1 reg_file_reg_23__2_ ( .D(n22182), .CLK(clk), .Q(reg_file[2946]) );
  DFFPOSX1 reg_file_reg_23__3_ ( .D(n22181), .CLK(clk), .Q(reg_file[2947]) );
  DFFPOSX1 reg_file_reg_23__4_ ( .D(n22180), .CLK(clk), .Q(reg_file[2948]) );
  DFFPOSX1 reg_file_reg_23__5_ ( .D(n22179), .CLK(clk), .Q(reg_file[2949]) );
  DFFPOSX1 reg_file_reg_23__6_ ( .D(n22178), .CLK(clk), .Q(reg_file[2950]) );
  DFFPOSX1 reg_file_reg_23__7_ ( .D(n22177), .CLK(clk), .Q(reg_file[2951]) );
  DFFPOSX1 reg_file_reg_23__8_ ( .D(n22176), .CLK(clk), .Q(reg_file[2952]) );
  DFFPOSX1 reg_file_reg_23__9_ ( .D(n22175), .CLK(clk), .Q(reg_file[2953]) );
  DFFPOSX1 reg_file_reg_23__10_ ( .D(n22174), .CLK(clk), .Q(reg_file[2954]) );
  DFFPOSX1 reg_file_reg_23__11_ ( .D(n22173), .CLK(clk), .Q(reg_file[2955]) );
  DFFPOSX1 reg_file_reg_23__12_ ( .D(n22172), .CLK(clk), .Q(reg_file[2956]) );
  DFFPOSX1 reg_file_reg_23__13_ ( .D(n22171), .CLK(clk), .Q(reg_file[2957]) );
  DFFPOSX1 reg_file_reg_23__14_ ( .D(n22170), .CLK(clk), .Q(reg_file[2958]) );
  DFFPOSX1 reg_file_reg_23__15_ ( .D(n22169), .CLK(clk), .Q(reg_file[2959]) );
  DFFPOSX1 reg_file_reg_23__16_ ( .D(n22168), .CLK(clk), .Q(reg_file[2960]) );
  DFFPOSX1 reg_file_reg_23__17_ ( .D(n22167), .CLK(clk), .Q(reg_file[2961]) );
  DFFPOSX1 reg_file_reg_23__18_ ( .D(n22166), .CLK(clk), .Q(reg_file[2962]) );
  DFFPOSX1 reg_file_reg_23__19_ ( .D(n22165), .CLK(clk), .Q(reg_file[2963]) );
  DFFPOSX1 reg_file_reg_23__20_ ( .D(n22164), .CLK(clk), .Q(reg_file[2964]) );
  DFFPOSX1 reg_file_reg_23__21_ ( .D(n22163), .CLK(clk), .Q(reg_file[2965]) );
  DFFPOSX1 reg_file_reg_23__22_ ( .D(n22162), .CLK(clk), .Q(reg_file[2966]) );
  DFFPOSX1 reg_file_reg_23__23_ ( .D(n22161), .CLK(clk), .Q(reg_file[2967]) );
  DFFPOSX1 reg_file_reg_23__24_ ( .D(n22160), .CLK(clk), .Q(reg_file[2968]) );
  DFFPOSX1 reg_file_reg_23__25_ ( .D(n22159), .CLK(clk), .Q(reg_file[2969]) );
  DFFPOSX1 reg_file_reg_23__26_ ( .D(n22158), .CLK(clk), .Q(reg_file[2970]) );
  DFFPOSX1 reg_file_reg_23__27_ ( .D(n22157), .CLK(clk), .Q(reg_file[2971]) );
  DFFPOSX1 reg_file_reg_23__28_ ( .D(n22156), .CLK(clk), .Q(reg_file[2972]) );
  DFFPOSX1 reg_file_reg_23__29_ ( .D(n22155), .CLK(clk), .Q(reg_file[2973]) );
  DFFPOSX1 reg_file_reg_23__30_ ( .D(n22154), .CLK(clk), .Q(reg_file[2974]) );
  DFFPOSX1 reg_file_reg_23__31_ ( .D(n22153), .CLK(clk), .Q(reg_file[2975]) );
  DFFPOSX1 reg_file_reg_23__32_ ( .D(n22152), .CLK(clk), .Q(reg_file[2976]) );
  DFFPOSX1 reg_file_reg_23__33_ ( .D(n22151), .CLK(clk), .Q(reg_file[2977]) );
  DFFPOSX1 reg_file_reg_23__34_ ( .D(n22150), .CLK(clk), .Q(reg_file[2978]) );
  DFFPOSX1 reg_file_reg_23__35_ ( .D(n22149), .CLK(clk), .Q(reg_file[2979]) );
  DFFPOSX1 reg_file_reg_23__36_ ( .D(n22148), .CLK(clk), .Q(reg_file[2980]) );
  DFFPOSX1 reg_file_reg_23__37_ ( .D(n22147), .CLK(clk), .Q(reg_file[2981]) );
  DFFPOSX1 reg_file_reg_23__38_ ( .D(n22146), .CLK(clk), .Q(reg_file[2982]) );
  DFFPOSX1 reg_file_reg_23__39_ ( .D(n22145), .CLK(clk), .Q(reg_file[2983]) );
  DFFPOSX1 reg_file_reg_23__40_ ( .D(n22144), .CLK(clk), .Q(reg_file[2984]) );
  DFFPOSX1 reg_file_reg_23__41_ ( .D(n22143), .CLK(clk), .Q(reg_file[2985]) );
  DFFPOSX1 reg_file_reg_23__42_ ( .D(n22142), .CLK(clk), .Q(reg_file[2986]) );
  DFFPOSX1 reg_file_reg_23__43_ ( .D(n22141), .CLK(clk), .Q(reg_file[2987]) );
  DFFPOSX1 reg_file_reg_23__44_ ( .D(n22140), .CLK(clk), .Q(reg_file[2988]) );
  DFFPOSX1 reg_file_reg_23__45_ ( .D(n22139), .CLK(clk), .Q(reg_file[2989]) );
  DFFPOSX1 reg_file_reg_23__46_ ( .D(n22138), .CLK(clk), .Q(reg_file[2990]) );
  DFFPOSX1 reg_file_reg_23__47_ ( .D(n22137), .CLK(clk), .Q(reg_file[2991]) );
  DFFPOSX1 reg_file_reg_23__48_ ( .D(n22136), .CLK(clk), .Q(reg_file[2992]) );
  DFFPOSX1 reg_file_reg_23__49_ ( .D(n22135), .CLK(clk), .Q(reg_file[2993]) );
  DFFPOSX1 reg_file_reg_23__50_ ( .D(n22134), .CLK(clk), .Q(reg_file[2994]) );
  DFFPOSX1 reg_file_reg_23__51_ ( .D(n22133), .CLK(clk), .Q(reg_file[2995]) );
  DFFPOSX1 reg_file_reg_23__52_ ( .D(n22132), .CLK(clk), .Q(reg_file[2996]) );
  DFFPOSX1 reg_file_reg_23__53_ ( .D(n22131), .CLK(clk), .Q(reg_file[2997]) );
  DFFPOSX1 reg_file_reg_23__54_ ( .D(n22130), .CLK(clk), .Q(reg_file[2998]) );
  DFFPOSX1 reg_file_reg_23__55_ ( .D(n22129), .CLK(clk), .Q(reg_file[2999]) );
  DFFPOSX1 reg_file_reg_23__56_ ( .D(n22128), .CLK(clk), .Q(reg_file[3000]) );
  DFFPOSX1 reg_file_reg_23__57_ ( .D(n22127), .CLK(clk), .Q(reg_file[3001]) );
  DFFPOSX1 reg_file_reg_23__58_ ( .D(n22126), .CLK(clk), .Q(reg_file[3002]) );
  DFFPOSX1 reg_file_reg_23__59_ ( .D(n22125), .CLK(clk), .Q(reg_file[3003]) );
  DFFPOSX1 reg_file_reg_23__60_ ( .D(n22124), .CLK(clk), .Q(reg_file[3004]) );
  DFFPOSX1 reg_file_reg_23__61_ ( .D(n22123), .CLK(clk), .Q(reg_file[3005]) );
  DFFPOSX1 reg_file_reg_23__62_ ( .D(n22122), .CLK(clk), .Q(reg_file[3006]) );
  DFFPOSX1 reg_file_reg_23__63_ ( .D(n22121), .CLK(clk), .Q(reg_file[3007]) );
  DFFPOSX1 reg_file_reg_23__64_ ( .D(n22120), .CLK(clk), .Q(reg_file[3008]) );
  DFFPOSX1 reg_file_reg_23__65_ ( .D(n22119), .CLK(clk), .Q(reg_file[3009]) );
  DFFPOSX1 reg_file_reg_23__66_ ( .D(n22118), .CLK(clk), .Q(reg_file[3010]) );
  DFFPOSX1 reg_file_reg_23__67_ ( .D(n22117), .CLK(clk), .Q(reg_file[3011]) );
  DFFPOSX1 reg_file_reg_23__68_ ( .D(n22116), .CLK(clk), .Q(reg_file[3012]) );
  DFFPOSX1 reg_file_reg_23__69_ ( .D(n22115), .CLK(clk), .Q(reg_file[3013]) );
  DFFPOSX1 reg_file_reg_23__70_ ( .D(n22114), .CLK(clk), .Q(reg_file[3014]) );
  DFFPOSX1 reg_file_reg_23__71_ ( .D(n22113), .CLK(clk), .Q(reg_file[3015]) );
  DFFPOSX1 reg_file_reg_23__72_ ( .D(n22112), .CLK(clk), .Q(reg_file[3016]) );
  DFFPOSX1 reg_file_reg_23__73_ ( .D(n22111), .CLK(clk), .Q(reg_file[3017]) );
  DFFPOSX1 reg_file_reg_23__74_ ( .D(n22110), .CLK(clk), .Q(reg_file[3018]) );
  DFFPOSX1 reg_file_reg_23__75_ ( .D(n22109), .CLK(clk), .Q(reg_file[3019]) );
  DFFPOSX1 reg_file_reg_23__76_ ( .D(n22108), .CLK(clk), .Q(reg_file[3020]) );
  DFFPOSX1 reg_file_reg_23__77_ ( .D(n22107), .CLK(clk), .Q(reg_file[3021]) );
  DFFPOSX1 reg_file_reg_23__78_ ( .D(n22106), .CLK(clk), .Q(reg_file[3022]) );
  DFFPOSX1 reg_file_reg_23__79_ ( .D(n22105), .CLK(clk), .Q(reg_file[3023]) );
  DFFPOSX1 reg_file_reg_23__80_ ( .D(n22104), .CLK(clk), .Q(reg_file[3024]) );
  DFFPOSX1 reg_file_reg_23__81_ ( .D(n22103), .CLK(clk), .Q(reg_file[3025]) );
  DFFPOSX1 reg_file_reg_23__82_ ( .D(n22102), .CLK(clk), .Q(reg_file[3026]) );
  DFFPOSX1 reg_file_reg_23__83_ ( .D(n22101), .CLK(clk), .Q(reg_file[3027]) );
  DFFPOSX1 reg_file_reg_23__84_ ( .D(n22100), .CLK(clk), .Q(reg_file[3028]) );
  DFFPOSX1 reg_file_reg_23__85_ ( .D(n22099), .CLK(clk), .Q(reg_file[3029]) );
  DFFPOSX1 reg_file_reg_23__86_ ( .D(n22098), .CLK(clk), .Q(reg_file[3030]) );
  DFFPOSX1 reg_file_reg_23__87_ ( .D(n22097), .CLK(clk), .Q(reg_file[3031]) );
  DFFPOSX1 reg_file_reg_23__88_ ( .D(n22096), .CLK(clk), .Q(reg_file[3032]) );
  DFFPOSX1 reg_file_reg_23__89_ ( .D(n22095), .CLK(clk), .Q(reg_file[3033]) );
  DFFPOSX1 reg_file_reg_23__90_ ( .D(n22094), .CLK(clk), .Q(reg_file[3034]) );
  DFFPOSX1 reg_file_reg_23__91_ ( .D(n22093), .CLK(clk), .Q(reg_file[3035]) );
  DFFPOSX1 reg_file_reg_23__92_ ( .D(n22092), .CLK(clk), .Q(reg_file[3036]) );
  DFFPOSX1 reg_file_reg_23__93_ ( .D(n22091), .CLK(clk), .Q(reg_file[3037]) );
  DFFPOSX1 reg_file_reg_23__94_ ( .D(n22090), .CLK(clk), .Q(reg_file[3038]) );
  DFFPOSX1 reg_file_reg_23__95_ ( .D(n22089), .CLK(clk), .Q(reg_file[3039]) );
  DFFPOSX1 reg_file_reg_23__96_ ( .D(n22088), .CLK(clk), .Q(reg_file[3040]) );
  DFFPOSX1 reg_file_reg_23__97_ ( .D(n22087), .CLK(clk), .Q(reg_file[3041]) );
  DFFPOSX1 reg_file_reg_23__98_ ( .D(n22086), .CLK(clk), .Q(reg_file[3042]) );
  DFFPOSX1 reg_file_reg_23__99_ ( .D(n22085), .CLK(clk), .Q(reg_file[3043]) );
  DFFPOSX1 reg_file_reg_23__100_ ( .D(n22084), .CLK(clk), .Q(reg_file[3044])
         );
  DFFPOSX1 reg_file_reg_23__101_ ( .D(n22083), .CLK(clk), .Q(reg_file[3045])
         );
  DFFPOSX1 reg_file_reg_23__102_ ( .D(n22082), .CLK(clk), .Q(reg_file[3046])
         );
  DFFPOSX1 reg_file_reg_23__103_ ( .D(n22081), .CLK(clk), .Q(reg_file[3047])
         );
  DFFPOSX1 reg_file_reg_23__104_ ( .D(n22080), .CLK(clk), .Q(reg_file[3048])
         );
  DFFPOSX1 reg_file_reg_23__105_ ( .D(n22079), .CLK(clk), .Q(reg_file[3049])
         );
  DFFPOSX1 reg_file_reg_23__106_ ( .D(n22078), .CLK(clk), .Q(reg_file[3050])
         );
  DFFPOSX1 reg_file_reg_23__107_ ( .D(n22077), .CLK(clk), .Q(reg_file[3051])
         );
  DFFPOSX1 reg_file_reg_23__108_ ( .D(n22076), .CLK(clk), .Q(reg_file[3052])
         );
  DFFPOSX1 reg_file_reg_23__109_ ( .D(n22075), .CLK(clk), .Q(reg_file[3053])
         );
  DFFPOSX1 reg_file_reg_23__110_ ( .D(n22074), .CLK(clk), .Q(reg_file[3054])
         );
  DFFPOSX1 reg_file_reg_23__111_ ( .D(n22073), .CLK(clk), .Q(reg_file[3055])
         );
  DFFPOSX1 reg_file_reg_23__112_ ( .D(n22072), .CLK(clk), .Q(reg_file[3056])
         );
  DFFPOSX1 reg_file_reg_23__113_ ( .D(n22071), .CLK(clk), .Q(reg_file[3057])
         );
  DFFPOSX1 reg_file_reg_23__114_ ( .D(n22070), .CLK(clk), .Q(reg_file[3058])
         );
  DFFPOSX1 reg_file_reg_23__115_ ( .D(n22069), .CLK(clk), .Q(reg_file[3059])
         );
  DFFPOSX1 reg_file_reg_23__116_ ( .D(n22068), .CLK(clk), .Q(reg_file[3060])
         );
  DFFPOSX1 reg_file_reg_23__117_ ( .D(n22067), .CLK(clk), .Q(reg_file[3061])
         );
  DFFPOSX1 reg_file_reg_23__118_ ( .D(n22066), .CLK(clk), .Q(reg_file[3062])
         );
  DFFPOSX1 reg_file_reg_23__119_ ( .D(n22065), .CLK(clk), .Q(reg_file[3063])
         );
  DFFPOSX1 reg_file_reg_23__120_ ( .D(n22064), .CLK(clk), .Q(reg_file[3064])
         );
  DFFPOSX1 reg_file_reg_23__121_ ( .D(n22063), .CLK(clk), .Q(reg_file[3065])
         );
  DFFPOSX1 reg_file_reg_23__122_ ( .D(n22062), .CLK(clk), .Q(reg_file[3066])
         );
  DFFPOSX1 reg_file_reg_23__123_ ( .D(n22061), .CLK(clk), .Q(reg_file[3067])
         );
  DFFPOSX1 reg_file_reg_23__124_ ( .D(n22060), .CLK(clk), .Q(reg_file[3068])
         );
  DFFPOSX1 reg_file_reg_23__125_ ( .D(n22059), .CLK(clk), .Q(reg_file[3069])
         );
  DFFPOSX1 reg_file_reg_23__126_ ( .D(n22058), .CLK(clk), .Q(reg_file[3070])
         );
  DFFPOSX1 reg_file_reg_23__127_ ( .D(n22057), .CLK(clk), .Q(reg_file[3071])
         );
  DFFPOSX1 reg_file_reg_24__0_ ( .D(n22056), .CLK(clk), .Q(reg_file[3072]) );
  DFFPOSX1 reg_file_reg_24__1_ ( .D(n22055), .CLK(clk), .Q(reg_file[3073]) );
  DFFPOSX1 reg_file_reg_24__2_ ( .D(n22054), .CLK(clk), .Q(reg_file[3074]) );
  DFFPOSX1 reg_file_reg_24__3_ ( .D(n22053), .CLK(clk), .Q(reg_file[3075]) );
  DFFPOSX1 reg_file_reg_24__4_ ( .D(n22052), .CLK(clk), .Q(reg_file[3076]) );
  DFFPOSX1 reg_file_reg_24__5_ ( .D(n22051), .CLK(clk), .Q(reg_file[3077]) );
  DFFPOSX1 reg_file_reg_24__6_ ( .D(n22050), .CLK(clk), .Q(reg_file[3078]) );
  DFFPOSX1 reg_file_reg_24__7_ ( .D(n22049), .CLK(clk), .Q(reg_file[3079]) );
  DFFPOSX1 reg_file_reg_24__8_ ( .D(n22048), .CLK(clk), .Q(reg_file[3080]) );
  DFFPOSX1 reg_file_reg_24__9_ ( .D(n22047), .CLK(clk), .Q(reg_file[3081]) );
  DFFPOSX1 reg_file_reg_24__10_ ( .D(n22046), .CLK(clk), .Q(reg_file[3082]) );
  DFFPOSX1 reg_file_reg_24__11_ ( .D(n22045), .CLK(clk), .Q(reg_file[3083]) );
  DFFPOSX1 reg_file_reg_24__12_ ( .D(n22044), .CLK(clk), .Q(reg_file[3084]) );
  DFFPOSX1 reg_file_reg_24__13_ ( .D(n22043), .CLK(clk), .Q(reg_file[3085]) );
  DFFPOSX1 reg_file_reg_24__14_ ( .D(n22042), .CLK(clk), .Q(reg_file[3086]) );
  DFFPOSX1 reg_file_reg_24__15_ ( .D(n22041), .CLK(clk), .Q(reg_file[3087]) );
  DFFPOSX1 reg_file_reg_24__16_ ( .D(n22040), .CLK(clk), .Q(reg_file[3088]) );
  DFFPOSX1 reg_file_reg_24__17_ ( .D(n22039), .CLK(clk), .Q(reg_file[3089]) );
  DFFPOSX1 reg_file_reg_24__18_ ( .D(n22038), .CLK(clk), .Q(reg_file[3090]) );
  DFFPOSX1 reg_file_reg_24__19_ ( .D(n22037), .CLK(clk), .Q(reg_file[3091]) );
  DFFPOSX1 reg_file_reg_24__20_ ( .D(n22036), .CLK(clk), .Q(reg_file[3092]) );
  DFFPOSX1 reg_file_reg_24__21_ ( .D(n22035), .CLK(clk), .Q(reg_file[3093]) );
  DFFPOSX1 reg_file_reg_24__22_ ( .D(n22034), .CLK(clk), .Q(reg_file[3094]) );
  DFFPOSX1 reg_file_reg_24__23_ ( .D(n22033), .CLK(clk), .Q(reg_file[3095]) );
  DFFPOSX1 reg_file_reg_24__24_ ( .D(n22032), .CLK(clk), .Q(reg_file[3096]) );
  DFFPOSX1 reg_file_reg_24__25_ ( .D(n22031), .CLK(clk), .Q(reg_file[3097]) );
  DFFPOSX1 reg_file_reg_24__26_ ( .D(n22030), .CLK(clk), .Q(reg_file[3098]) );
  DFFPOSX1 reg_file_reg_24__27_ ( .D(n22029), .CLK(clk), .Q(reg_file[3099]) );
  DFFPOSX1 reg_file_reg_24__28_ ( .D(n22028), .CLK(clk), .Q(reg_file[3100]) );
  DFFPOSX1 reg_file_reg_24__29_ ( .D(n22027), .CLK(clk), .Q(reg_file[3101]) );
  DFFPOSX1 reg_file_reg_24__30_ ( .D(n22026), .CLK(clk), .Q(reg_file[3102]) );
  DFFPOSX1 reg_file_reg_24__31_ ( .D(n22025), .CLK(clk), .Q(reg_file[3103]) );
  DFFPOSX1 reg_file_reg_24__32_ ( .D(n22024), .CLK(clk), .Q(reg_file[3104]) );
  DFFPOSX1 reg_file_reg_24__33_ ( .D(n22023), .CLK(clk), .Q(reg_file[3105]) );
  DFFPOSX1 reg_file_reg_24__34_ ( .D(n22022), .CLK(clk), .Q(reg_file[3106]) );
  DFFPOSX1 reg_file_reg_24__35_ ( .D(n22021), .CLK(clk), .Q(reg_file[3107]) );
  DFFPOSX1 reg_file_reg_24__36_ ( .D(n22020), .CLK(clk), .Q(reg_file[3108]) );
  DFFPOSX1 reg_file_reg_24__37_ ( .D(n22019), .CLK(clk), .Q(reg_file[3109]) );
  DFFPOSX1 reg_file_reg_24__38_ ( .D(n22018), .CLK(clk), .Q(reg_file[3110]) );
  DFFPOSX1 reg_file_reg_24__39_ ( .D(n22017), .CLK(clk), .Q(reg_file[3111]) );
  DFFPOSX1 reg_file_reg_24__40_ ( .D(n22016), .CLK(clk), .Q(reg_file[3112]) );
  DFFPOSX1 reg_file_reg_24__41_ ( .D(n22015), .CLK(clk), .Q(reg_file[3113]) );
  DFFPOSX1 reg_file_reg_24__42_ ( .D(n22014), .CLK(clk), .Q(reg_file[3114]) );
  DFFPOSX1 reg_file_reg_24__43_ ( .D(n22013), .CLK(clk), .Q(reg_file[3115]) );
  DFFPOSX1 reg_file_reg_24__44_ ( .D(n22012), .CLK(clk), .Q(reg_file[3116]) );
  DFFPOSX1 reg_file_reg_24__45_ ( .D(n22011), .CLK(clk), .Q(reg_file[3117]) );
  DFFPOSX1 reg_file_reg_24__46_ ( .D(n22010), .CLK(clk), .Q(reg_file[3118]) );
  DFFPOSX1 reg_file_reg_24__47_ ( .D(n22009), .CLK(clk), .Q(reg_file[3119]) );
  DFFPOSX1 reg_file_reg_24__48_ ( .D(n22008), .CLK(clk), .Q(reg_file[3120]) );
  DFFPOSX1 reg_file_reg_24__49_ ( .D(n22007), .CLK(clk), .Q(reg_file[3121]) );
  DFFPOSX1 reg_file_reg_24__50_ ( .D(n22006), .CLK(clk), .Q(reg_file[3122]) );
  DFFPOSX1 reg_file_reg_24__51_ ( .D(n22005), .CLK(clk), .Q(reg_file[3123]) );
  DFFPOSX1 reg_file_reg_24__52_ ( .D(n22004), .CLK(clk), .Q(reg_file[3124]) );
  DFFPOSX1 reg_file_reg_24__53_ ( .D(n22003), .CLK(clk), .Q(reg_file[3125]) );
  DFFPOSX1 reg_file_reg_24__54_ ( .D(n22002), .CLK(clk), .Q(reg_file[3126]) );
  DFFPOSX1 reg_file_reg_24__55_ ( .D(n22001), .CLK(clk), .Q(reg_file[3127]) );
  DFFPOSX1 reg_file_reg_24__56_ ( .D(n22000), .CLK(clk), .Q(reg_file[3128]) );
  DFFPOSX1 reg_file_reg_24__57_ ( .D(n21999), .CLK(clk), .Q(reg_file[3129]) );
  DFFPOSX1 reg_file_reg_24__58_ ( .D(n21998), .CLK(clk), .Q(reg_file[3130]) );
  DFFPOSX1 reg_file_reg_24__59_ ( .D(n21997), .CLK(clk), .Q(reg_file[3131]) );
  DFFPOSX1 reg_file_reg_24__60_ ( .D(n21996), .CLK(clk), .Q(reg_file[3132]) );
  DFFPOSX1 reg_file_reg_24__61_ ( .D(n21995), .CLK(clk), .Q(reg_file[3133]) );
  DFFPOSX1 reg_file_reg_24__62_ ( .D(n21994), .CLK(clk), .Q(reg_file[3134]) );
  DFFPOSX1 reg_file_reg_24__63_ ( .D(n21993), .CLK(clk), .Q(reg_file[3135]) );
  DFFPOSX1 reg_file_reg_24__64_ ( .D(n21992), .CLK(clk), .Q(reg_file[3136]) );
  DFFPOSX1 reg_file_reg_24__65_ ( .D(n21991), .CLK(clk), .Q(reg_file[3137]) );
  DFFPOSX1 reg_file_reg_24__66_ ( .D(n21990), .CLK(clk), .Q(reg_file[3138]) );
  DFFPOSX1 reg_file_reg_24__67_ ( .D(n21989), .CLK(clk), .Q(reg_file[3139]) );
  DFFPOSX1 reg_file_reg_24__68_ ( .D(n21988), .CLK(clk), .Q(reg_file[3140]) );
  DFFPOSX1 reg_file_reg_24__69_ ( .D(n21987), .CLK(clk), .Q(reg_file[3141]) );
  DFFPOSX1 reg_file_reg_24__70_ ( .D(n21986), .CLK(clk), .Q(reg_file[3142]) );
  DFFPOSX1 reg_file_reg_24__71_ ( .D(n21985), .CLK(clk), .Q(reg_file[3143]) );
  DFFPOSX1 reg_file_reg_24__72_ ( .D(n21984), .CLK(clk), .Q(reg_file[3144]) );
  DFFPOSX1 reg_file_reg_24__73_ ( .D(n21983), .CLK(clk), .Q(reg_file[3145]) );
  DFFPOSX1 reg_file_reg_24__74_ ( .D(n21982), .CLK(clk), .Q(reg_file[3146]) );
  DFFPOSX1 reg_file_reg_24__75_ ( .D(n21981), .CLK(clk), .Q(reg_file[3147]) );
  DFFPOSX1 reg_file_reg_24__76_ ( .D(n21980), .CLK(clk), .Q(reg_file[3148]) );
  DFFPOSX1 reg_file_reg_24__77_ ( .D(n21979), .CLK(clk), .Q(reg_file[3149]) );
  DFFPOSX1 reg_file_reg_24__78_ ( .D(n21978), .CLK(clk), .Q(reg_file[3150]) );
  DFFPOSX1 reg_file_reg_24__79_ ( .D(n21977), .CLK(clk), .Q(reg_file[3151]) );
  DFFPOSX1 reg_file_reg_24__80_ ( .D(n21976), .CLK(clk), .Q(reg_file[3152]) );
  DFFPOSX1 reg_file_reg_24__81_ ( .D(n21975), .CLK(clk), .Q(reg_file[3153]) );
  DFFPOSX1 reg_file_reg_24__82_ ( .D(n21974), .CLK(clk), .Q(reg_file[3154]) );
  DFFPOSX1 reg_file_reg_24__83_ ( .D(n21973), .CLK(clk), .Q(reg_file[3155]) );
  DFFPOSX1 reg_file_reg_24__84_ ( .D(n21972), .CLK(clk), .Q(reg_file[3156]) );
  DFFPOSX1 reg_file_reg_24__85_ ( .D(n21971), .CLK(clk), .Q(reg_file[3157]) );
  DFFPOSX1 reg_file_reg_24__86_ ( .D(n21970), .CLK(clk), .Q(reg_file[3158]) );
  DFFPOSX1 reg_file_reg_24__87_ ( .D(n21969), .CLK(clk), .Q(reg_file[3159]) );
  DFFPOSX1 reg_file_reg_24__88_ ( .D(n21968), .CLK(clk), .Q(reg_file[3160]) );
  DFFPOSX1 reg_file_reg_24__89_ ( .D(n21967), .CLK(clk), .Q(reg_file[3161]) );
  DFFPOSX1 reg_file_reg_24__90_ ( .D(n21966), .CLK(clk), .Q(reg_file[3162]) );
  DFFPOSX1 reg_file_reg_24__91_ ( .D(n21965), .CLK(clk), .Q(reg_file[3163]) );
  DFFPOSX1 reg_file_reg_24__92_ ( .D(n21964), .CLK(clk), .Q(reg_file[3164]) );
  DFFPOSX1 reg_file_reg_24__93_ ( .D(n21963), .CLK(clk), .Q(reg_file[3165]) );
  DFFPOSX1 reg_file_reg_24__94_ ( .D(n21962), .CLK(clk), .Q(reg_file[3166]) );
  DFFPOSX1 reg_file_reg_24__95_ ( .D(n21961), .CLK(clk), .Q(reg_file[3167]) );
  DFFPOSX1 reg_file_reg_24__96_ ( .D(n21960), .CLK(clk), .Q(reg_file[3168]) );
  DFFPOSX1 reg_file_reg_24__97_ ( .D(n21959), .CLK(clk), .Q(reg_file[3169]) );
  DFFPOSX1 reg_file_reg_24__98_ ( .D(n21958), .CLK(clk), .Q(reg_file[3170]) );
  DFFPOSX1 reg_file_reg_24__99_ ( .D(n21957), .CLK(clk), .Q(reg_file[3171]) );
  DFFPOSX1 reg_file_reg_24__100_ ( .D(n21956), .CLK(clk), .Q(reg_file[3172])
         );
  DFFPOSX1 reg_file_reg_24__101_ ( .D(n21955), .CLK(clk), .Q(reg_file[3173])
         );
  DFFPOSX1 reg_file_reg_24__102_ ( .D(n21954), .CLK(clk), .Q(reg_file[3174])
         );
  DFFPOSX1 reg_file_reg_24__103_ ( .D(n21953), .CLK(clk), .Q(reg_file[3175])
         );
  DFFPOSX1 reg_file_reg_24__104_ ( .D(n21952), .CLK(clk), .Q(reg_file[3176])
         );
  DFFPOSX1 reg_file_reg_24__105_ ( .D(n21951), .CLK(clk), .Q(reg_file[3177])
         );
  DFFPOSX1 reg_file_reg_24__106_ ( .D(n21950), .CLK(clk), .Q(reg_file[3178])
         );
  DFFPOSX1 reg_file_reg_24__107_ ( .D(n21949), .CLK(clk), .Q(reg_file[3179])
         );
  DFFPOSX1 reg_file_reg_24__108_ ( .D(n21948), .CLK(clk), .Q(reg_file[3180])
         );
  DFFPOSX1 reg_file_reg_24__109_ ( .D(n21947), .CLK(clk), .Q(reg_file[3181])
         );
  DFFPOSX1 reg_file_reg_24__110_ ( .D(n21946), .CLK(clk), .Q(reg_file[3182])
         );
  DFFPOSX1 reg_file_reg_24__111_ ( .D(n21945), .CLK(clk), .Q(reg_file[3183])
         );
  DFFPOSX1 reg_file_reg_24__112_ ( .D(n21944), .CLK(clk), .Q(reg_file[3184])
         );
  DFFPOSX1 reg_file_reg_24__113_ ( .D(n21943), .CLK(clk), .Q(reg_file[3185])
         );
  DFFPOSX1 reg_file_reg_24__114_ ( .D(n21942), .CLK(clk), .Q(reg_file[3186])
         );
  DFFPOSX1 reg_file_reg_24__115_ ( .D(n21941), .CLK(clk), .Q(reg_file[3187])
         );
  DFFPOSX1 reg_file_reg_24__116_ ( .D(n21940), .CLK(clk), .Q(reg_file[3188])
         );
  DFFPOSX1 reg_file_reg_24__117_ ( .D(n21939), .CLK(clk), .Q(reg_file[3189])
         );
  DFFPOSX1 reg_file_reg_24__118_ ( .D(n21938), .CLK(clk), .Q(reg_file[3190])
         );
  DFFPOSX1 reg_file_reg_24__119_ ( .D(n21937), .CLK(clk), .Q(reg_file[3191])
         );
  DFFPOSX1 reg_file_reg_24__120_ ( .D(n21936), .CLK(clk), .Q(reg_file[3192])
         );
  DFFPOSX1 reg_file_reg_24__121_ ( .D(n21935), .CLK(clk), .Q(reg_file[3193])
         );
  DFFPOSX1 reg_file_reg_24__122_ ( .D(n21934), .CLK(clk), .Q(reg_file[3194])
         );
  DFFPOSX1 reg_file_reg_24__123_ ( .D(n21933), .CLK(clk), .Q(reg_file[3195])
         );
  DFFPOSX1 reg_file_reg_24__124_ ( .D(n21932), .CLK(clk), .Q(reg_file[3196])
         );
  DFFPOSX1 reg_file_reg_24__125_ ( .D(n21931), .CLK(clk), .Q(reg_file[3197])
         );
  DFFPOSX1 reg_file_reg_24__126_ ( .D(n21930), .CLK(clk), .Q(reg_file[3198])
         );
  DFFPOSX1 reg_file_reg_24__127_ ( .D(n21929), .CLK(clk), .Q(reg_file[3199])
         );
  DFFPOSX1 reg_file_reg_25__0_ ( .D(n21928), .CLK(clk), .Q(reg_file[3200]) );
  DFFPOSX1 reg_file_reg_25__1_ ( .D(n21927), .CLK(clk), .Q(reg_file[3201]) );
  DFFPOSX1 reg_file_reg_25__2_ ( .D(n21926), .CLK(clk), .Q(reg_file[3202]) );
  DFFPOSX1 reg_file_reg_25__3_ ( .D(n21925), .CLK(clk), .Q(reg_file[3203]) );
  DFFPOSX1 reg_file_reg_25__4_ ( .D(n21924), .CLK(clk), .Q(reg_file[3204]) );
  DFFPOSX1 reg_file_reg_25__5_ ( .D(n21923), .CLK(clk), .Q(reg_file[3205]) );
  DFFPOSX1 reg_file_reg_25__6_ ( .D(n21922), .CLK(clk), .Q(reg_file[3206]) );
  DFFPOSX1 reg_file_reg_25__7_ ( .D(n21921), .CLK(clk), .Q(reg_file[3207]) );
  DFFPOSX1 reg_file_reg_25__8_ ( .D(n21920), .CLK(clk), .Q(reg_file[3208]) );
  DFFPOSX1 reg_file_reg_25__9_ ( .D(n21919), .CLK(clk), .Q(reg_file[3209]) );
  DFFPOSX1 reg_file_reg_25__10_ ( .D(n21918), .CLK(clk), .Q(reg_file[3210]) );
  DFFPOSX1 reg_file_reg_25__11_ ( .D(n21917), .CLK(clk), .Q(reg_file[3211]) );
  DFFPOSX1 reg_file_reg_25__12_ ( .D(n21916), .CLK(clk), .Q(reg_file[3212]) );
  DFFPOSX1 reg_file_reg_25__13_ ( .D(n21915), .CLK(clk), .Q(reg_file[3213]) );
  DFFPOSX1 reg_file_reg_25__14_ ( .D(n21914), .CLK(clk), .Q(reg_file[3214]) );
  DFFPOSX1 reg_file_reg_25__15_ ( .D(n21913), .CLK(clk), .Q(reg_file[3215]) );
  DFFPOSX1 reg_file_reg_25__16_ ( .D(n21912), .CLK(clk), .Q(reg_file[3216]) );
  DFFPOSX1 reg_file_reg_25__17_ ( .D(n21911), .CLK(clk), .Q(reg_file[3217]) );
  DFFPOSX1 reg_file_reg_25__18_ ( .D(n21910), .CLK(clk), .Q(reg_file[3218]) );
  DFFPOSX1 reg_file_reg_25__19_ ( .D(n21909), .CLK(clk), .Q(reg_file[3219]) );
  DFFPOSX1 reg_file_reg_25__20_ ( .D(n21908), .CLK(clk), .Q(reg_file[3220]) );
  DFFPOSX1 reg_file_reg_25__21_ ( .D(n21907), .CLK(clk), .Q(reg_file[3221]) );
  DFFPOSX1 reg_file_reg_25__22_ ( .D(n21906), .CLK(clk), .Q(reg_file[3222]) );
  DFFPOSX1 reg_file_reg_25__23_ ( .D(n21905), .CLK(clk), .Q(reg_file[3223]) );
  DFFPOSX1 reg_file_reg_25__24_ ( .D(n21904), .CLK(clk), .Q(reg_file[3224]) );
  DFFPOSX1 reg_file_reg_25__25_ ( .D(n21903), .CLK(clk), .Q(reg_file[3225]) );
  DFFPOSX1 reg_file_reg_25__26_ ( .D(n21902), .CLK(clk), .Q(reg_file[3226]) );
  DFFPOSX1 reg_file_reg_25__27_ ( .D(n21901), .CLK(clk), .Q(reg_file[3227]) );
  DFFPOSX1 reg_file_reg_25__28_ ( .D(n21900), .CLK(clk), .Q(reg_file[3228]) );
  DFFPOSX1 reg_file_reg_25__29_ ( .D(n21899), .CLK(clk), .Q(reg_file[3229]) );
  DFFPOSX1 reg_file_reg_25__30_ ( .D(n21898), .CLK(clk), .Q(reg_file[3230]) );
  DFFPOSX1 reg_file_reg_25__31_ ( .D(n21897), .CLK(clk), .Q(reg_file[3231]) );
  DFFPOSX1 reg_file_reg_25__32_ ( .D(n21896), .CLK(clk), .Q(reg_file[3232]) );
  DFFPOSX1 reg_file_reg_25__33_ ( .D(n21895), .CLK(clk), .Q(reg_file[3233]) );
  DFFPOSX1 reg_file_reg_25__34_ ( .D(n21894), .CLK(clk), .Q(reg_file[3234]) );
  DFFPOSX1 reg_file_reg_25__35_ ( .D(n21893), .CLK(clk), .Q(reg_file[3235]) );
  DFFPOSX1 reg_file_reg_25__36_ ( .D(n21892), .CLK(clk), .Q(reg_file[3236]) );
  DFFPOSX1 reg_file_reg_25__37_ ( .D(n21891), .CLK(clk), .Q(reg_file[3237]) );
  DFFPOSX1 reg_file_reg_25__38_ ( .D(n21890), .CLK(clk), .Q(reg_file[3238]) );
  DFFPOSX1 reg_file_reg_25__39_ ( .D(n21889), .CLK(clk), .Q(reg_file[3239]) );
  DFFPOSX1 reg_file_reg_25__40_ ( .D(n21888), .CLK(clk), .Q(reg_file[3240]) );
  DFFPOSX1 reg_file_reg_25__41_ ( .D(n21887), .CLK(clk), .Q(reg_file[3241]) );
  DFFPOSX1 reg_file_reg_25__42_ ( .D(n21886), .CLK(clk), .Q(reg_file[3242]) );
  DFFPOSX1 reg_file_reg_25__43_ ( .D(n21885), .CLK(clk), .Q(reg_file[3243]) );
  DFFPOSX1 reg_file_reg_25__44_ ( .D(n21884), .CLK(clk), .Q(reg_file[3244]) );
  DFFPOSX1 reg_file_reg_25__45_ ( .D(n21883), .CLK(clk), .Q(reg_file[3245]) );
  DFFPOSX1 reg_file_reg_25__46_ ( .D(n21882), .CLK(clk), .Q(reg_file[3246]) );
  DFFPOSX1 reg_file_reg_25__47_ ( .D(n21881), .CLK(clk), .Q(reg_file[3247]) );
  DFFPOSX1 reg_file_reg_25__48_ ( .D(n21880), .CLK(clk), .Q(reg_file[3248]) );
  DFFPOSX1 reg_file_reg_25__49_ ( .D(n21879), .CLK(clk), .Q(reg_file[3249]) );
  DFFPOSX1 reg_file_reg_25__50_ ( .D(n21878), .CLK(clk), .Q(reg_file[3250]) );
  DFFPOSX1 reg_file_reg_25__51_ ( .D(n21877), .CLK(clk), .Q(reg_file[3251]) );
  DFFPOSX1 reg_file_reg_25__52_ ( .D(n21876), .CLK(clk), .Q(reg_file[3252]) );
  DFFPOSX1 reg_file_reg_25__53_ ( .D(n21875), .CLK(clk), .Q(reg_file[3253]) );
  DFFPOSX1 reg_file_reg_25__54_ ( .D(n21874), .CLK(clk), .Q(reg_file[3254]) );
  DFFPOSX1 reg_file_reg_25__55_ ( .D(n21873), .CLK(clk), .Q(reg_file[3255]) );
  DFFPOSX1 reg_file_reg_25__56_ ( .D(n21872), .CLK(clk), .Q(reg_file[3256]) );
  DFFPOSX1 reg_file_reg_25__57_ ( .D(n21871), .CLK(clk), .Q(reg_file[3257]) );
  DFFPOSX1 reg_file_reg_25__58_ ( .D(n21870), .CLK(clk), .Q(reg_file[3258]) );
  DFFPOSX1 reg_file_reg_25__59_ ( .D(n21869), .CLK(clk), .Q(reg_file[3259]) );
  DFFPOSX1 reg_file_reg_25__60_ ( .D(n21868), .CLK(clk), .Q(reg_file[3260]) );
  DFFPOSX1 reg_file_reg_25__61_ ( .D(n21867), .CLK(clk), .Q(reg_file[3261]) );
  DFFPOSX1 reg_file_reg_25__62_ ( .D(n21866), .CLK(clk), .Q(reg_file[3262]) );
  DFFPOSX1 reg_file_reg_25__63_ ( .D(n21865), .CLK(clk), .Q(reg_file[3263]) );
  DFFPOSX1 reg_file_reg_25__64_ ( .D(n21864), .CLK(clk), .Q(reg_file[3264]) );
  DFFPOSX1 reg_file_reg_25__65_ ( .D(n21863), .CLK(clk), .Q(reg_file[3265]) );
  DFFPOSX1 reg_file_reg_25__66_ ( .D(n21862), .CLK(clk), .Q(reg_file[3266]) );
  DFFPOSX1 reg_file_reg_25__67_ ( .D(n21861), .CLK(clk), .Q(reg_file[3267]) );
  DFFPOSX1 reg_file_reg_25__68_ ( .D(n21860), .CLK(clk), .Q(reg_file[3268]) );
  DFFPOSX1 reg_file_reg_25__69_ ( .D(n21859), .CLK(clk), .Q(reg_file[3269]) );
  DFFPOSX1 reg_file_reg_25__70_ ( .D(n21858), .CLK(clk), .Q(reg_file[3270]) );
  DFFPOSX1 reg_file_reg_25__71_ ( .D(n21857), .CLK(clk), .Q(reg_file[3271]) );
  DFFPOSX1 reg_file_reg_25__72_ ( .D(n21856), .CLK(clk), .Q(reg_file[3272]) );
  DFFPOSX1 reg_file_reg_25__73_ ( .D(n21855), .CLK(clk), .Q(reg_file[3273]) );
  DFFPOSX1 reg_file_reg_25__74_ ( .D(n21854), .CLK(clk), .Q(reg_file[3274]) );
  DFFPOSX1 reg_file_reg_25__75_ ( .D(n21853), .CLK(clk), .Q(reg_file[3275]) );
  DFFPOSX1 reg_file_reg_25__76_ ( .D(n21852), .CLK(clk), .Q(reg_file[3276]) );
  DFFPOSX1 reg_file_reg_25__77_ ( .D(n21851), .CLK(clk), .Q(reg_file[3277]) );
  DFFPOSX1 reg_file_reg_25__78_ ( .D(n21850), .CLK(clk), .Q(reg_file[3278]) );
  DFFPOSX1 reg_file_reg_25__79_ ( .D(n21849), .CLK(clk), .Q(reg_file[3279]) );
  DFFPOSX1 reg_file_reg_25__80_ ( .D(n21848), .CLK(clk), .Q(reg_file[3280]) );
  DFFPOSX1 reg_file_reg_25__81_ ( .D(n21847), .CLK(clk), .Q(reg_file[3281]) );
  DFFPOSX1 reg_file_reg_25__82_ ( .D(n21846), .CLK(clk), .Q(reg_file[3282]) );
  DFFPOSX1 reg_file_reg_25__83_ ( .D(n21845), .CLK(clk), .Q(reg_file[3283]) );
  DFFPOSX1 reg_file_reg_25__84_ ( .D(n21844), .CLK(clk), .Q(reg_file[3284]) );
  DFFPOSX1 reg_file_reg_25__85_ ( .D(n21843), .CLK(clk), .Q(reg_file[3285]) );
  DFFPOSX1 reg_file_reg_25__86_ ( .D(n21842), .CLK(clk), .Q(reg_file[3286]) );
  DFFPOSX1 reg_file_reg_25__87_ ( .D(n21841), .CLK(clk), .Q(reg_file[3287]) );
  DFFPOSX1 reg_file_reg_25__88_ ( .D(n21840), .CLK(clk), .Q(reg_file[3288]) );
  DFFPOSX1 reg_file_reg_25__89_ ( .D(n21839), .CLK(clk), .Q(reg_file[3289]) );
  DFFPOSX1 reg_file_reg_25__90_ ( .D(n21838), .CLK(clk), .Q(reg_file[3290]) );
  DFFPOSX1 reg_file_reg_25__91_ ( .D(n21837), .CLK(clk), .Q(reg_file[3291]) );
  DFFPOSX1 reg_file_reg_25__92_ ( .D(n21836), .CLK(clk), .Q(reg_file[3292]) );
  DFFPOSX1 reg_file_reg_25__93_ ( .D(n21835), .CLK(clk), .Q(reg_file[3293]) );
  DFFPOSX1 reg_file_reg_25__94_ ( .D(n21834), .CLK(clk), .Q(reg_file[3294]) );
  DFFPOSX1 reg_file_reg_25__95_ ( .D(n21833), .CLK(clk), .Q(reg_file[3295]) );
  DFFPOSX1 reg_file_reg_25__96_ ( .D(n21832), .CLK(clk), .Q(reg_file[3296]) );
  DFFPOSX1 reg_file_reg_25__97_ ( .D(n21831), .CLK(clk), .Q(reg_file[3297]) );
  DFFPOSX1 reg_file_reg_25__98_ ( .D(n21830), .CLK(clk), .Q(reg_file[3298]) );
  DFFPOSX1 reg_file_reg_25__99_ ( .D(n21829), .CLK(clk), .Q(reg_file[3299]) );
  DFFPOSX1 reg_file_reg_25__100_ ( .D(n21828), .CLK(clk), .Q(reg_file[3300])
         );
  DFFPOSX1 reg_file_reg_25__101_ ( .D(n21827), .CLK(clk), .Q(reg_file[3301])
         );
  DFFPOSX1 reg_file_reg_25__102_ ( .D(n21826), .CLK(clk), .Q(reg_file[3302])
         );
  DFFPOSX1 reg_file_reg_25__103_ ( .D(n21825), .CLK(clk), .Q(reg_file[3303])
         );
  DFFPOSX1 reg_file_reg_25__104_ ( .D(n21824), .CLK(clk), .Q(reg_file[3304])
         );
  DFFPOSX1 reg_file_reg_25__105_ ( .D(n21823), .CLK(clk), .Q(reg_file[3305])
         );
  DFFPOSX1 reg_file_reg_25__106_ ( .D(n21822), .CLK(clk), .Q(reg_file[3306])
         );
  DFFPOSX1 reg_file_reg_25__107_ ( .D(n21821), .CLK(clk), .Q(reg_file[3307])
         );
  DFFPOSX1 reg_file_reg_25__108_ ( .D(n21820), .CLK(clk), .Q(reg_file[3308])
         );
  DFFPOSX1 reg_file_reg_25__109_ ( .D(n21819), .CLK(clk), .Q(reg_file[3309])
         );
  DFFPOSX1 reg_file_reg_25__110_ ( .D(n21818), .CLK(clk), .Q(reg_file[3310])
         );
  DFFPOSX1 reg_file_reg_25__111_ ( .D(n21817), .CLK(clk), .Q(reg_file[3311])
         );
  DFFPOSX1 reg_file_reg_25__112_ ( .D(n21816), .CLK(clk), .Q(reg_file[3312])
         );
  DFFPOSX1 reg_file_reg_25__113_ ( .D(n21815), .CLK(clk), .Q(reg_file[3313])
         );
  DFFPOSX1 reg_file_reg_25__114_ ( .D(n21814), .CLK(clk), .Q(reg_file[3314])
         );
  DFFPOSX1 reg_file_reg_25__115_ ( .D(n21813), .CLK(clk), .Q(reg_file[3315])
         );
  DFFPOSX1 reg_file_reg_25__116_ ( .D(n21812), .CLK(clk), .Q(reg_file[3316])
         );
  DFFPOSX1 reg_file_reg_25__117_ ( .D(n21811), .CLK(clk), .Q(reg_file[3317])
         );
  DFFPOSX1 reg_file_reg_25__118_ ( .D(n21810), .CLK(clk), .Q(reg_file[3318])
         );
  DFFPOSX1 reg_file_reg_25__119_ ( .D(n21809), .CLK(clk), .Q(reg_file[3319])
         );
  DFFPOSX1 reg_file_reg_25__120_ ( .D(n21808), .CLK(clk), .Q(reg_file[3320])
         );
  DFFPOSX1 reg_file_reg_25__121_ ( .D(n21807), .CLK(clk), .Q(reg_file[3321])
         );
  DFFPOSX1 reg_file_reg_25__122_ ( .D(n21806), .CLK(clk), .Q(reg_file[3322])
         );
  DFFPOSX1 reg_file_reg_25__123_ ( .D(n21805), .CLK(clk), .Q(reg_file[3323])
         );
  DFFPOSX1 reg_file_reg_25__124_ ( .D(n21804), .CLK(clk), .Q(reg_file[3324])
         );
  DFFPOSX1 reg_file_reg_25__125_ ( .D(n21803), .CLK(clk), .Q(reg_file[3325])
         );
  DFFPOSX1 reg_file_reg_25__126_ ( .D(n21802), .CLK(clk), .Q(reg_file[3326])
         );
  DFFPOSX1 reg_file_reg_25__127_ ( .D(n21801), .CLK(clk), .Q(reg_file[3327])
         );
  DFFPOSX1 reg_file_reg_26__0_ ( .D(n21800), .CLK(clk), .Q(reg_file[3328]) );
  DFFPOSX1 reg_file_reg_26__1_ ( .D(n21799), .CLK(clk), .Q(reg_file[3329]) );
  DFFPOSX1 reg_file_reg_26__2_ ( .D(n21798), .CLK(clk), .Q(reg_file[3330]) );
  DFFPOSX1 reg_file_reg_26__3_ ( .D(n21797), .CLK(clk), .Q(reg_file[3331]) );
  DFFPOSX1 reg_file_reg_26__4_ ( .D(n21796), .CLK(clk), .Q(reg_file[3332]) );
  DFFPOSX1 reg_file_reg_26__5_ ( .D(n21795), .CLK(clk), .Q(reg_file[3333]) );
  DFFPOSX1 reg_file_reg_26__6_ ( .D(n21794), .CLK(clk), .Q(reg_file[3334]) );
  DFFPOSX1 reg_file_reg_26__7_ ( .D(n21793), .CLK(clk), .Q(reg_file[3335]) );
  DFFPOSX1 reg_file_reg_26__8_ ( .D(n21792), .CLK(clk), .Q(reg_file[3336]) );
  DFFPOSX1 reg_file_reg_26__9_ ( .D(n21791), .CLK(clk), .Q(reg_file[3337]) );
  DFFPOSX1 reg_file_reg_26__10_ ( .D(n21790), .CLK(clk), .Q(reg_file[3338]) );
  DFFPOSX1 reg_file_reg_26__11_ ( .D(n21789), .CLK(clk), .Q(reg_file[3339]) );
  DFFPOSX1 reg_file_reg_26__12_ ( .D(n21788), .CLK(clk), .Q(reg_file[3340]) );
  DFFPOSX1 reg_file_reg_26__13_ ( .D(n21787), .CLK(clk), .Q(reg_file[3341]) );
  DFFPOSX1 reg_file_reg_26__14_ ( .D(n21786), .CLK(clk), .Q(reg_file[3342]) );
  DFFPOSX1 reg_file_reg_26__15_ ( .D(n21785), .CLK(clk), .Q(reg_file[3343]) );
  DFFPOSX1 reg_file_reg_26__16_ ( .D(n21784), .CLK(clk), .Q(reg_file[3344]) );
  DFFPOSX1 reg_file_reg_26__17_ ( .D(n21783), .CLK(clk), .Q(reg_file[3345]) );
  DFFPOSX1 reg_file_reg_26__18_ ( .D(n21782), .CLK(clk), .Q(reg_file[3346]) );
  DFFPOSX1 reg_file_reg_26__19_ ( .D(n21781), .CLK(clk), .Q(reg_file[3347]) );
  DFFPOSX1 reg_file_reg_26__20_ ( .D(n21780), .CLK(clk), .Q(reg_file[3348]) );
  DFFPOSX1 reg_file_reg_26__21_ ( .D(n21779), .CLK(clk), .Q(reg_file[3349]) );
  DFFPOSX1 reg_file_reg_26__22_ ( .D(n21778), .CLK(clk), .Q(reg_file[3350]) );
  DFFPOSX1 reg_file_reg_26__23_ ( .D(n21777), .CLK(clk), .Q(reg_file[3351]) );
  DFFPOSX1 reg_file_reg_26__24_ ( .D(n21776), .CLK(clk), .Q(reg_file[3352]) );
  DFFPOSX1 reg_file_reg_26__25_ ( .D(n21775), .CLK(clk), .Q(reg_file[3353]) );
  DFFPOSX1 reg_file_reg_26__26_ ( .D(n21774), .CLK(clk), .Q(reg_file[3354]) );
  DFFPOSX1 reg_file_reg_26__27_ ( .D(n21773), .CLK(clk), .Q(reg_file[3355]) );
  DFFPOSX1 reg_file_reg_26__28_ ( .D(n21772), .CLK(clk), .Q(reg_file[3356]) );
  DFFPOSX1 reg_file_reg_26__29_ ( .D(n21771), .CLK(clk), .Q(reg_file[3357]) );
  DFFPOSX1 reg_file_reg_26__30_ ( .D(n21770), .CLK(clk), .Q(reg_file[3358]) );
  DFFPOSX1 reg_file_reg_26__31_ ( .D(n21769), .CLK(clk), .Q(reg_file[3359]) );
  DFFPOSX1 reg_file_reg_26__32_ ( .D(n21768), .CLK(clk), .Q(reg_file[3360]) );
  DFFPOSX1 reg_file_reg_26__33_ ( .D(n21767), .CLK(clk), .Q(reg_file[3361]) );
  DFFPOSX1 reg_file_reg_26__34_ ( .D(n21766), .CLK(clk), .Q(reg_file[3362]) );
  DFFPOSX1 reg_file_reg_26__35_ ( .D(n21765), .CLK(clk), .Q(reg_file[3363]) );
  DFFPOSX1 reg_file_reg_26__36_ ( .D(n21764), .CLK(clk), .Q(reg_file[3364]) );
  DFFPOSX1 reg_file_reg_26__37_ ( .D(n21763), .CLK(clk), .Q(reg_file[3365]) );
  DFFPOSX1 reg_file_reg_26__38_ ( .D(n21762), .CLK(clk), .Q(reg_file[3366]) );
  DFFPOSX1 reg_file_reg_26__39_ ( .D(n21761), .CLK(clk), .Q(reg_file[3367]) );
  DFFPOSX1 reg_file_reg_26__40_ ( .D(n21760), .CLK(clk), .Q(reg_file[3368]) );
  DFFPOSX1 reg_file_reg_26__41_ ( .D(n21759), .CLK(clk), .Q(reg_file[3369]) );
  DFFPOSX1 reg_file_reg_26__42_ ( .D(n21758), .CLK(clk), .Q(reg_file[3370]) );
  DFFPOSX1 reg_file_reg_26__43_ ( .D(n21757), .CLK(clk), .Q(reg_file[3371]) );
  DFFPOSX1 reg_file_reg_26__44_ ( .D(n21756), .CLK(clk), .Q(reg_file[3372]) );
  DFFPOSX1 reg_file_reg_26__45_ ( .D(n21755), .CLK(clk), .Q(reg_file[3373]) );
  DFFPOSX1 reg_file_reg_26__46_ ( .D(n21754), .CLK(clk), .Q(reg_file[3374]) );
  DFFPOSX1 reg_file_reg_26__47_ ( .D(n21753), .CLK(clk), .Q(reg_file[3375]) );
  DFFPOSX1 reg_file_reg_26__48_ ( .D(n21752), .CLK(clk), .Q(reg_file[3376]) );
  DFFPOSX1 reg_file_reg_26__49_ ( .D(n21751), .CLK(clk), .Q(reg_file[3377]) );
  DFFPOSX1 reg_file_reg_26__50_ ( .D(n21750), .CLK(clk), .Q(reg_file[3378]) );
  DFFPOSX1 reg_file_reg_26__51_ ( .D(n21749), .CLK(clk), .Q(reg_file[3379]) );
  DFFPOSX1 reg_file_reg_26__52_ ( .D(n21748), .CLK(clk), .Q(reg_file[3380]) );
  DFFPOSX1 reg_file_reg_26__53_ ( .D(n21747), .CLK(clk), .Q(reg_file[3381]) );
  DFFPOSX1 reg_file_reg_26__54_ ( .D(n21746), .CLK(clk), .Q(reg_file[3382]) );
  DFFPOSX1 reg_file_reg_26__55_ ( .D(n21745), .CLK(clk), .Q(reg_file[3383]) );
  DFFPOSX1 reg_file_reg_26__56_ ( .D(n21744), .CLK(clk), .Q(reg_file[3384]) );
  DFFPOSX1 reg_file_reg_26__57_ ( .D(n21743), .CLK(clk), .Q(reg_file[3385]) );
  DFFPOSX1 reg_file_reg_26__58_ ( .D(n21742), .CLK(clk), .Q(reg_file[3386]) );
  DFFPOSX1 reg_file_reg_26__59_ ( .D(n21741), .CLK(clk), .Q(reg_file[3387]) );
  DFFPOSX1 reg_file_reg_26__60_ ( .D(n21740), .CLK(clk), .Q(reg_file[3388]) );
  DFFPOSX1 reg_file_reg_26__61_ ( .D(n21739), .CLK(clk), .Q(reg_file[3389]) );
  DFFPOSX1 reg_file_reg_26__62_ ( .D(n21738), .CLK(clk), .Q(reg_file[3390]) );
  DFFPOSX1 reg_file_reg_26__63_ ( .D(n21737), .CLK(clk), .Q(reg_file[3391]) );
  DFFPOSX1 reg_file_reg_26__64_ ( .D(n21736), .CLK(clk), .Q(reg_file[3392]) );
  DFFPOSX1 reg_file_reg_26__65_ ( .D(n21735), .CLK(clk), .Q(reg_file[3393]) );
  DFFPOSX1 reg_file_reg_26__66_ ( .D(n21734), .CLK(clk), .Q(reg_file[3394]) );
  DFFPOSX1 reg_file_reg_26__67_ ( .D(n21733), .CLK(clk), .Q(reg_file[3395]) );
  DFFPOSX1 reg_file_reg_26__68_ ( .D(n21732), .CLK(clk), .Q(reg_file[3396]) );
  DFFPOSX1 reg_file_reg_26__69_ ( .D(n21731), .CLK(clk), .Q(reg_file[3397]) );
  DFFPOSX1 reg_file_reg_26__70_ ( .D(n21730), .CLK(clk), .Q(reg_file[3398]) );
  DFFPOSX1 reg_file_reg_26__71_ ( .D(n21729), .CLK(clk), .Q(reg_file[3399]) );
  DFFPOSX1 reg_file_reg_26__72_ ( .D(n21728), .CLK(clk), .Q(reg_file[3400]) );
  DFFPOSX1 reg_file_reg_26__73_ ( .D(n21727), .CLK(clk), .Q(reg_file[3401]) );
  DFFPOSX1 reg_file_reg_26__74_ ( .D(n21726), .CLK(clk), .Q(reg_file[3402]) );
  DFFPOSX1 reg_file_reg_26__75_ ( .D(n21725), .CLK(clk), .Q(reg_file[3403]) );
  DFFPOSX1 reg_file_reg_26__76_ ( .D(n21724), .CLK(clk), .Q(reg_file[3404]) );
  DFFPOSX1 reg_file_reg_26__77_ ( .D(n21723), .CLK(clk), .Q(reg_file[3405]) );
  DFFPOSX1 reg_file_reg_26__78_ ( .D(n21722), .CLK(clk), .Q(reg_file[3406]) );
  DFFPOSX1 reg_file_reg_26__79_ ( .D(n21721), .CLK(clk), .Q(reg_file[3407]) );
  DFFPOSX1 reg_file_reg_26__80_ ( .D(n21720), .CLK(clk), .Q(reg_file[3408]) );
  DFFPOSX1 reg_file_reg_26__81_ ( .D(n21719), .CLK(clk), .Q(reg_file[3409]) );
  DFFPOSX1 reg_file_reg_26__82_ ( .D(n21718), .CLK(clk), .Q(reg_file[3410]) );
  DFFPOSX1 reg_file_reg_26__83_ ( .D(n21717), .CLK(clk), .Q(reg_file[3411]) );
  DFFPOSX1 reg_file_reg_26__84_ ( .D(n21716), .CLK(clk), .Q(reg_file[3412]) );
  DFFPOSX1 reg_file_reg_26__85_ ( .D(n21715), .CLK(clk), .Q(reg_file[3413]) );
  DFFPOSX1 reg_file_reg_26__86_ ( .D(n21714), .CLK(clk), .Q(reg_file[3414]) );
  DFFPOSX1 reg_file_reg_26__87_ ( .D(n21713), .CLK(clk), .Q(reg_file[3415]) );
  DFFPOSX1 reg_file_reg_26__88_ ( .D(n21712), .CLK(clk), .Q(reg_file[3416]) );
  DFFPOSX1 reg_file_reg_26__89_ ( .D(n21711), .CLK(clk), .Q(reg_file[3417]) );
  DFFPOSX1 reg_file_reg_26__90_ ( .D(n21710), .CLK(clk), .Q(reg_file[3418]) );
  DFFPOSX1 reg_file_reg_26__91_ ( .D(n21709), .CLK(clk), .Q(reg_file[3419]) );
  DFFPOSX1 reg_file_reg_26__92_ ( .D(n21708), .CLK(clk), .Q(reg_file[3420]) );
  DFFPOSX1 reg_file_reg_26__93_ ( .D(n21707), .CLK(clk), .Q(reg_file[3421]) );
  DFFPOSX1 reg_file_reg_26__94_ ( .D(n21706), .CLK(clk), .Q(reg_file[3422]) );
  DFFPOSX1 reg_file_reg_26__95_ ( .D(n21705), .CLK(clk), .Q(reg_file[3423]) );
  DFFPOSX1 reg_file_reg_26__96_ ( .D(n21704), .CLK(clk), .Q(reg_file[3424]) );
  DFFPOSX1 reg_file_reg_26__97_ ( .D(n21703), .CLK(clk), .Q(reg_file[3425]) );
  DFFPOSX1 reg_file_reg_26__98_ ( .D(n21702), .CLK(clk), .Q(reg_file[3426]) );
  DFFPOSX1 reg_file_reg_26__99_ ( .D(n21701), .CLK(clk), .Q(reg_file[3427]) );
  DFFPOSX1 reg_file_reg_26__100_ ( .D(n21700), .CLK(clk), .Q(reg_file[3428])
         );
  DFFPOSX1 reg_file_reg_26__101_ ( .D(n21699), .CLK(clk), .Q(reg_file[3429])
         );
  DFFPOSX1 reg_file_reg_26__102_ ( .D(n21698), .CLK(clk), .Q(reg_file[3430])
         );
  DFFPOSX1 reg_file_reg_26__103_ ( .D(n21697), .CLK(clk), .Q(reg_file[3431])
         );
  DFFPOSX1 reg_file_reg_26__104_ ( .D(n21696), .CLK(clk), .Q(reg_file[3432])
         );
  DFFPOSX1 reg_file_reg_26__105_ ( .D(n21695), .CLK(clk), .Q(reg_file[3433])
         );
  DFFPOSX1 reg_file_reg_26__106_ ( .D(n21694), .CLK(clk), .Q(reg_file[3434])
         );
  DFFPOSX1 reg_file_reg_26__107_ ( .D(n21693), .CLK(clk), .Q(reg_file[3435])
         );
  DFFPOSX1 reg_file_reg_26__108_ ( .D(n21692), .CLK(clk), .Q(reg_file[3436])
         );
  DFFPOSX1 reg_file_reg_26__109_ ( .D(n21691), .CLK(clk), .Q(reg_file[3437])
         );
  DFFPOSX1 reg_file_reg_26__110_ ( .D(n21690), .CLK(clk), .Q(reg_file[3438])
         );
  DFFPOSX1 reg_file_reg_26__111_ ( .D(n21689), .CLK(clk), .Q(reg_file[3439])
         );
  DFFPOSX1 reg_file_reg_26__112_ ( .D(n21688), .CLK(clk), .Q(reg_file[3440])
         );
  DFFPOSX1 reg_file_reg_26__113_ ( .D(n21687), .CLK(clk), .Q(reg_file[3441])
         );
  DFFPOSX1 reg_file_reg_26__114_ ( .D(n21686), .CLK(clk), .Q(reg_file[3442])
         );
  DFFPOSX1 reg_file_reg_26__115_ ( .D(n21685), .CLK(clk), .Q(reg_file[3443])
         );
  DFFPOSX1 reg_file_reg_26__116_ ( .D(n21684), .CLK(clk), .Q(reg_file[3444])
         );
  DFFPOSX1 reg_file_reg_26__117_ ( .D(n21683), .CLK(clk), .Q(reg_file[3445])
         );
  DFFPOSX1 reg_file_reg_26__118_ ( .D(n21682), .CLK(clk), .Q(reg_file[3446])
         );
  DFFPOSX1 reg_file_reg_26__119_ ( .D(n21681), .CLK(clk), .Q(reg_file[3447])
         );
  DFFPOSX1 reg_file_reg_26__120_ ( .D(n21680), .CLK(clk), .Q(reg_file[3448])
         );
  DFFPOSX1 reg_file_reg_26__121_ ( .D(n21679), .CLK(clk), .Q(reg_file[3449])
         );
  DFFPOSX1 reg_file_reg_26__122_ ( .D(n21678), .CLK(clk), .Q(reg_file[3450])
         );
  DFFPOSX1 reg_file_reg_26__123_ ( .D(n21677), .CLK(clk), .Q(reg_file[3451])
         );
  DFFPOSX1 reg_file_reg_26__124_ ( .D(n21676), .CLK(clk), .Q(reg_file[3452])
         );
  DFFPOSX1 reg_file_reg_26__125_ ( .D(n21675), .CLK(clk), .Q(reg_file[3453])
         );
  DFFPOSX1 reg_file_reg_26__126_ ( .D(n21674), .CLK(clk), .Q(reg_file[3454])
         );
  DFFPOSX1 reg_file_reg_26__127_ ( .D(n21673), .CLK(clk), .Q(reg_file[3455])
         );
  DFFPOSX1 reg_file_reg_27__0_ ( .D(n21672), .CLK(clk), .Q(reg_file[3456]) );
  DFFPOSX1 reg_file_reg_27__1_ ( .D(n21671), .CLK(clk), .Q(reg_file[3457]) );
  DFFPOSX1 reg_file_reg_27__2_ ( .D(n21670), .CLK(clk), .Q(reg_file[3458]) );
  DFFPOSX1 reg_file_reg_27__3_ ( .D(n21669), .CLK(clk), .Q(reg_file[3459]) );
  DFFPOSX1 reg_file_reg_27__4_ ( .D(n21668), .CLK(clk), .Q(reg_file[3460]) );
  DFFPOSX1 reg_file_reg_27__5_ ( .D(n21667), .CLK(clk), .Q(reg_file[3461]) );
  DFFPOSX1 reg_file_reg_27__6_ ( .D(n21666), .CLK(clk), .Q(reg_file[3462]) );
  DFFPOSX1 reg_file_reg_27__7_ ( .D(n21665), .CLK(clk), .Q(reg_file[3463]) );
  DFFPOSX1 reg_file_reg_27__8_ ( .D(n21664), .CLK(clk), .Q(reg_file[3464]) );
  DFFPOSX1 reg_file_reg_27__9_ ( .D(n21663), .CLK(clk), .Q(reg_file[3465]) );
  DFFPOSX1 reg_file_reg_27__10_ ( .D(n21662), .CLK(clk), .Q(reg_file[3466]) );
  DFFPOSX1 reg_file_reg_27__11_ ( .D(n21661), .CLK(clk), .Q(reg_file[3467]) );
  DFFPOSX1 reg_file_reg_27__12_ ( .D(n21660), .CLK(clk), .Q(reg_file[3468]) );
  DFFPOSX1 reg_file_reg_27__13_ ( .D(n21659), .CLK(clk), .Q(reg_file[3469]) );
  DFFPOSX1 reg_file_reg_27__14_ ( .D(n21658), .CLK(clk), .Q(reg_file[3470]) );
  DFFPOSX1 reg_file_reg_27__15_ ( .D(n21657), .CLK(clk), .Q(reg_file[3471]) );
  DFFPOSX1 reg_file_reg_27__16_ ( .D(n21656), .CLK(clk), .Q(reg_file[3472]) );
  DFFPOSX1 reg_file_reg_27__17_ ( .D(n21655), .CLK(clk), .Q(reg_file[3473]) );
  DFFPOSX1 reg_file_reg_27__18_ ( .D(n21654), .CLK(clk), .Q(reg_file[3474]) );
  DFFPOSX1 reg_file_reg_27__19_ ( .D(n21653), .CLK(clk), .Q(reg_file[3475]) );
  DFFPOSX1 reg_file_reg_27__20_ ( .D(n21652), .CLK(clk), .Q(reg_file[3476]) );
  DFFPOSX1 reg_file_reg_27__21_ ( .D(n21651), .CLK(clk), .Q(reg_file[3477]) );
  DFFPOSX1 reg_file_reg_27__22_ ( .D(n21650), .CLK(clk), .Q(reg_file[3478]) );
  DFFPOSX1 reg_file_reg_27__23_ ( .D(n21649), .CLK(clk), .Q(reg_file[3479]) );
  DFFPOSX1 reg_file_reg_27__24_ ( .D(n21648), .CLK(clk), .Q(reg_file[3480]) );
  DFFPOSX1 reg_file_reg_27__25_ ( .D(n21647), .CLK(clk), .Q(reg_file[3481]) );
  DFFPOSX1 reg_file_reg_27__26_ ( .D(n21646), .CLK(clk), .Q(reg_file[3482]) );
  DFFPOSX1 reg_file_reg_27__27_ ( .D(n21645), .CLK(clk), .Q(reg_file[3483]) );
  DFFPOSX1 reg_file_reg_27__28_ ( .D(n21644), .CLK(clk), .Q(reg_file[3484]) );
  DFFPOSX1 reg_file_reg_27__29_ ( .D(n21643), .CLK(clk), .Q(reg_file[3485]) );
  DFFPOSX1 reg_file_reg_27__30_ ( .D(n21642), .CLK(clk), .Q(reg_file[3486]) );
  DFFPOSX1 reg_file_reg_27__31_ ( .D(n21641), .CLK(clk), .Q(reg_file[3487]) );
  DFFPOSX1 reg_file_reg_27__32_ ( .D(n21640), .CLK(clk), .Q(reg_file[3488]) );
  DFFPOSX1 reg_file_reg_27__33_ ( .D(n21639), .CLK(clk), .Q(reg_file[3489]) );
  DFFPOSX1 reg_file_reg_27__34_ ( .D(n21638), .CLK(clk), .Q(reg_file[3490]) );
  DFFPOSX1 reg_file_reg_27__35_ ( .D(n21637), .CLK(clk), .Q(reg_file[3491]) );
  DFFPOSX1 reg_file_reg_27__36_ ( .D(n21636), .CLK(clk), .Q(reg_file[3492]) );
  DFFPOSX1 reg_file_reg_27__37_ ( .D(n21635), .CLK(clk), .Q(reg_file[3493]) );
  DFFPOSX1 reg_file_reg_27__38_ ( .D(n21634), .CLK(clk), .Q(reg_file[3494]) );
  DFFPOSX1 reg_file_reg_27__39_ ( .D(n21633), .CLK(clk), .Q(reg_file[3495]) );
  DFFPOSX1 reg_file_reg_27__40_ ( .D(n21632), .CLK(clk), .Q(reg_file[3496]) );
  DFFPOSX1 reg_file_reg_27__41_ ( .D(n21631), .CLK(clk), .Q(reg_file[3497]) );
  DFFPOSX1 reg_file_reg_27__42_ ( .D(n21630), .CLK(clk), .Q(reg_file[3498]) );
  DFFPOSX1 reg_file_reg_27__43_ ( .D(n21629), .CLK(clk), .Q(reg_file[3499]) );
  DFFPOSX1 reg_file_reg_27__44_ ( .D(n21628), .CLK(clk), .Q(reg_file[3500]) );
  DFFPOSX1 reg_file_reg_27__45_ ( .D(n21627), .CLK(clk), .Q(reg_file[3501]) );
  DFFPOSX1 reg_file_reg_27__46_ ( .D(n21626), .CLK(clk), .Q(reg_file[3502]) );
  DFFPOSX1 reg_file_reg_27__47_ ( .D(n21625), .CLK(clk), .Q(reg_file[3503]) );
  DFFPOSX1 reg_file_reg_27__48_ ( .D(n21624), .CLK(clk), .Q(reg_file[3504]) );
  DFFPOSX1 reg_file_reg_27__49_ ( .D(n21623), .CLK(clk), .Q(reg_file[3505]) );
  DFFPOSX1 reg_file_reg_27__50_ ( .D(n21622), .CLK(clk), .Q(reg_file[3506]) );
  DFFPOSX1 reg_file_reg_27__51_ ( .D(n21621), .CLK(clk), .Q(reg_file[3507]) );
  DFFPOSX1 reg_file_reg_27__52_ ( .D(n21620), .CLK(clk), .Q(reg_file[3508]) );
  DFFPOSX1 reg_file_reg_27__53_ ( .D(n21619), .CLK(clk), .Q(reg_file[3509]) );
  DFFPOSX1 reg_file_reg_27__54_ ( .D(n21618), .CLK(clk), .Q(reg_file[3510]) );
  DFFPOSX1 reg_file_reg_27__55_ ( .D(n21617), .CLK(clk), .Q(reg_file[3511]) );
  DFFPOSX1 reg_file_reg_27__56_ ( .D(n21616), .CLK(clk), .Q(reg_file[3512]) );
  DFFPOSX1 reg_file_reg_27__57_ ( .D(n21615), .CLK(clk), .Q(reg_file[3513]) );
  DFFPOSX1 reg_file_reg_27__58_ ( .D(n21614), .CLK(clk), .Q(reg_file[3514]) );
  DFFPOSX1 reg_file_reg_27__59_ ( .D(n21613), .CLK(clk), .Q(reg_file[3515]) );
  DFFPOSX1 reg_file_reg_27__60_ ( .D(n21612), .CLK(clk), .Q(reg_file[3516]) );
  DFFPOSX1 reg_file_reg_27__61_ ( .D(n21611), .CLK(clk), .Q(reg_file[3517]) );
  DFFPOSX1 reg_file_reg_27__62_ ( .D(n21610), .CLK(clk), .Q(reg_file[3518]) );
  DFFPOSX1 reg_file_reg_27__63_ ( .D(n21609), .CLK(clk), .Q(reg_file[3519]) );
  DFFPOSX1 reg_file_reg_27__64_ ( .D(n21608), .CLK(clk), .Q(reg_file[3520]) );
  DFFPOSX1 reg_file_reg_27__65_ ( .D(n21607), .CLK(clk), .Q(reg_file[3521]) );
  DFFPOSX1 reg_file_reg_27__66_ ( .D(n21606), .CLK(clk), .Q(reg_file[3522]) );
  DFFPOSX1 reg_file_reg_27__67_ ( .D(n21605), .CLK(clk), .Q(reg_file[3523]) );
  DFFPOSX1 reg_file_reg_27__68_ ( .D(n21604), .CLK(clk), .Q(reg_file[3524]) );
  DFFPOSX1 reg_file_reg_27__69_ ( .D(n21603), .CLK(clk), .Q(reg_file[3525]) );
  DFFPOSX1 reg_file_reg_27__70_ ( .D(n21602), .CLK(clk), .Q(reg_file[3526]) );
  DFFPOSX1 reg_file_reg_27__71_ ( .D(n21601), .CLK(clk), .Q(reg_file[3527]) );
  DFFPOSX1 reg_file_reg_27__72_ ( .D(n21600), .CLK(clk), .Q(reg_file[3528]) );
  DFFPOSX1 reg_file_reg_27__73_ ( .D(n21599), .CLK(clk), .Q(reg_file[3529]) );
  DFFPOSX1 reg_file_reg_27__74_ ( .D(n21598), .CLK(clk), .Q(reg_file[3530]) );
  DFFPOSX1 reg_file_reg_27__75_ ( .D(n21597), .CLK(clk), .Q(reg_file[3531]) );
  DFFPOSX1 reg_file_reg_27__76_ ( .D(n21596), .CLK(clk), .Q(reg_file[3532]) );
  DFFPOSX1 reg_file_reg_27__77_ ( .D(n21595), .CLK(clk), .Q(reg_file[3533]) );
  DFFPOSX1 reg_file_reg_27__78_ ( .D(n21594), .CLK(clk), .Q(reg_file[3534]) );
  DFFPOSX1 reg_file_reg_27__79_ ( .D(n21593), .CLK(clk), .Q(reg_file[3535]) );
  DFFPOSX1 reg_file_reg_27__80_ ( .D(n21592), .CLK(clk), .Q(reg_file[3536]) );
  DFFPOSX1 reg_file_reg_27__81_ ( .D(n21591), .CLK(clk), .Q(reg_file[3537]) );
  DFFPOSX1 reg_file_reg_27__82_ ( .D(n21590), .CLK(clk), .Q(reg_file[3538]) );
  DFFPOSX1 reg_file_reg_27__83_ ( .D(n21589), .CLK(clk), .Q(reg_file[3539]) );
  DFFPOSX1 reg_file_reg_27__84_ ( .D(n21588), .CLK(clk), .Q(reg_file[3540]) );
  DFFPOSX1 reg_file_reg_27__85_ ( .D(n21587), .CLK(clk), .Q(reg_file[3541]) );
  DFFPOSX1 reg_file_reg_27__86_ ( .D(n21586), .CLK(clk), .Q(reg_file[3542]) );
  DFFPOSX1 reg_file_reg_27__87_ ( .D(n21585), .CLK(clk), .Q(reg_file[3543]) );
  DFFPOSX1 reg_file_reg_27__88_ ( .D(n21584), .CLK(clk), .Q(reg_file[3544]) );
  DFFPOSX1 reg_file_reg_27__89_ ( .D(n21583), .CLK(clk), .Q(reg_file[3545]) );
  DFFPOSX1 reg_file_reg_27__90_ ( .D(n21582), .CLK(clk), .Q(reg_file[3546]) );
  DFFPOSX1 reg_file_reg_27__91_ ( .D(n21581), .CLK(clk), .Q(reg_file[3547]) );
  DFFPOSX1 reg_file_reg_27__92_ ( .D(n21580), .CLK(clk), .Q(reg_file[3548]) );
  DFFPOSX1 reg_file_reg_27__93_ ( .D(n21579), .CLK(clk), .Q(reg_file[3549]) );
  DFFPOSX1 reg_file_reg_27__94_ ( .D(n21578), .CLK(clk), .Q(reg_file[3550]) );
  DFFPOSX1 reg_file_reg_27__95_ ( .D(n21577), .CLK(clk), .Q(reg_file[3551]) );
  DFFPOSX1 reg_file_reg_27__96_ ( .D(n21576), .CLK(clk), .Q(reg_file[3552]) );
  DFFPOSX1 reg_file_reg_27__97_ ( .D(n21575), .CLK(clk), .Q(reg_file[3553]) );
  DFFPOSX1 reg_file_reg_27__98_ ( .D(n21574), .CLK(clk), .Q(reg_file[3554]) );
  DFFPOSX1 reg_file_reg_27__99_ ( .D(n21573), .CLK(clk), .Q(reg_file[3555]) );
  DFFPOSX1 reg_file_reg_27__100_ ( .D(n21572), .CLK(clk), .Q(reg_file[3556])
         );
  DFFPOSX1 reg_file_reg_27__101_ ( .D(n21571), .CLK(clk), .Q(reg_file[3557])
         );
  DFFPOSX1 reg_file_reg_27__102_ ( .D(n21570), .CLK(clk), .Q(reg_file[3558])
         );
  DFFPOSX1 reg_file_reg_27__103_ ( .D(n21569), .CLK(clk), .Q(reg_file[3559])
         );
  DFFPOSX1 reg_file_reg_27__104_ ( .D(n21568), .CLK(clk), .Q(reg_file[3560])
         );
  DFFPOSX1 reg_file_reg_27__105_ ( .D(n21567), .CLK(clk), .Q(reg_file[3561])
         );
  DFFPOSX1 reg_file_reg_27__106_ ( .D(n21566), .CLK(clk), .Q(reg_file[3562])
         );
  DFFPOSX1 reg_file_reg_27__107_ ( .D(n21565), .CLK(clk), .Q(reg_file[3563])
         );
  DFFPOSX1 reg_file_reg_27__108_ ( .D(n21564), .CLK(clk), .Q(reg_file[3564])
         );
  DFFPOSX1 reg_file_reg_27__109_ ( .D(n21563), .CLK(clk), .Q(reg_file[3565])
         );
  DFFPOSX1 reg_file_reg_27__110_ ( .D(n21562), .CLK(clk), .Q(reg_file[3566])
         );
  DFFPOSX1 reg_file_reg_27__111_ ( .D(n21561), .CLK(clk), .Q(reg_file[3567])
         );
  DFFPOSX1 reg_file_reg_27__112_ ( .D(n21560), .CLK(clk), .Q(reg_file[3568])
         );
  DFFPOSX1 reg_file_reg_27__113_ ( .D(n21559), .CLK(clk), .Q(reg_file[3569])
         );
  DFFPOSX1 reg_file_reg_27__114_ ( .D(n21558), .CLK(clk), .Q(reg_file[3570])
         );
  DFFPOSX1 reg_file_reg_27__115_ ( .D(n21557), .CLK(clk), .Q(reg_file[3571])
         );
  DFFPOSX1 reg_file_reg_27__116_ ( .D(n21556), .CLK(clk), .Q(reg_file[3572])
         );
  DFFPOSX1 reg_file_reg_27__117_ ( .D(n21555), .CLK(clk), .Q(reg_file[3573])
         );
  DFFPOSX1 reg_file_reg_27__118_ ( .D(n21554), .CLK(clk), .Q(reg_file[3574])
         );
  DFFPOSX1 reg_file_reg_27__119_ ( .D(n21553), .CLK(clk), .Q(reg_file[3575])
         );
  DFFPOSX1 reg_file_reg_27__120_ ( .D(n21552), .CLK(clk), .Q(reg_file[3576])
         );
  DFFPOSX1 reg_file_reg_27__121_ ( .D(n21551), .CLK(clk), .Q(reg_file[3577])
         );
  DFFPOSX1 reg_file_reg_27__122_ ( .D(n21550), .CLK(clk), .Q(reg_file[3578])
         );
  DFFPOSX1 reg_file_reg_27__123_ ( .D(n21549), .CLK(clk), .Q(reg_file[3579])
         );
  DFFPOSX1 reg_file_reg_27__124_ ( .D(n21548), .CLK(clk), .Q(reg_file[3580])
         );
  DFFPOSX1 reg_file_reg_27__125_ ( .D(n21547), .CLK(clk), .Q(reg_file[3581])
         );
  DFFPOSX1 reg_file_reg_27__126_ ( .D(n21546), .CLK(clk), .Q(reg_file[3582])
         );
  DFFPOSX1 reg_file_reg_27__127_ ( .D(n21545), .CLK(clk), .Q(reg_file[3583])
         );
  DFFPOSX1 reg_file_reg_28__0_ ( .D(n21544), .CLK(clk), .Q(reg_file[3584]) );
  DFFPOSX1 reg_file_reg_28__1_ ( .D(n21543), .CLK(clk), .Q(reg_file[3585]) );
  DFFPOSX1 reg_file_reg_28__2_ ( .D(n21542), .CLK(clk), .Q(reg_file[3586]) );
  DFFPOSX1 reg_file_reg_28__3_ ( .D(n21541), .CLK(clk), .Q(reg_file[3587]) );
  DFFPOSX1 reg_file_reg_28__4_ ( .D(n21540), .CLK(clk), .Q(reg_file[3588]) );
  DFFPOSX1 reg_file_reg_28__5_ ( .D(n21539), .CLK(clk), .Q(reg_file[3589]) );
  DFFPOSX1 reg_file_reg_28__6_ ( .D(n21538), .CLK(clk), .Q(reg_file[3590]) );
  DFFPOSX1 reg_file_reg_28__7_ ( .D(n21537), .CLK(clk), .Q(reg_file[3591]) );
  DFFPOSX1 reg_file_reg_28__8_ ( .D(n21536), .CLK(clk), .Q(reg_file[3592]) );
  DFFPOSX1 reg_file_reg_28__9_ ( .D(n21535), .CLK(clk), .Q(reg_file[3593]) );
  DFFPOSX1 reg_file_reg_28__10_ ( .D(n21534), .CLK(clk), .Q(reg_file[3594]) );
  DFFPOSX1 reg_file_reg_28__11_ ( .D(n21533), .CLK(clk), .Q(reg_file[3595]) );
  DFFPOSX1 reg_file_reg_28__12_ ( .D(n21532), .CLK(clk), .Q(reg_file[3596]) );
  DFFPOSX1 reg_file_reg_28__13_ ( .D(n21531), .CLK(clk), .Q(reg_file[3597]) );
  DFFPOSX1 reg_file_reg_28__14_ ( .D(n21530), .CLK(clk), .Q(reg_file[3598]) );
  DFFPOSX1 reg_file_reg_28__15_ ( .D(n21529), .CLK(clk), .Q(reg_file[3599]) );
  DFFPOSX1 reg_file_reg_28__16_ ( .D(n21528), .CLK(clk), .Q(reg_file[3600]) );
  DFFPOSX1 reg_file_reg_28__17_ ( .D(n21527), .CLK(clk), .Q(reg_file[3601]) );
  DFFPOSX1 reg_file_reg_28__18_ ( .D(n21526), .CLK(clk), .Q(reg_file[3602]) );
  DFFPOSX1 reg_file_reg_28__19_ ( .D(n21525), .CLK(clk), .Q(reg_file[3603]) );
  DFFPOSX1 reg_file_reg_28__20_ ( .D(n21524), .CLK(clk), .Q(reg_file[3604]) );
  DFFPOSX1 reg_file_reg_28__21_ ( .D(n21523), .CLK(clk), .Q(reg_file[3605]) );
  DFFPOSX1 reg_file_reg_28__22_ ( .D(n21522), .CLK(clk), .Q(reg_file[3606]) );
  DFFPOSX1 reg_file_reg_28__23_ ( .D(n21521), .CLK(clk), .Q(reg_file[3607]) );
  DFFPOSX1 reg_file_reg_28__24_ ( .D(n21520), .CLK(clk), .Q(reg_file[3608]) );
  DFFPOSX1 reg_file_reg_28__25_ ( .D(n21519), .CLK(clk), .Q(reg_file[3609]) );
  DFFPOSX1 reg_file_reg_28__26_ ( .D(n21518), .CLK(clk), .Q(reg_file[3610]) );
  DFFPOSX1 reg_file_reg_28__27_ ( .D(n21517), .CLK(clk), .Q(reg_file[3611]) );
  DFFPOSX1 reg_file_reg_28__28_ ( .D(n21516), .CLK(clk), .Q(reg_file[3612]) );
  DFFPOSX1 reg_file_reg_28__29_ ( .D(n21515), .CLK(clk), .Q(reg_file[3613]) );
  DFFPOSX1 reg_file_reg_28__30_ ( .D(n21514), .CLK(clk), .Q(reg_file[3614]) );
  DFFPOSX1 reg_file_reg_28__31_ ( .D(n21513), .CLK(clk), .Q(reg_file[3615]) );
  DFFPOSX1 reg_file_reg_28__32_ ( .D(n21512), .CLK(clk), .Q(reg_file[3616]) );
  DFFPOSX1 reg_file_reg_28__33_ ( .D(n21511), .CLK(clk), .Q(reg_file[3617]) );
  DFFPOSX1 reg_file_reg_28__34_ ( .D(n21510), .CLK(clk), .Q(reg_file[3618]) );
  DFFPOSX1 reg_file_reg_28__35_ ( .D(n21509), .CLK(clk), .Q(reg_file[3619]) );
  DFFPOSX1 reg_file_reg_28__36_ ( .D(n21508), .CLK(clk), .Q(reg_file[3620]) );
  DFFPOSX1 reg_file_reg_28__37_ ( .D(n21507), .CLK(clk), .Q(reg_file[3621]) );
  DFFPOSX1 reg_file_reg_28__38_ ( .D(n21506), .CLK(clk), .Q(reg_file[3622]) );
  DFFPOSX1 reg_file_reg_28__39_ ( .D(n21505), .CLK(clk), .Q(reg_file[3623]) );
  DFFPOSX1 reg_file_reg_28__40_ ( .D(n21504), .CLK(clk), .Q(reg_file[3624]) );
  DFFPOSX1 reg_file_reg_28__41_ ( .D(n21503), .CLK(clk), .Q(reg_file[3625]) );
  DFFPOSX1 reg_file_reg_28__42_ ( .D(n21502), .CLK(clk), .Q(reg_file[3626]) );
  DFFPOSX1 reg_file_reg_28__43_ ( .D(n21501), .CLK(clk), .Q(reg_file[3627]) );
  DFFPOSX1 reg_file_reg_28__44_ ( .D(n21500), .CLK(clk), .Q(reg_file[3628]) );
  DFFPOSX1 reg_file_reg_28__45_ ( .D(n21499), .CLK(clk), .Q(reg_file[3629]) );
  DFFPOSX1 reg_file_reg_28__46_ ( .D(n21498), .CLK(clk), .Q(reg_file[3630]) );
  DFFPOSX1 reg_file_reg_28__47_ ( .D(n21497), .CLK(clk), .Q(reg_file[3631]) );
  DFFPOSX1 reg_file_reg_28__48_ ( .D(n21496), .CLK(clk), .Q(reg_file[3632]) );
  DFFPOSX1 reg_file_reg_28__49_ ( .D(n21495), .CLK(clk), .Q(reg_file[3633]) );
  DFFPOSX1 reg_file_reg_28__50_ ( .D(n21494), .CLK(clk), .Q(reg_file[3634]) );
  DFFPOSX1 reg_file_reg_28__51_ ( .D(n21493), .CLK(clk), .Q(reg_file[3635]) );
  DFFPOSX1 reg_file_reg_28__52_ ( .D(n21492), .CLK(clk), .Q(reg_file[3636]) );
  DFFPOSX1 reg_file_reg_28__53_ ( .D(n21491), .CLK(clk), .Q(reg_file[3637]) );
  DFFPOSX1 reg_file_reg_28__54_ ( .D(n21490), .CLK(clk), .Q(reg_file[3638]) );
  DFFPOSX1 reg_file_reg_28__55_ ( .D(n21489), .CLK(clk), .Q(reg_file[3639]) );
  DFFPOSX1 reg_file_reg_28__56_ ( .D(n21488), .CLK(clk), .Q(reg_file[3640]) );
  DFFPOSX1 reg_file_reg_28__57_ ( .D(n21487), .CLK(clk), .Q(reg_file[3641]) );
  DFFPOSX1 reg_file_reg_28__58_ ( .D(n21486), .CLK(clk), .Q(reg_file[3642]) );
  DFFPOSX1 reg_file_reg_28__59_ ( .D(n21485), .CLK(clk), .Q(reg_file[3643]) );
  DFFPOSX1 reg_file_reg_28__60_ ( .D(n21484), .CLK(clk), .Q(reg_file[3644]) );
  DFFPOSX1 reg_file_reg_28__61_ ( .D(n21483), .CLK(clk), .Q(reg_file[3645]) );
  DFFPOSX1 reg_file_reg_28__62_ ( .D(n21482), .CLK(clk), .Q(reg_file[3646]) );
  DFFPOSX1 reg_file_reg_28__63_ ( .D(n21481), .CLK(clk), .Q(reg_file[3647]) );
  DFFPOSX1 reg_file_reg_28__64_ ( .D(n21480), .CLK(clk), .Q(reg_file[3648]) );
  DFFPOSX1 reg_file_reg_28__65_ ( .D(n21479), .CLK(clk), .Q(reg_file[3649]) );
  DFFPOSX1 reg_file_reg_28__66_ ( .D(n21478), .CLK(clk), .Q(reg_file[3650]) );
  DFFPOSX1 reg_file_reg_28__67_ ( .D(n21477), .CLK(clk), .Q(reg_file[3651]) );
  DFFPOSX1 reg_file_reg_28__68_ ( .D(n21476), .CLK(clk), .Q(reg_file[3652]) );
  DFFPOSX1 reg_file_reg_28__69_ ( .D(n21475), .CLK(clk), .Q(reg_file[3653]) );
  DFFPOSX1 reg_file_reg_28__70_ ( .D(n21474), .CLK(clk), .Q(reg_file[3654]) );
  DFFPOSX1 reg_file_reg_28__71_ ( .D(n21473), .CLK(clk), .Q(reg_file[3655]) );
  DFFPOSX1 reg_file_reg_28__72_ ( .D(n21472), .CLK(clk), .Q(reg_file[3656]) );
  DFFPOSX1 reg_file_reg_28__73_ ( .D(n21471), .CLK(clk), .Q(reg_file[3657]) );
  DFFPOSX1 reg_file_reg_28__74_ ( .D(n21470), .CLK(clk), .Q(reg_file[3658]) );
  DFFPOSX1 reg_file_reg_28__75_ ( .D(n21469), .CLK(clk), .Q(reg_file[3659]) );
  DFFPOSX1 reg_file_reg_28__76_ ( .D(n21468), .CLK(clk), .Q(reg_file[3660]) );
  DFFPOSX1 reg_file_reg_28__77_ ( .D(n21467), .CLK(clk), .Q(reg_file[3661]) );
  DFFPOSX1 reg_file_reg_28__78_ ( .D(n21466), .CLK(clk), .Q(reg_file[3662]) );
  DFFPOSX1 reg_file_reg_28__79_ ( .D(n21465), .CLK(clk), .Q(reg_file[3663]) );
  DFFPOSX1 reg_file_reg_28__80_ ( .D(n21464), .CLK(clk), .Q(reg_file[3664]) );
  DFFPOSX1 reg_file_reg_28__81_ ( .D(n21463), .CLK(clk), .Q(reg_file[3665]) );
  DFFPOSX1 reg_file_reg_28__82_ ( .D(n21462), .CLK(clk), .Q(reg_file[3666]) );
  DFFPOSX1 reg_file_reg_28__83_ ( .D(n21461), .CLK(clk), .Q(reg_file[3667]) );
  DFFPOSX1 reg_file_reg_28__84_ ( .D(n21460), .CLK(clk), .Q(reg_file[3668]) );
  DFFPOSX1 reg_file_reg_28__85_ ( .D(n21459), .CLK(clk), .Q(reg_file[3669]) );
  DFFPOSX1 reg_file_reg_28__86_ ( .D(n21458), .CLK(clk), .Q(reg_file[3670]) );
  DFFPOSX1 reg_file_reg_28__87_ ( .D(n21457), .CLK(clk), .Q(reg_file[3671]) );
  DFFPOSX1 reg_file_reg_28__88_ ( .D(n21456), .CLK(clk), .Q(reg_file[3672]) );
  DFFPOSX1 reg_file_reg_28__89_ ( .D(n21455), .CLK(clk), .Q(reg_file[3673]) );
  DFFPOSX1 reg_file_reg_28__90_ ( .D(n21454), .CLK(clk), .Q(reg_file[3674]) );
  DFFPOSX1 reg_file_reg_28__91_ ( .D(n21453), .CLK(clk), .Q(reg_file[3675]) );
  DFFPOSX1 reg_file_reg_28__92_ ( .D(n21452), .CLK(clk), .Q(reg_file[3676]) );
  DFFPOSX1 reg_file_reg_28__93_ ( .D(n21451), .CLK(clk), .Q(reg_file[3677]) );
  DFFPOSX1 reg_file_reg_28__94_ ( .D(n21450), .CLK(clk), .Q(reg_file[3678]) );
  DFFPOSX1 reg_file_reg_28__95_ ( .D(n21449), .CLK(clk), .Q(reg_file[3679]) );
  DFFPOSX1 reg_file_reg_28__96_ ( .D(n21448), .CLK(clk), .Q(reg_file[3680]) );
  DFFPOSX1 reg_file_reg_28__97_ ( .D(n21447), .CLK(clk), .Q(reg_file[3681]) );
  DFFPOSX1 reg_file_reg_28__98_ ( .D(n21446), .CLK(clk), .Q(reg_file[3682]) );
  DFFPOSX1 reg_file_reg_28__99_ ( .D(n21445), .CLK(clk), .Q(reg_file[3683]) );
  DFFPOSX1 reg_file_reg_28__100_ ( .D(n21444), .CLK(clk), .Q(reg_file[3684])
         );
  DFFPOSX1 reg_file_reg_28__101_ ( .D(n21443), .CLK(clk), .Q(reg_file[3685])
         );
  DFFPOSX1 reg_file_reg_28__102_ ( .D(n21442), .CLK(clk), .Q(reg_file[3686])
         );
  DFFPOSX1 reg_file_reg_28__103_ ( .D(n21441), .CLK(clk), .Q(reg_file[3687])
         );
  DFFPOSX1 reg_file_reg_28__104_ ( .D(n21440), .CLK(clk), .Q(reg_file[3688])
         );
  DFFPOSX1 reg_file_reg_28__105_ ( .D(n21439), .CLK(clk), .Q(reg_file[3689])
         );
  DFFPOSX1 reg_file_reg_28__106_ ( .D(n21438), .CLK(clk), .Q(reg_file[3690])
         );
  DFFPOSX1 reg_file_reg_28__107_ ( .D(n21437), .CLK(clk), .Q(reg_file[3691])
         );
  DFFPOSX1 reg_file_reg_28__108_ ( .D(n21436), .CLK(clk), .Q(reg_file[3692])
         );
  DFFPOSX1 reg_file_reg_28__109_ ( .D(n21435), .CLK(clk), .Q(reg_file[3693])
         );
  DFFPOSX1 reg_file_reg_28__110_ ( .D(n21434), .CLK(clk), .Q(reg_file[3694])
         );
  DFFPOSX1 reg_file_reg_28__111_ ( .D(n21433), .CLK(clk), .Q(reg_file[3695])
         );
  DFFPOSX1 reg_file_reg_28__112_ ( .D(n21432), .CLK(clk), .Q(reg_file[3696])
         );
  DFFPOSX1 reg_file_reg_28__113_ ( .D(n21431), .CLK(clk), .Q(reg_file[3697])
         );
  DFFPOSX1 reg_file_reg_28__114_ ( .D(n21430), .CLK(clk), .Q(reg_file[3698])
         );
  DFFPOSX1 reg_file_reg_28__115_ ( .D(n21429), .CLK(clk), .Q(reg_file[3699])
         );
  DFFPOSX1 reg_file_reg_28__116_ ( .D(n21428), .CLK(clk), .Q(reg_file[3700])
         );
  DFFPOSX1 reg_file_reg_28__117_ ( .D(n21427), .CLK(clk), .Q(reg_file[3701])
         );
  DFFPOSX1 reg_file_reg_28__118_ ( .D(n21426), .CLK(clk), .Q(reg_file[3702])
         );
  DFFPOSX1 reg_file_reg_28__119_ ( .D(n21425), .CLK(clk), .Q(reg_file[3703])
         );
  DFFPOSX1 reg_file_reg_28__120_ ( .D(n21424), .CLK(clk), .Q(reg_file[3704])
         );
  DFFPOSX1 reg_file_reg_28__121_ ( .D(n21423), .CLK(clk), .Q(reg_file[3705])
         );
  DFFPOSX1 reg_file_reg_28__122_ ( .D(n21422), .CLK(clk), .Q(reg_file[3706])
         );
  DFFPOSX1 reg_file_reg_28__123_ ( .D(n21421), .CLK(clk), .Q(reg_file[3707])
         );
  DFFPOSX1 reg_file_reg_28__124_ ( .D(n21420), .CLK(clk), .Q(reg_file[3708])
         );
  DFFPOSX1 reg_file_reg_28__125_ ( .D(n21419), .CLK(clk), .Q(reg_file[3709])
         );
  DFFPOSX1 reg_file_reg_28__126_ ( .D(n21418), .CLK(clk), .Q(reg_file[3710])
         );
  DFFPOSX1 reg_file_reg_28__127_ ( .D(n21417), .CLK(clk), .Q(reg_file[3711])
         );
  DFFPOSX1 reg_file_reg_29__0_ ( .D(n21416), .CLK(clk), .Q(reg_file[3712]) );
  DFFPOSX1 reg_file_reg_29__1_ ( .D(n21415), .CLK(clk), .Q(reg_file[3713]) );
  DFFPOSX1 reg_file_reg_29__2_ ( .D(n21414), .CLK(clk), .Q(reg_file[3714]) );
  DFFPOSX1 reg_file_reg_29__3_ ( .D(n21413), .CLK(clk), .Q(reg_file[3715]) );
  DFFPOSX1 reg_file_reg_29__4_ ( .D(n21412), .CLK(clk), .Q(reg_file[3716]) );
  DFFPOSX1 reg_file_reg_29__5_ ( .D(n21411), .CLK(clk), .Q(reg_file[3717]) );
  DFFPOSX1 reg_file_reg_29__6_ ( .D(n21410), .CLK(clk), .Q(reg_file[3718]) );
  DFFPOSX1 reg_file_reg_29__7_ ( .D(n21409), .CLK(clk), .Q(reg_file[3719]) );
  DFFPOSX1 reg_file_reg_29__8_ ( .D(n21408), .CLK(clk), .Q(reg_file[3720]) );
  DFFPOSX1 reg_file_reg_29__9_ ( .D(n21407), .CLK(clk), .Q(reg_file[3721]) );
  DFFPOSX1 reg_file_reg_29__10_ ( .D(n21406), .CLK(clk), .Q(reg_file[3722]) );
  DFFPOSX1 reg_file_reg_29__11_ ( .D(n21405), .CLK(clk), .Q(reg_file[3723]) );
  DFFPOSX1 reg_file_reg_29__12_ ( .D(n21404), .CLK(clk), .Q(reg_file[3724]) );
  DFFPOSX1 reg_file_reg_29__13_ ( .D(n21403), .CLK(clk), .Q(reg_file[3725]) );
  DFFPOSX1 reg_file_reg_29__14_ ( .D(n21402), .CLK(clk), .Q(reg_file[3726]) );
  DFFPOSX1 reg_file_reg_29__15_ ( .D(n21401), .CLK(clk), .Q(reg_file[3727]) );
  DFFPOSX1 reg_file_reg_29__16_ ( .D(n21400), .CLK(clk), .Q(reg_file[3728]) );
  DFFPOSX1 reg_file_reg_29__17_ ( .D(n21399), .CLK(clk), .Q(reg_file[3729]) );
  DFFPOSX1 reg_file_reg_29__18_ ( .D(n21398), .CLK(clk), .Q(reg_file[3730]) );
  DFFPOSX1 reg_file_reg_29__19_ ( .D(n21397), .CLK(clk), .Q(reg_file[3731]) );
  DFFPOSX1 reg_file_reg_29__20_ ( .D(n21396), .CLK(clk), .Q(reg_file[3732]) );
  DFFPOSX1 reg_file_reg_29__21_ ( .D(n21395), .CLK(clk), .Q(reg_file[3733]) );
  DFFPOSX1 reg_file_reg_29__22_ ( .D(n21394), .CLK(clk), .Q(reg_file[3734]) );
  DFFPOSX1 reg_file_reg_29__23_ ( .D(n21393), .CLK(clk), .Q(reg_file[3735]) );
  DFFPOSX1 reg_file_reg_29__24_ ( .D(n21392), .CLK(clk), .Q(reg_file[3736]) );
  DFFPOSX1 reg_file_reg_29__25_ ( .D(n21391), .CLK(clk), .Q(reg_file[3737]) );
  DFFPOSX1 reg_file_reg_29__26_ ( .D(n21390), .CLK(clk), .Q(reg_file[3738]) );
  DFFPOSX1 reg_file_reg_29__27_ ( .D(n21389), .CLK(clk), .Q(reg_file[3739]) );
  DFFPOSX1 reg_file_reg_29__28_ ( .D(n21388), .CLK(clk), .Q(reg_file[3740]) );
  DFFPOSX1 reg_file_reg_29__29_ ( .D(n21387), .CLK(clk), .Q(reg_file[3741]) );
  DFFPOSX1 reg_file_reg_29__30_ ( .D(n21386), .CLK(clk), .Q(reg_file[3742]) );
  DFFPOSX1 reg_file_reg_29__31_ ( .D(n21385), .CLK(clk), .Q(reg_file[3743]) );
  DFFPOSX1 reg_file_reg_29__32_ ( .D(n21384), .CLK(clk), .Q(reg_file[3744]) );
  DFFPOSX1 reg_file_reg_29__33_ ( .D(n21383), .CLK(clk), .Q(reg_file[3745]) );
  DFFPOSX1 reg_file_reg_29__34_ ( .D(n21382), .CLK(clk), .Q(reg_file[3746]) );
  DFFPOSX1 reg_file_reg_29__35_ ( .D(n21381), .CLK(clk), .Q(reg_file[3747]) );
  DFFPOSX1 reg_file_reg_29__36_ ( .D(n21380), .CLK(clk), .Q(reg_file[3748]) );
  DFFPOSX1 reg_file_reg_29__37_ ( .D(n21379), .CLK(clk), .Q(reg_file[3749]) );
  DFFPOSX1 reg_file_reg_29__38_ ( .D(n21378), .CLK(clk), .Q(reg_file[3750]) );
  DFFPOSX1 reg_file_reg_29__39_ ( .D(n21377), .CLK(clk), .Q(reg_file[3751]) );
  DFFPOSX1 reg_file_reg_29__40_ ( .D(n21376), .CLK(clk), .Q(reg_file[3752]) );
  DFFPOSX1 reg_file_reg_29__41_ ( .D(n21375), .CLK(clk), .Q(reg_file[3753]) );
  DFFPOSX1 reg_file_reg_29__42_ ( .D(n21374), .CLK(clk), .Q(reg_file[3754]) );
  DFFPOSX1 reg_file_reg_29__43_ ( .D(n21373), .CLK(clk), .Q(reg_file[3755]) );
  DFFPOSX1 reg_file_reg_29__44_ ( .D(n21372), .CLK(clk), .Q(reg_file[3756]) );
  DFFPOSX1 reg_file_reg_29__45_ ( .D(n21371), .CLK(clk), .Q(reg_file[3757]) );
  DFFPOSX1 reg_file_reg_29__46_ ( .D(n21370), .CLK(clk), .Q(reg_file[3758]) );
  DFFPOSX1 reg_file_reg_29__47_ ( .D(n21369), .CLK(clk), .Q(reg_file[3759]) );
  DFFPOSX1 reg_file_reg_29__48_ ( .D(n21368), .CLK(clk), .Q(reg_file[3760]) );
  DFFPOSX1 reg_file_reg_29__49_ ( .D(n21367), .CLK(clk), .Q(reg_file[3761]) );
  DFFPOSX1 reg_file_reg_29__50_ ( .D(n21366), .CLK(clk), .Q(reg_file[3762]) );
  DFFPOSX1 reg_file_reg_29__51_ ( .D(n21365), .CLK(clk), .Q(reg_file[3763]) );
  DFFPOSX1 reg_file_reg_29__52_ ( .D(n21364), .CLK(clk), .Q(reg_file[3764]) );
  DFFPOSX1 reg_file_reg_29__53_ ( .D(n21363), .CLK(clk), .Q(reg_file[3765]) );
  DFFPOSX1 reg_file_reg_29__54_ ( .D(n21362), .CLK(clk), .Q(reg_file[3766]) );
  DFFPOSX1 reg_file_reg_29__55_ ( .D(n21361), .CLK(clk), .Q(reg_file[3767]) );
  DFFPOSX1 reg_file_reg_29__56_ ( .D(n21360), .CLK(clk), .Q(reg_file[3768]) );
  DFFPOSX1 reg_file_reg_29__57_ ( .D(n21359), .CLK(clk), .Q(reg_file[3769]) );
  DFFPOSX1 reg_file_reg_29__58_ ( .D(n21358), .CLK(clk), .Q(reg_file[3770]) );
  DFFPOSX1 reg_file_reg_29__59_ ( .D(n21357), .CLK(clk), .Q(reg_file[3771]) );
  DFFPOSX1 reg_file_reg_29__60_ ( .D(n21356), .CLK(clk), .Q(reg_file[3772]) );
  DFFPOSX1 reg_file_reg_29__61_ ( .D(n21355), .CLK(clk), .Q(reg_file[3773]) );
  DFFPOSX1 reg_file_reg_29__62_ ( .D(n21354), .CLK(clk), .Q(reg_file[3774]) );
  DFFPOSX1 reg_file_reg_29__63_ ( .D(n21353), .CLK(clk), .Q(reg_file[3775]) );
  DFFPOSX1 reg_file_reg_29__64_ ( .D(n21352), .CLK(clk), .Q(reg_file[3776]) );
  DFFPOSX1 reg_file_reg_29__65_ ( .D(n21351), .CLK(clk), .Q(reg_file[3777]) );
  DFFPOSX1 reg_file_reg_29__66_ ( .D(n21350), .CLK(clk), .Q(reg_file[3778]) );
  DFFPOSX1 reg_file_reg_29__67_ ( .D(n21349), .CLK(clk), .Q(reg_file[3779]) );
  DFFPOSX1 reg_file_reg_29__68_ ( .D(n21348), .CLK(clk), .Q(reg_file[3780]) );
  DFFPOSX1 reg_file_reg_29__69_ ( .D(n21347), .CLK(clk), .Q(reg_file[3781]) );
  DFFPOSX1 reg_file_reg_29__70_ ( .D(n21346), .CLK(clk), .Q(reg_file[3782]) );
  DFFPOSX1 reg_file_reg_29__71_ ( .D(n21345), .CLK(clk), .Q(reg_file[3783]) );
  DFFPOSX1 reg_file_reg_29__72_ ( .D(n21344), .CLK(clk), .Q(reg_file[3784]) );
  DFFPOSX1 reg_file_reg_29__73_ ( .D(n21343), .CLK(clk), .Q(reg_file[3785]) );
  DFFPOSX1 reg_file_reg_29__74_ ( .D(n21342), .CLK(clk), .Q(reg_file[3786]) );
  DFFPOSX1 reg_file_reg_29__75_ ( .D(n21341), .CLK(clk), .Q(reg_file[3787]) );
  DFFPOSX1 reg_file_reg_29__76_ ( .D(n21340), .CLK(clk), .Q(reg_file[3788]) );
  DFFPOSX1 reg_file_reg_29__77_ ( .D(n21339), .CLK(clk), .Q(reg_file[3789]) );
  DFFPOSX1 reg_file_reg_29__78_ ( .D(n21338), .CLK(clk), .Q(reg_file[3790]) );
  DFFPOSX1 reg_file_reg_29__79_ ( .D(n21337), .CLK(clk), .Q(reg_file[3791]) );
  DFFPOSX1 reg_file_reg_29__80_ ( .D(n21336), .CLK(clk), .Q(reg_file[3792]) );
  DFFPOSX1 reg_file_reg_29__81_ ( .D(n21335), .CLK(clk), .Q(reg_file[3793]) );
  DFFPOSX1 reg_file_reg_29__82_ ( .D(n21334), .CLK(clk), .Q(reg_file[3794]) );
  DFFPOSX1 reg_file_reg_29__83_ ( .D(n21333), .CLK(clk), .Q(reg_file[3795]) );
  DFFPOSX1 reg_file_reg_29__84_ ( .D(n21332), .CLK(clk), .Q(reg_file[3796]) );
  DFFPOSX1 reg_file_reg_29__85_ ( .D(n21331), .CLK(clk), .Q(reg_file[3797]) );
  DFFPOSX1 reg_file_reg_29__86_ ( .D(n21330), .CLK(clk), .Q(reg_file[3798]) );
  DFFPOSX1 reg_file_reg_29__87_ ( .D(n21329), .CLK(clk), .Q(reg_file[3799]) );
  DFFPOSX1 reg_file_reg_29__88_ ( .D(n21328), .CLK(clk), .Q(reg_file[3800]) );
  DFFPOSX1 reg_file_reg_29__89_ ( .D(n21327), .CLK(clk), .Q(reg_file[3801]) );
  DFFPOSX1 reg_file_reg_29__90_ ( .D(n21326), .CLK(clk), .Q(reg_file[3802]) );
  DFFPOSX1 reg_file_reg_29__91_ ( .D(n21325), .CLK(clk), .Q(reg_file[3803]) );
  DFFPOSX1 reg_file_reg_29__92_ ( .D(n21324), .CLK(clk), .Q(reg_file[3804]) );
  DFFPOSX1 reg_file_reg_29__93_ ( .D(n21323), .CLK(clk), .Q(reg_file[3805]) );
  DFFPOSX1 reg_file_reg_29__94_ ( .D(n21322), .CLK(clk), .Q(reg_file[3806]) );
  DFFPOSX1 reg_file_reg_29__95_ ( .D(n21321), .CLK(clk), .Q(reg_file[3807]) );
  DFFPOSX1 reg_file_reg_29__96_ ( .D(n21320), .CLK(clk), .Q(reg_file[3808]) );
  DFFPOSX1 reg_file_reg_29__97_ ( .D(n21319), .CLK(clk), .Q(reg_file[3809]) );
  DFFPOSX1 reg_file_reg_29__98_ ( .D(n21318), .CLK(clk), .Q(reg_file[3810]) );
  DFFPOSX1 reg_file_reg_29__99_ ( .D(n21317), .CLK(clk), .Q(reg_file[3811]) );
  DFFPOSX1 reg_file_reg_29__100_ ( .D(n21316), .CLK(clk), .Q(reg_file[3812])
         );
  DFFPOSX1 reg_file_reg_29__101_ ( .D(n21315), .CLK(clk), .Q(reg_file[3813])
         );
  DFFPOSX1 reg_file_reg_29__102_ ( .D(n21314), .CLK(clk), .Q(reg_file[3814])
         );
  DFFPOSX1 reg_file_reg_29__103_ ( .D(n21313), .CLK(clk), .Q(reg_file[3815])
         );
  DFFPOSX1 reg_file_reg_29__104_ ( .D(n21312), .CLK(clk), .Q(reg_file[3816])
         );
  DFFPOSX1 reg_file_reg_29__105_ ( .D(n21311), .CLK(clk), .Q(reg_file[3817])
         );
  DFFPOSX1 reg_file_reg_29__106_ ( .D(n21310), .CLK(clk), .Q(reg_file[3818])
         );
  DFFPOSX1 reg_file_reg_29__107_ ( .D(n21309), .CLK(clk), .Q(reg_file[3819])
         );
  DFFPOSX1 reg_file_reg_29__108_ ( .D(n21308), .CLK(clk), .Q(reg_file[3820])
         );
  DFFPOSX1 reg_file_reg_29__109_ ( .D(n21307), .CLK(clk), .Q(reg_file[3821])
         );
  DFFPOSX1 reg_file_reg_29__110_ ( .D(n21306), .CLK(clk), .Q(reg_file[3822])
         );
  DFFPOSX1 reg_file_reg_29__111_ ( .D(n21305), .CLK(clk), .Q(reg_file[3823])
         );
  DFFPOSX1 reg_file_reg_29__112_ ( .D(n21304), .CLK(clk), .Q(reg_file[3824])
         );
  DFFPOSX1 reg_file_reg_29__113_ ( .D(n21303), .CLK(clk), .Q(reg_file[3825])
         );
  DFFPOSX1 reg_file_reg_29__114_ ( .D(n21302), .CLK(clk), .Q(reg_file[3826])
         );
  DFFPOSX1 reg_file_reg_29__115_ ( .D(n21301), .CLK(clk), .Q(reg_file[3827])
         );
  DFFPOSX1 reg_file_reg_29__116_ ( .D(n21300), .CLK(clk), .Q(reg_file[3828])
         );
  DFFPOSX1 reg_file_reg_29__117_ ( .D(n21299), .CLK(clk), .Q(reg_file[3829])
         );
  DFFPOSX1 reg_file_reg_29__118_ ( .D(n21298), .CLK(clk), .Q(reg_file[3830])
         );
  DFFPOSX1 reg_file_reg_29__119_ ( .D(n21297), .CLK(clk), .Q(reg_file[3831])
         );
  DFFPOSX1 reg_file_reg_29__120_ ( .D(n21296), .CLK(clk), .Q(reg_file[3832])
         );
  DFFPOSX1 reg_file_reg_29__121_ ( .D(n21295), .CLK(clk), .Q(reg_file[3833])
         );
  DFFPOSX1 reg_file_reg_29__122_ ( .D(n21294), .CLK(clk), .Q(reg_file[3834])
         );
  DFFPOSX1 reg_file_reg_29__123_ ( .D(n21293), .CLK(clk), .Q(reg_file[3835])
         );
  DFFPOSX1 reg_file_reg_29__124_ ( .D(n21292), .CLK(clk), .Q(reg_file[3836])
         );
  DFFPOSX1 reg_file_reg_29__125_ ( .D(n21291), .CLK(clk), .Q(reg_file[3837])
         );
  DFFPOSX1 reg_file_reg_29__126_ ( .D(n21290), .CLK(clk), .Q(reg_file[3838])
         );
  DFFPOSX1 reg_file_reg_29__127_ ( .D(n21289), .CLK(clk), .Q(reg_file[3839])
         );
  DFFPOSX1 reg_file_reg_30__0_ ( .D(n21288), .CLK(clk), .Q(reg_file[3840]) );
  DFFPOSX1 reg_file_reg_30__1_ ( .D(n21287), .CLK(clk), .Q(reg_file[3841]) );
  DFFPOSX1 reg_file_reg_30__2_ ( .D(n21286), .CLK(clk), .Q(reg_file[3842]) );
  DFFPOSX1 reg_file_reg_30__3_ ( .D(n21285), .CLK(clk), .Q(reg_file[3843]) );
  DFFPOSX1 reg_file_reg_30__4_ ( .D(n21284), .CLK(clk), .Q(reg_file[3844]) );
  DFFPOSX1 reg_file_reg_30__5_ ( .D(n21283), .CLK(clk), .Q(reg_file[3845]) );
  DFFPOSX1 reg_file_reg_30__6_ ( .D(n21282), .CLK(clk), .Q(reg_file[3846]) );
  DFFPOSX1 reg_file_reg_30__7_ ( .D(n21281), .CLK(clk), .Q(reg_file[3847]) );
  DFFPOSX1 reg_file_reg_30__8_ ( .D(n21280), .CLK(clk), .Q(reg_file[3848]) );
  DFFPOSX1 reg_file_reg_30__9_ ( .D(n21279), .CLK(clk), .Q(reg_file[3849]) );
  DFFPOSX1 reg_file_reg_30__10_ ( .D(n21278), .CLK(clk), .Q(reg_file[3850]) );
  DFFPOSX1 reg_file_reg_30__11_ ( .D(n21277), .CLK(clk), .Q(reg_file[3851]) );
  DFFPOSX1 reg_file_reg_30__12_ ( .D(n21276), .CLK(clk), .Q(reg_file[3852]) );
  DFFPOSX1 reg_file_reg_30__13_ ( .D(n21275), .CLK(clk), .Q(reg_file[3853]) );
  DFFPOSX1 reg_file_reg_30__14_ ( .D(n21274), .CLK(clk), .Q(reg_file[3854]) );
  DFFPOSX1 reg_file_reg_30__15_ ( .D(n21273), .CLK(clk), .Q(reg_file[3855]) );
  DFFPOSX1 reg_file_reg_30__16_ ( .D(n21272), .CLK(clk), .Q(reg_file[3856]) );
  DFFPOSX1 reg_file_reg_30__17_ ( .D(n21271), .CLK(clk), .Q(reg_file[3857]) );
  DFFPOSX1 reg_file_reg_30__18_ ( .D(n21270), .CLK(clk), .Q(reg_file[3858]) );
  DFFPOSX1 reg_file_reg_30__19_ ( .D(n21269), .CLK(clk), .Q(reg_file[3859]) );
  DFFPOSX1 reg_file_reg_30__20_ ( .D(n21268), .CLK(clk), .Q(reg_file[3860]) );
  DFFPOSX1 reg_file_reg_30__21_ ( .D(n21267), .CLK(clk), .Q(reg_file[3861]) );
  DFFPOSX1 reg_file_reg_30__22_ ( .D(n21266), .CLK(clk), .Q(reg_file[3862]) );
  DFFPOSX1 reg_file_reg_30__23_ ( .D(n21265), .CLK(clk), .Q(reg_file[3863]) );
  DFFPOSX1 reg_file_reg_30__24_ ( .D(n21264), .CLK(clk), .Q(reg_file[3864]) );
  DFFPOSX1 reg_file_reg_30__25_ ( .D(n21263), .CLK(clk), .Q(reg_file[3865]) );
  DFFPOSX1 reg_file_reg_30__26_ ( .D(n21262), .CLK(clk), .Q(reg_file[3866]) );
  DFFPOSX1 reg_file_reg_30__27_ ( .D(n21261), .CLK(clk), .Q(reg_file[3867]) );
  DFFPOSX1 reg_file_reg_30__28_ ( .D(n21260), .CLK(clk), .Q(reg_file[3868]) );
  DFFPOSX1 reg_file_reg_30__29_ ( .D(n21259), .CLK(clk), .Q(reg_file[3869]) );
  DFFPOSX1 reg_file_reg_30__30_ ( .D(n21258), .CLK(clk), .Q(reg_file[3870]) );
  DFFPOSX1 reg_file_reg_30__31_ ( .D(n21257), .CLK(clk), .Q(reg_file[3871]) );
  DFFPOSX1 reg_file_reg_30__32_ ( .D(n21256), .CLK(clk), .Q(reg_file[3872]) );
  DFFPOSX1 reg_file_reg_30__33_ ( .D(n21255), .CLK(clk), .Q(reg_file[3873]) );
  DFFPOSX1 reg_file_reg_30__34_ ( .D(n21254), .CLK(clk), .Q(reg_file[3874]) );
  DFFPOSX1 reg_file_reg_30__35_ ( .D(n21253), .CLK(clk), .Q(reg_file[3875]) );
  DFFPOSX1 reg_file_reg_30__36_ ( .D(n21252), .CLK(clk), .Q(reg_file[3876]) );
  DFFPOSX1 reg_file_reg_30__37_ ( .D(n21251), .CLK(clk), .Q(reg_file[3877]) );
  DFFPOSX1 reg_file_reg_30__38_ ( .D(n21250), .CLK(clk), .Q(reg_file[3878]) );
  DFFPOSX1 reg_file_reg_30__39_ ( .D(n21249), .CLK(clk), .Q(reg_file[3879]) );
  DFFPOSX1 reg_file_reg_30__40_ ( .D(n21248), .CLK(clk), .Q(reg_file[3880]) );
  DFFPOSX1 reg_file_reg_30__41_ ( .D(n21247), .CLK(clk), .Q(reg_file[3881]) );
  DFFPOSX1 reg_file_reg_30__42_ ( .D(n21246), .CLK(clk), .Q(reg_file[3882]) );
  DFFPOSX1 reg_file_reg_30__43_ ( .D(n21245), .CLK(clk), .Q(reg_file[3883]) );
  DFFPOSX1 reg_file_reg_30__44_ ( .D(n21244), .CLK(clk), .Q(reg_file[3884]) );
  DFFPOSX1 reg_file_reg_30__45_ ( .D(n21243), .CLK(clk), .Q(reg_file[3885]) );
  DFFPOSX1 reg_file_reg_30__46_ ( .D(n21242), .CLK(clk), .Q(reg_file[3886]) );
  DFFPOSX1 reg_file_reg_30__47_ ( .D(n21241), .CLK(clk), .Q(reg_file[3887]) );
  DFFPOSX1 reg_file_reg_30__48_ ( .D(n21240), .CLK(clk), .Q(reg_file[3888]) );
  DFFPOSX1 reg_file_reg_30__49_ ( .D(n21239), .CLK(clk), .Q(reg_file[3889]) );
  DFFPOSX1 reg_file_reg_30__50_ ( .D(n21238), .CLK(clk), .Q(reg_file[3890]) );
  DFFPOSX1 reg_file_reg_30__51_ ( .D(n21237), .CLK(clk), .Q(reg_file[3891]) );
  DFFPOSX1 reg_file_reg_30__52_ ( .D(n21236), .CLK(clk), .Q(reg_file[3892]) );
  DFFPOSX1 reg_file_reg_30__53_ ( .D(n21235), .CLK(clk), .Q(reg_file[3893]) );
  DFFPOSX1 reg_file_reg_30__54_ ( .D(n21234), .CLK(clk), .Q(reg_file[3894]) );
  DFFPOSX1 reg_file_reg_30__55_ ( .D(n21233), .CLK(clk), .Q(reg_file[3895]) );
  DFFPOSX1 reg_file_reg_30__56_ ( .D(n21232), .CLK(clk), .Q(reg_file[3896]) );
  DFFPOSX1 reg_file_reg_30__57_ ( .D(n21231), .CLK(clk), .Q(reg_file[3897]) );
  DFFPOSX1 reg_file_reg_30__58_ ( .D(n21230), .CLK(clk), .Q(reg_file[3898]) );
  DFFPOSX1 reg_file_reg_30__59_ ( .D(n21229), .CLK(clk), .Q(reg_file[3899]) );
  DFFPOSX1 reg_file_reg_30__60_ ( .D(n21228), .CLK(clk), .Q(reg_file[3900]) );
  DFFPOSX1 reg_file_reg_30__61_ ( .D(n21227), .CLK(clk), .Q(reg_file[3901]) );
  DFFPOSX1 reg_file_reg_30__62_ ( .D(n21226), .CLK(clk), .Q(reg_file[3902]) );
  DFFPOSX1 reg_file_reg_30__63_ ( .D(n21225), .CLK(clk), .Q(reg_file[3903]) );
  DFFPOSX1 reg_file_reg_30__64_ ( .D(n21224), .CLK(clk), .Q(reg_file[3904]) );
  DFFPOSX1 reg_file_reg_30__65_ ( .D(n21223), .CLK(clk), .Q(reg_file[3905]) );
  DFFPOSX1 reg_file_reg_30__66_ ( .D(n21222), .CLK(clk), .Q(reg_file[3906]) );
  DFFPOSX1 reg_file_reg_30__67_ ( .D(n21221), .CLK(clk), .Q(reg_file[3907]) );
  DFFPOSX1 reg_file_reg_30__68_ ( .D(n21220), .CLK(clk), .Q(reg_file[3908]) );
  DFFPOSX1 reg_file_reg_30__69_ ( .D(n21219), .CLK(clk), .Q(reg_file[3909]) );
  DFFPOSX1 reg_file_reg_30__70_ ( .D(n21218), .CLK(clk), .Q(reg_file[3910]) );
  DFFPOSX1 reg_file_reg_30__71_ ( .D(n21217), .CLK(clk), .Q(reg_file[3911]) );
  DFFPOSX1 reg_file_reg_30__72_ ( .D(n21216), .CLK(clk), .Q(reg_file[3912]) );
  DFFPOSX1 reg_file_reg_30__73_ ( .D(n21215), .CLK(clk), .Q(reg_file[3913]) );
  DFFPOSX1 reg_file_reg_30__74_ ( .D(n21214), .CLK(clk), .Q(reg_file[3914]) );
  DFFPOSX1 reg_file_reg_30__75_ ( .D(n21213), .CLK(clk), .Q(reg_file[3915]) );
  DFFPOSX1 reg_file_reg_30__76_ ( .D(n21212), .CLK(clk), .Q(reg_file[3916]) );
  DFFPOSX1 reg_file_reg_30__77_ ( .D(n21211), .CLK(clk), .Q(reg_file[3917]) );
  DFFPOSX1 reg_file_reg_30__78_ ( .D(n21210), .CLK(clk), .Q(reg_file[3918]) );
  DFFPOSX1 reg_file_reg_30__79_ ( .D(n21209), .CLK(clk), .Q(reg_file[3919]) );
  DFFPOSX1 reg_file_reg_30__80_ ( .D(n21208), .CLK(clk), .Q(reg_file[3920]) );
  DFFPOSX1 reg_file_reg_30__81_ ( .D(n21207), .CLK(clk), .Q(reg_file[3921]) );
  DFFPOSX1 reg_file_reg_30__82_ ( .D(n21206), .CLK(clk), .Q(reg_file[3922]) );
  DFFPOSX1 reg_file_reg_30__83_ ( .D(n21205), .CLK(clk), .Q(reg_file[3923]) );
  DFFPOSX1 reg_file_reg_30__84_ ( .D(n21204), .CLK(clk), .Q(reg_file[3924]) );
  DFFPOSX1 reg_file_reg_30__85_ ( .D(n21203), .CLK(clk), .Q(reg_file[3925]) );
  DFFPOSX1 reg_file_reg_30__86_ ( .D(n21202), .CLK(clk), .Q(reg_file[3926]) );
  DFFPOSX1 reg_file_reg_30__87_ ( .D(n21201), .CLK(clk), .Q(reg_file[3927]) );
  DFFPOSX1 reg_file_reg_30__88_ ( .D(n21200), .CLK(clk), .Q(reg_file[3928]) );
  DFFPOSX1 reg_file_reg_30__89_ ( .D(n21199), .CLK(clk), .Q(reg_file[3929]) );
  DFFPOSX1 reg_file_reg_30__90_ ( .D(n21198), .CLK(clk), .Q(reg_file[3930]) );
  DFFPOSX1 reg_file_reg_30__91_ ( .D(n21197), .CLK(clk), .Q(reg_file[3931]) );
  DFFPOSX1 reg_file_reg_30__92_ ( .D(n21196), .CLK(clk), .Q(reg_file[3932]) );
  DFFPOSX1 reg_file_reg_30__93_ ( .D(n21195), .CLK(clk), .Q(reg_file[3933]) );
  DFFPOSX1 reg_file_reg_30__94_ ( .D(n21194), .CLK(clk), .Q(reg_file[3934]) );
  DFFPOSX1 reg_file_reg_30__95_ ( .D(n21193), .CLK(clk), .Q(reg_file[3935]) );
  DFFPOSX1 reg_file_reg_30__96_ ( .D(n21192), .CLK(clk), .Q(reg_file[3936]) );
  DFFPOSX1 reg_file_reg_30__97_ ( .D(n21191), .CLK(clk), .Q(reg_file[3937]) );
  DFFPOSX1 reg_file_reg_30__98_ ( .D(n21190), .CLK(clk), .Q(reg_file[3938]) );
  DFFPOSX1 reg_file_reg_30__99_ ( .D(n21189), .CLK(clk), .Q(reg_file[3939]) );
  DFFPOSX1 reg_file_reg_30__100_ ( .D(n21188), .CLK(clk), .Q(reg_file[3940])
         );
  DFFPOSX1 reg_file_reg_30__101_ ( .D(n21187), .CLK(clk), .Q(reg_file[3941])
         );
  DFFPOSX1 reg_file_reg_30__102_ ( .D(n21186), .CLK(clk), .Q(reg_file[3942])
         );
  DFFPOSX1 reg_file_reg_30__103_ ( .D(n21185), .CLK(clk), .Q(reg_file[3943])
         );
  DFFPOSX1 reg_file_reg_30__104_ ( .D(n21184), .CLK(clk), .Q(reg_file[3944])
         );
  DFFPOSX1 reg_file_reg_30__105_ ( .D(n21183), .CLK(clk), .Q(reg_file[3945])
         );
  DFFPOSX1 reg_file_reg_30__106_ ( .D(n21182), .CLK(clk), .Q(reg_file[3946])
         );
  DFFPOSX1 reg_file_reg_30__107_ ( .D(n21181), .CLK(clk), .Q(reg_file[3947])
         );
  DFFPOSX1 reg_file_reg_30__108_ ( .D(n21180), .CLK(clk), .Q(reg_file[3948])
         );
  DFFPOSX1 reg_file_reg_30__109_ ( .D(n21179), .CLK(clk), .Q(reg_file[3949])
         );
  DFFPOSX1 reg_file_reg_30__110_ ( .D(n21178), .CLK(clk), .Q(reg_file[3950])
         );
  DFFPOSX1 reg_file_reg_30__111_ ( .D(n21177), .CLK(clk), .Q(reg_file[3951])
         );
  DFFPOSX1 reg_file_reg_30__112_ ( .D(n21176), .CLK(clk), .Q(reg_file[3952])
         );
  DFFPOSX1 reg_file_reg_30__113_ ( .D(n21175), .CLK(clk), .Q(reg_file[3953])
         );
  DFFPOSX1 reg_file_reg_30__114_ ( .D(n21174), .CLK(clk), .Q(reg_file[3954])
         );
  DFFPOSX1 reg_file_reg_30__115_ ( .D(n21173), .CLK(clk), .Q(reg_file[3955])
         );
  DFFPOSX1 reg_file_reg_30__116_ ( .D(n21172), .CLK(clk), .Q(reg_file[3956])
         );
  DFFPOSX1 reg_file_reg_30__117_ ( .D(n21171), .CLK(clk), .Q(reg_file[3957])
         );
  DFFPOSX1 reg_file_reg_30__118_ ( .D(n21170), .CLK(clk), .Q(reg_file[3958])
         );
  DFFPOSX1 reg_file_reg_30__119_ ( .D(n21169), .CLK(clk), .Q(reg_file[3959])
         );
  DFFPOSX1 reg_file_reg_30__120_ ( .D(n21168), .CLK(clk), .Q(reg_file[3960])
         );
  DFFPOSX1 reg_file_reg_30__121_ ( .D(n21167), .CLK(clk), .Q(reg_file[3961])
         );
  DFFPOSX1 reg_file_reg_30__122_ ( .D(n21166), .CLK(clk), .Q(reg_file[3962])
         );
  DFFPOSX1 reg_file_reg_30__123_ ( .D(n21165), .CLK(clk), .Q(reg_file[3963])
         );
  DFFPOSX1 reg_file_reg_30__124_ ( .D(n21164), .CLK(clk), .Q(reg_file[3964])
         );
  DFFPOSX1 reg_file_reg_30__125_ ( .D(n21163), .CLK(clk), .Q(reg_file[3965])
         );
  DFFPOSX1 reg_file_reg_30__126_ ( .D(n21162), .CLK(clk), .Q(reg_file[3966])
         );
  DFFPOSX1 reg_file_reg_30__127_ ( .D(n21161), .CLK(clk), .Q(reg_file[3967])
         );
  DFFPOSX1 reg_file_reg_31__0_ ( .D(n21160), .CLK(clk), .Q(reg_file[3968]) );
  DFFPOSX1 rd1data_reg_0_ ( .D(rd1data1033_0_), .CLK(clk), .Q(rd1data[0]) );
  DFFPOSX1 rd2data_reg_0_ ( .D(rd2data1040_0_), .CLK(clk), .Q(rd2data[0]) );
  DFFPOSX1 reg_file_reg_31__1_ ( .D(n21159), .CLK(clk), .Q(reg_file[3969]) );
  DFFPOSX1 rd1data_reg_1_ ( .D(rd1data1033_1_), .CLK(clk), .Q(rd1data[1]) );
  DFFPOSX1 rd2data_reg_1_ ( .D(rd2data1040_1_), .CLK(clk), .Q(rd2data[1]) );
  DFFPOSX1 reg_file_reg_31__2_ ( .D(n21158), .CLK(clk), .Q(reg_file[3970]) );
  DFFPOSX1 rd1data_reg_2_ ( .D(rd1data1033_2_), .CLK(clk), .Q(rd1data[2]) );
  DFFPOSX1 rd2data_reg_2_ ( .D(rd2data1040_2_), .CLK(clk), .Q(rd2data[2]) );
  DFFPOSX1 reg_file_reg_31__3_ ( .D(n21157), .CLK(clk), .Q(reg_file[3971]) );
  DFFPOSX1 rd1data_reg_3_ ( .D(rd1data1033_3_), .CLK(clk), .Q(rd1data[3]) );
  DFFPOSX1 rd2data_reg_3_ ( .D(rd2data1040_3_), .CLK(clk), .Q(rd2data[3]) );
  DFFPOSX1 reg_file_reg_31__4_ ( .D(n21156), .CLK(clk), .Q(reg_file[3972]) );
  DFFPOSX1 rd1data_reg_4_ ( .D(rd1data1033_4_), .CLK(clk), .Q(rd1data[4]) );
  DFFPOSX1 rd2data_reg_4_ ( .D(rd2data1040_4_), .CLK(clk), .Q(rd2data[4]) );
  DFFPOSX1 reg_file_reg_31__5_ ( .D(n21155), .CLK(clk), .Q(reg_file[3973]) );
  DFFPOSX1 rd1data_reg_5_ ( .D(rd1data1033_5_), .CLK(clk), .Q(rd1data[5]) );
  DFFPOSX1 rd2data_reg_5_ ( .D(rd2data1040_5_), .CLK(clk), .Q(rd2data[5]) );
  DFFPOSX1 reg_file_reg_31__6_ ( .D(n21154), .CLK(clk), .Q(reg_file[3974]) );
  DFFPOSX1 rd1data_reg_6_ ( .D(rd1data1033_6_), .CLK(clk), .Q(rd1data[6]) );
  DFFPOSX1 rd2data_reg_6_ ( .D(rd2data1040_6_), .CLK(clk), .Q(rd2data[6]) );
  DFFPOSX1 reg_file_reg_31__7_ ( .D(n21153), .CLK(clk), .Q(reg_file[3975]) );
  DFFPOSX1 rd1data_reg_7_ ( .D(rd1data1033_7_), .CLK(clk), .Q(rd1data[7]) );
  DFFPOSX1 rd2data_reg_7_ ( .D(rd2data1040_7_), .CLK(clk), .Q(rd2data[7]) );
  DFFPOSX1 reg_file_reg_31__8_ ( .D(n21152), .CLK(clk), .Q(reg_file[3976]) );
  DFFPOSX1 rd1data_reg_8_ ( .D(rd1data1033_8_), .CLK(clk), .Q(rd1data[8]) );
  DFFPOSX1 rd2data_reg_8_ ( .D(rd2data1040_8_), .CLK(clk), .Q(rd2data[8]) );
  DFFPOSX1 reg_file_reg_31__9_ ( .D(n21151), .CLK(clk), .Q(reg_file[3977]) );
  DFFPOSX1 rd1data_reg_9_ ( .D(rd1data1033_9_), .CLK(clk), .Q(rd1data[9]) );
  DFFPOSX1 rd2data_reg_9_ ( .D(rd2data1040_9_), .CLK(clk), .Q(rd2data[9]) );
  DFFPOSX1 reg_file_reg_31__10_ ( .D(n21150), .CLK(clk), .Q(reg_file[3978]) );
  DFFPOSX1 rd1data_reg_10_ ( .D(rd1data1033_10_), .CLK(clk), .Q(rd1data[10])
         );
  DFFPOSX1 rd2data_reg_10_ ( .D(rd2data1040_10_), .CLK(clk), .Q(rd2data[10])
         );
  DFFPOSX1 reg_file_reg_31__11_ ( .D(n21149), .CLK(clk), .Q(reg_file[3979]) );
  DFFPOSX1 rd1data_reg_11_ ( .D(rd1data1033_11_), .CLK(clk), .Q(rd1data[11])
         );
  DFFPOSX1 rd2data_reg_11_ ( .D(rd2data1040_11_), .CLK(clk), .Q(rd2data[11])
         );
  DFFPOSX1 reg_file_reg_31__12_ ( .D(n21148), .CLK(clk), .Q(reg_file[3980]) );
  DFFPOSX1 rd1data_reg_12_ ( .D(rd1data1033_12_), .CLK(clk), .Q(rd1data[12])
         );
  DFFPOSX1 rd2data_reg_12_ ( .D(rd2data1040_12_), .CLK(clk), .Q(rd2data[12])
         );
  DFFPOSX1 reg_file_reg_31__13_ ( .D(n21147), .CLK(clk), .Q(reg_file[3981]) );
  DFFPOSX1 rd1data_reg_13_ ( .D(rd1data1033_13_), .CLK(clk), .Q(rd1data[13])
         );
  DFFPOSX1 rd2data_reg_13_ ( .D(rd2data1040_13_), .CLK(clk), .Q(rd2data[13])
         );
  DFFPOSX1 reg_file_reg_31__14_ ( .D(n21146), .CLK(clk), .Q(reg_file[3982]) );
  DFFPOSX1 rd1data_reg_14_ ( .D(rd1data1033_14_), .CLK(clk), .Q(rd1data[14])
         );
  DFFPOSX1 rd2data_reg_14_ ( .D(rd2data1040_14_), .CLK(clk), .Q(rd2data[14])
         );
  DFFPOSX1 reg_file_reg_31__15_ ( .D(n21145), .CLK(clk), .Q(reg_file[3983]) );
  DFFPOSX1 rd1data_reg_15_ ( .D(rd1data1033_15_), .CLK(clk), .Q(rd1data[15])
         );
  DFFPOSX1 rd2data_reg_15_ ( .D(rd2data1040_15_), .CLK(clk), .Q(rd2data[15])
         );
  DFFPOSX1 reg_file_reg_31__16_ ( .D(n21144), .CLK(clk), .Q(reg_file[3984]) );
  DFFPOSX1 rd1data_reg_16_ ( .D(rd1data1033_16_), .CLK(clk), .Q(rd1data[16])
         );
  DFFPOSX1 rd2data_reg_16_ ( .D(rd2data1040_16_), .CLK(clk), .Q(rd2data[16])
         );
  DFFPOSX1 reg_file_reg_31__17_ ( .D(n21143), .CLK(clk), .Q(reg_file[3985]) );
  DFFPOSX1 rd1data_reg_17_ ( .D(rd1data1033_17_), .CLK(clk), .Q(rd1data[17])
         );
  DFFPOSX1 rd2data_reg_17_ ( .D(rd2data1040_17_), .CLK(clk), .Q(rd2data[17])
         );
  DFFPOSX1 reg_file_reg_31__18_ ( .D(n21142), .CLK(clk), .Q(reg_file[3986]) );
  DFFPOSX1 rd1data_reg_18_ ( .D(rd1data1033_18_), .CLK(clk), .Q(rd1data[18])
         );
  DFFPOSX1 rd2data_reg_18_ ( .D(rd2data1040_18_), .CLK(clk), .Q(rd2data[18])
         );
  DFFPOSX1 reg_file_reg_31__19_ ( .D(n21141), .CLK(clk), .Q(reg_file[3987]) );
  DFFPOSX1 rd1data_reg_19_ ( .D(rd1data1033_19_), .CLK(clk), .Q(rd1data[19])
         );
  DFFPOSX1 rd2data_reg_19_ ( .D(rd2data1040_19_), .CLK(clk), .Q(rd2data[19])
         );
  DFFPOSX1 reg_file_reg_31__20_ ( .D(n21140), .CLK(clk), .Q(reg_file[3988]) );
  DFFPOSX1 rd1data_reg_20_ ( .D(rd1data1033_20_), .CLK(clk), .Q(rd1data[20])
         );
  DFFPOSX1 rd2data_reg_20_ ( .D(rd2data1040_20_), .CLK(clk), .Q(rd2data[20])
         );
  DFFPOSX1 reg_file_reg_31__21_ ( .D(n21139), .CLK(clk), .Q(reg_file[3989]) );
  DFFPOSX1 rd1data_reg_21_ ( .D(rd1data1033_21_), .CLK(clk), .Q(rd1data[21])
         );
  DFFPOSX1 rd2data_reg_21_ ( .D(rd2data1040_21_), .CLK(clk), .Q(rd2data[21])
         );
  DFFPOSX1 reg_file_reg_31__22_ ( .D(n21138), .CLK(clk), .Q(reg_file[3990]) );
  DFFPOSX1 rd1data_reg_22_ ( .D(rd1data1033_22_), .CLK(clk), .Q(rd1data[22])
         );
  DFFPOSX1 rd2data_reg_22_ ( .D(rd2data1040_22_), .CLK(clk), .Q(rd2data[22])
         );
  DFFPOSX1 reg_file_reg_31__23_ ( .D(n21137), .CLK(clk), .Q(reg_file[3991]) );
  DFFPOSX1 rd1data_reg_23_ ( .D(rd1data1033_23_), .CLK(clk), .Q(rd1data[23])
         );
  DFFPOSX1 rd2data_reg_23_ ( .D(rd2data1040_23_), .CLK(clk), .Q(rd2data[23])
         );
  DFFPOSX1 reg_file_reg_31__24_ ( .D(n21136), .CLK(clk), .Q(reg_file[3992]) );
  DFFPOSX1 rd1data_reg_24_ ( .D(rd1data1033_24_), .CLK(clk), .Q(rd1data[24])
         );
  DFFPOSX1 rd2data_reg_24_ ( .D(rd2data1040_24_), .CLK(clk), .Q(rd2data[24])
         );
  DFFPOSX1 reg_file_reg_31__25_ ( .D(n21135), .CLK(clk), .Q(reg_file[3993]) );
  DFFPOSX1 rd1data_reg_25_ ( .D(rd1data1033_25_), .CLK(clk), .Q(rd1data[25])
         );
  DFFPOSX1 rd2data_reg_25_ ( .D(rd2data1040_25_), .CLK(clk), .Q(rd2data[25])
         );
  DFFPOSX1 reg_file_reg_31__26_ ( .D(n21134), .CLK(clk), .Q(reg_file[3994]) );
  DFFPOSX1 rd1data_reg_26_ ( .D(rd1data1033_26_), .CLK(clk), .Q(rd1data[26])
         );
  DFFPOSX1 rd2data_reg_26_ ( .D(rd2data1040_26_), .CLK(clk), .Q(rd2data[26])
         );
  DFFPOSX1 reg_file_reg_31__27_ ( .D(n21133), .CLK(clk), .Q(reg_file[3995]) );
  DFFPOSX1 rd1data_reg_27_ ( .D(rd1data1033_27_), .CLK(clk), .Q(rd1data[27])
         );
  DFFPOSX1 rd2data_reg_27_ ( .D(rd2data1040_27_), .CLK(clk), .Q(rd2data[27])
         );
  DFFPOSX1 reg_file_reg_31__28_ ( .D(n21132), .CLK(clk), .Q(reg_file[3996]) );
  DFFPOSX1 rd1data_reg_28_ ( .D(rd1data1033_28_), .CLK(clk), .Q(rd1data[28])
         );
  DFFPOSX1 rd2data_reg_28_ ( .D(rd2data1040_28_), .CLK(clk), .Q(rd2data[28])
         );
  DFFPOSX1 reg_file_reg_31__29_ ( .D(n21131), .CLK(clk), .Q(reg_file[3997]) );
  DFFPOSX1 rd1data_reg_29_ ( .D(rd1data1033_29_), .CLK(clk), .Q(rd1data[29])
         );
  DFFPOSX1 rd2data_reg_29_ ( .D(rd2data1040_29_), .CLK(clk), .Q(rd2data[29])
         );
  DFFPOSX1 reg_file_reg_31__30_ ( .D(n21130), .CLK(clk), .Q(reg_file[3998]) );
  DFFPOSX1 rd1data_reg_30_ ( .D(rd1data1033_30_), .CLK(clk), .Q(rd1data[30])
         );
  DFFPOSX1 rd2data_reg_30_ ( .D(rd2data1040_30_), .CLK(clk), .Q(rd2data[30])
         );
  DFFPOSX1 reg_file_reg_31__31_ ( .D(n21129), .CLK(clk), .Q(reg_file[3999]) );
  DFFPOSX1 rd1data_reg_31_ ( .D(rd1data1033_31_), .CLK(clk), .Q(rd1data[31])
         );
  DFFPOSX1 rd2data_reg_31_ ( .D(rd2data1040_31_), .CLK(clk), .Q(rd2data[31])
         );
  DFFPOSX1 reg_file_reg_31__32_ ( .D(n21128), .CLK(clk), .Q(reg_file[4000]) );
  DFFPOSX1 rd1data_reg_32_ ( .D(rd1data1033_32_), .CLK(clk), .Q(rd1data[32])
         );
  DFFPOSX1 rd2data_reg_32_ ( .D(rd2data1040_32_), .CLK(clk), .Q(rd2data[32])
         );
  DFFPOSX1 reg_file_reg_31__33_ ( .D(n21127), .CLK(clk), .Q(reg_file[4001]) );
  DFFPOSX1 rd1data_reg_33_ ( .D(rd1data1033_33_), .CLK(clk), .Q(rd1data[33])
         );
  DFFPOSX1 rd2data_reg_33_ ( .D(rd2data1040_33_), .CLK(clk), .Q(rd2data[33])
         );
  DFFPOSX1 reg_file_reg_31__34_ ( .D(n21126), .CLK(clk), .Q(reg_file[4002]) );
  DFFPOSX1 rd1data_reg_34_ ( .D(rd1data1033_34_), .CLK(clk), .Q(rd1data[34])
         );
  DFFPOSX1 rd2data_reg_34_ ( .D(rd2data1040_34_), .CLK(clk), .Q(rd2data[34])
         );
  DFFPOSX1 reg_file_reg_31__35_ ( .D(n21125), .CLK(clk), .Q(reg_file[4003]) );
  DFFPOSX1 rd1data_reg_35_ ( .D(rd1data1033_35_), .CLK(clk), .Q(rd1data[35])
         );
  DFFPOSX1 rd2data_reg_35_ ( .D(rd2data1040_35_), .CLK(clk), .Q(rd2data[35])
         );
  DFFPOSX1 reg_file_reg_31__36_ ( .D(n21124), .CLK(clk), .Q(reg_file[4004]) );
  DFFPOSX1 rd1data_reg_36_ ( .D(rd1data1033_36_), .CLK(clk), .Q(rd1data[36])
         );
  DFFPOSX1 rd2data_reg_36_ ( .D(rd2data1040_36_), .CLK(clk), .Q(rd2data[36])
         );
  DFFPOSX1 reg_file_reg_31__37_ ( .D(n21123), .CLK(clk), .Q(reg_file[4005]) );
  DFFPOSX1 rd1data_reg_37_ ( .D(rd1data1033_37_), .CLK(clk), .Q(rd1data[37])
         );
  DFFPOSX1 rd2data_reg_37_ ( .D(rd2data1040_37_), .CLK(clk), .Q(rd2data[37])
         );
  DFFPOSX1 reg_file_reg_31__38_ ( .D(n21122), .CLK(clk), .Q(reg_file[4006]) );
  DFFPOSX1 rd1data_reg_38_ ( .D(rd1data1033_38_), .CLK(clk), .Q(rd1data[38])
         );
  DFFPOSX1 rd2data_reg_38_ ( .D(rd2data1040_38_), .CLK(clk), .Q(rd2data[38])
         );
  DFFPOSX1 reg_file_reg_31__39_ ( .D(n21121), .CLK(clk), .Q(reg_file[4007]) );
  DFFPOSX1 rd1data_reg_39_ ( .D(rd1data1033_39_), .CLK(clk), .Q(rd1data[39])
         );
  DFFPOSX1 rd2data_reg_39_ ( .D(rd2data1040_39_), .CLK(clk), .Q(rd2data[39])
         );
  DFFPOSX1 reg_file_reg_31__40_ ( .D(n21120), .CLK(clk), .Q(reg_file[4008]) );
  DFFPOSX1 rd1data_reg_40_ ( .D(rd1data1033_40_), .CLK(clk), .Q(rd1data[40])
         );
  DFFPOSX1 rd2data_reg_40_ ( .D(rd2data1040_40_), .CLK(clk), .Q(rd2data[40])
         );
  DFFPOSX1 reg_file_reg_31__41_ ( .D(n21119), .CLK(clk), .Q(reg_file[4009]) );
  DFFPOSX1 rd1data_reg_41_ ( .D(rd1data1033_41_), .CLK(clk), .Q(rd1data[41])
         );
  DFFPOSX1 rd2data_reg_41_ ( .D(rd2data1040_41_), .CLK(clk), .Q(rd2data[41])
         );
  DFFPOSX1 reg_file_reg_31__42_ ( .D(n21118), .CLK(clk), .Q(reg_file[4010]) );
  DFFPOSX1 rd1data_reg_42_ ( .D(rd1data1033_42_), .CLK(clk), .Q(rd1data[42])
         );
  DFFPOSX1 rd2data_reg_42_ ( .D(rd2data1040_42_), .CLK(clk), .Q(rd2data[42])
         );
  DFFPOSX1 reg_file_reg_31__43_ ( .D(n21117), .CLK(clk), .Q(reg_file[4011]) );
  DFFPOSX1 rd1data_reg_43_ ( .D(rd1data1033_43_), .CLK(clk), .Q(rd1data[43])
         );
  DFFPOSX1 rd2data_reg_43_ ( .D(rd2data1040_43_), .CLK(clk), .Q(rd2data[43])
         );
  DFFPOSX1 reg_file_reg_31__44_ ( .D(n21116), .CLK(clk), .Q(reg_file[4012]) );
  DFFPOSX1 rd1data_reg_44_ ( .D(rd1data1033_44_), .CLK(clk), .Q(rd1data[44])
         );
  DFFPOSX1 rd2data_reg_44_ ( .D(rd2data1040_44_), .CLK(clk), .Q(rd2data[44])
         );
  DFFPOSX1 reg_file_reg_31__45_ ( .D(n21115), .CLK(clk), .Q(reg_file[4013]) );
  DFFPOSX1 rd1data_reg_45_ ( .D(rd1data1033_45_), .CLK(clk), .Q(rd1data[45])
         );
  DFFPOSX1 rd2data_reg_45_ ( .D(rd2data1040_45_), .CLK(clk), .Q(rd2data[45])
         );
  DFFPOSX1 reg_file_reg_31__46_ ( .D(n21114), .CLK(clk), .Q(reg_file[4014]) );
  DFFPOSX1 rd1data_reg_46_ ( .D(rd1data1033_46_), .CLK(clk), .Q(rd1data[46])
         );
  DFFPOSX1 rd2data_reg_46_ ( .D(rd2data1040_46_), .CLK(clk), .Q(rd2data[46])
         );
  DFFPOSX1 reg_file_reg_31__47_ ( .D(n21113), .CLK(clk), .Q(reg_file[4015]) );
  DFFPOSX1 rd1data_reg_47_ ( .D(rd1data1033_47_), .CLK(clk), .Q(rd1data[47])
         );
  DFFPOSX1 rd2data_reg_47_ ( .D(rd2data1040_47_), .CLK(clk), .Q(rd2data[47])
         );
  DFFPOSX1 reg_file_reg_31__48_ ( .D(n21112), .CLK(clk), .Q(reg_file[4016]) );
  DFFPOSX1 rd1data_reg_48_ ( .D(rd1data1033_48_), .CLK(clk), .Q(rd1data[48])
         );
  DFFPOSX1 rd2data_reg_48_ ( .D(rd2data1040_48_), .CLK(clk), .Q(rd2data[48])
         );
  DFFPOSX1 reg_file_reg_31__49_ ( .D(n21111), .CLK(clk), .Q(reg_file[4017]) );
  DFFPOSX1 rd1data_reg_49_ ( .D(rd1data1033_49_), .CLK(clk), .Q(rd1data[49])
         );
  DFFPOSX1 rd2data_reg_49_ ( .D(rd2data1040_49_), .CLK(clk), .Q(rd2data[49])
         );
  DFFPOSX1 reg_file_reg_31__50_ ( .D(n21110), .CLK(clk), .Q(reg_file[4018]) );
  DFFPOSX1 rd1data_reg_50_ ( .D(rd1data1033_50_), .CLK(clk), .Q(rd1data[50])
         );
  DFFPOSX1 rd2data_reg_50_ ( .D(rd2data1040_50_), .CLK(clk), .Q(rd2data[50])
         );
  DFFPOSX1 reg_file_reg_31__51_ ( .D(n21109), .CLK(clk), .Q(reg_file[4019]) );
  DFFPOSX1 rd1data_reg_51_ ( .D(rd1data1033_51_), .CLK(clk), .Q(rd1data[51])
         );
  DFFPOSX1 rd2data_reg_51_ ( .D(rd2data1040_51_), .CLK(clk), .Q(rd2data[51])
         );
  DFFPOSX1 reg_file_reg_31__52_ ( .D(n21108), .CLK(clk), .Q(reg_file[4020]) );
  DFFPOSX1 rd1data_reg_52_ ( .D(rd1data1033_52_), .CLK(clk), .Q(rd1data[52])
         );
  DFFPOSX1 rd2data_reg_52_ ( .D(rd2data1040_52_), .CLK(clk), .Q(rd2data[52])
         );
  DFFPOSX1 reg_file_reg_31__53_ ( .D(n21107), .CLK(clk), .Q(reg_file[4021]) );
  DFFPOSX1 rd1data_reg_53_ ( .D(rd1data1033_53_), .CLK(clk), .Q(rd1data[53])
         );
  DFFPOSX1 rd2data_reg_53_ ( .D(rd2data1040_53_), .CLK(clk), .Q(rd2data[53])
         );
  DFFPOSX1 reg_file_reg_31__54_ ( .D(n21106), .CLK(clk), .Q(reg_file[4022]) );
  DFFPOSX1 rd1data_reg_54_ ( .D(rd1data1033_54_), .CLK(clk), .Q(rd1data[54])
         );
  DFFPOSX1 rd2data_reg_54_ ( .D(rd2data1040_54_), .CLK(clk), .Q(rd2data[54])
         );
  DFFPOSX1 reg_file_reg_31__55_ ( .D(n21105), .CLK(clk), .Q(reg_file[4023]) );
  DFFPOSX1 rd1data_reg_55_ ( .D(rd1data1033_55_), .CLK(clk), .Q(rd1data[55])
         );
  DFFPOSX1 rd2data_reg_55_ ( .D(rd2data1040_55_), .CLK(clk), .Q(rd2data[55])
         );
  DFFPOSX1 reg_file_reg_31__56_ ( .D(n21104), .CLK(clk), .Q(reg_file[4024]) );
  DFFPOSX1 rd1data_reg_56_ ( .D(rd1data1033_56_), .CLK(clk), .Q(rd1data[56])
         );
  DFFPOSX1 rd2data_reg_56_ ( .D(rd2data1040_56_), .CLK(clk), .Q(rd2data[56])
         );
  DFFPOSX1 reg_file_reg_31__57_ ( .D(n21103), .CLK(clk), .Q(reg_file[4025]) );
  DFFPOSX1 rd1data_reg_57_ ( .D(rd1data1033_57_), .CLK(clk), .Q(rd1data[57])
         );
  DFFPOSX1 rd2data_reg_57_ ( .D(rd2data1040_57_), .CLK(clk), .Q(rd2data[57])
         );
  DFFPOSX1 reg_file_reg_31__58_ ( .D(n21102), .CLK(clk), .Q(reg_file[4026]) );
  DFFPOSX1 rd1data_reg_58_ ( .D(rd1data1033_58_), .CLK(clk), .Q(rd1data[58])
         );
  DFFPOSX1 rd2data_reg_58_ ( .D(rd2data1040_58_), .CLK(clk), .Q(rd2data[58])
         );
  DFFPOSX1 reg_file_reg_31__59_ ( .D(n21101), .CLK(clk), .Q(reg_file[4027]) );
  DFFPOSX1 rd1data_reg_59_ ( .D(rd1data1033_59_), .CLK(clk), .Q(rd1data[59])
         );
  DFFPOSX1 rd2data_reg_59_ ( .D(rd2data1040_59_), .CLK(clk), .Q(rd2data[59])
         );
  DFFPOSX1 reg_file_reg_31__60_ ( .D(n21100), .CLK(clk), .Q(reg_file[4028]) );
  DFFPOSX1 rd1data_reg_60_ ( .D(rd1data1033_60_), .CLK(clk), .Q(rd1data[60])
         );
  DFFPOSX1 rd2data_reg_60_ ( .D(rd2data1040_60_), .CLK(clk), .Q(rd2data[60])
         );
  DFFPOSX1 reg_file_reg_31__61_ ( .D(n21099), .CLK(clk), .Q(reg_file[4029]) );
  DFFPOSX1 rd1data_reg_61_ ( .D(rd1data1033_61_), .CLK(clk), .Q(rd1data[61])
         );
  DFFPOSX1 rd2data_reg_61_ ( .D(rd2data1040_61_), .CLK(clk), .Q(rd2data[61])
         );
  DFFPOSX1 reg_file_reg_31__62_ ( .D(n21098), .CLK(clk), .Q(reg_file[4030]) );
  DFFPOSX1 rd1data_reg_62_ ( .D(rd1data1033_62_), .CLK(clk), .Q(rd1data[62])
         );
  DFFPOSX1 rd2data_reg_62_ ( .D(rd2data1040_62_), .CLK(clk), .Q(rd2data[62])
         );
  DFFPOSX1 reg_file_reg_31__63_ ( .D(n21097), .CLK(clk), .Q(reg_file[4031]) );
  DFFPOSX1 rd1data_reg_63_ ( .D(rd1data1033_63_), .CLK(clk), .Q(rd1data[63])
         );
  DFFPOSX1 rd2data_reg_63_ ( .D(rd2data1040_63_), .CLK(clk), .Q(rd2data[63])
         );
  DFFPOSX1 reg_file_reg_31__64_ ( .D(n21096), .CLK(clk), .Q(reg_file[4032]) );
  DFFPOSX1 rd1data_reg_64_ ( .D(rd1data1033_64_), .CLK(clk), .Q(rd1data[64])
         );
  DFFPOSX1 rd2data_reg_64_ ( .D(rd2data1040_64_), .CLK(clk), .Q(rd2data[64])
         );
  DFFPOSX1 reg_file_reg_31__65_ ( .D(n21095), .CLK(clk), .Q(reg_file[4033]) );
  DFFPOSX1 rd1data_reg_65_ ( .D(rd1data1033_65_), .CLK(clk), .Q(rd1data[65])
         );
  DFFPOSX1 rd2data_reg_65_ ( .D(rd2data1040_65_), .CLK(clk), .Q(rd2data[65])
         );
  DFFPOSX1 reg_file_reg_31__66_ ( .D(n21094), .CLK(clk), .Q(reg_file[4034]) );
  DFFPOSX1 rd1data_reg_66_ ( .D(rd1data1033_66_), .CLK(clk), .Q(rd1data[66])
         );
  DFFPOSX1 rd2data_reg_66_ ( .D(rd2data1040_66_), .CLK(clk), .Q(rd2data[66])
         );
  DFFPOSX1 reg_file_reg_31__67_ ( .D(n21093), .CLK(clk), .Q(reg_file[4035]) );
  DFFPOSX1 rd1data_reg_67_ ( .D(rd1data1033_67_), .CLK(clk), .Q(rd1data[67])
         );
  DFFPOSX1 rd2data_reg_67_ ( .D(rd2data1040_67_), .CLK(clk), .Q(rd2data[67])
         );
  DFFPOSX1 reg_file_reg_31__68_ ( .D(n21092), .CLK(clk), .Q(reg_file[4036]) );
  DFFPOSX1 rd1data_reg_68_ ( .D(rd1data1033_68_), .CLK(clk), .Q(rd1data[68])
         );
  DFFPOSX1 rd2data_reg_68_ ( .D(rd2data1040_68_), .CLK(clk), .Q(rd2data[68])
         );
  DFFPOSX1 reg_file_reg_31__69_ ( .D(n21091), .CLK(clk), .Q(reg_file[4037]) );
  DFFPOSX1 rd1data_reg_69_ ( .D(rd1data1033_69_), .CLK(clk), .Q(rd1data[69])
         );
  DFFPOSX1 rd2data_reg_69_ ( .D(rd2data1040_69_), .CLK(clk), .Q(rd2data[69])
         );
  DFFPOSX1 reg_file_reg_31__70_ ( .D(n21090), .CLK(clk), .Q(reg_file[4038]) );
  DFFPOSX1 rd1data_reg_70_ ( .D(rd1data1033_70_), .CLK(clk), .Q(rd1data[70])
         );
  DFFPOSX1 rd2data_reg_70_ ( .D(rd2data1040_70_), .CLK(clk), .Q(rd2data[70])
         );
  DFFPOSX1 reg_file_reg_31__71_ ( .D(n21089), .CLK(clk), .Q(reg_file[4039]) );
  DFFPOSX1 rd1data_reg_71_ ( .D(rd1data1033_71_), .CLK(clk), .Q(rd1data[71])
         );
  DFFPOSX1 rd2data_reg_71_ ( .D(rd2data1040_71_), .CLK(clk), .Q(rd2data[71])
         );
  DFFPOSX1 reg_file_reg_31__72_ ( .D(n21088), .CLK(clk), .Q(reg_file[4040]) );
  DFFPOSX1 rd1data_reg_72_ ( .D(rd1data1033_72_), .CLK(clk), .Q(rd1data[72])
         );
  DFFPOSX1 rd2data_reg_72_ ( .D(rd2data1040_72_), .CLK(clk), .Q(rd2data[72])
         );
  DFFPOSX1 reg_file_reg_31__73_ ( .D(n21087), .CLK(clk), .Q(reg_file[4041]) );
  DFFPOSX1 rd1data_reg_73_ ( .D(rd1data1033_73_), .CLK(clk), .Q(rd1data[73])
         );
  DFFPOSX1 rd2data_reg_73_ ( .D(rd2data1040_73_), .CLK(clk), .Q(rd2data[73])
         );
  DFFPOSX1 reg_file_reg_31__74_ ( .D(n21086), .CLK(clk), .Q(reg_file[4042]) );
  DFFPOSX1 rd1data_reg_74_ ( .D(rd1data1033_74_), .CLK(clk), .Q(rd1data[74])
         );
  DFFPOSX1 rd2data_reg_74_ ( .D(rd2data1040_74_), .CLK(clk), .Q(rd2data[74])
         );
  DFFPOSX1 reg_file_reg_31__75_ ( .D(n21085), .CLK(clk), .Q(reg_file[4043]) );
  DFFPOSX1 rd1data_reg_75_ ( .D(rd1data1033_75_), .CLK(clk), .Q(rd1data[75])
         );
  DFFPOSX1 rd2data_reg_75_ ( .D(rd2data1040_75_), .CLK(clk), .Q(rd2data[75])
         );
  DFFPOSX1 reg_file_reg_31__76_ ( .D(n21084), .CLK(clk), .Q(reg_file[4044]) );
  DFFPOSX1 rd1data_reg_76_ ( .D(rd1data1033_76_), .CLK(clk), .Q(rd1data[76])
         );
  DFFPOSX1 rd2data_reg_76_ ( .D(rd2data1040_76_), .CLK(clk), .Q(rd2data[76])
         );
  DFFPOSX1 reg_file_reg_31__77_ ( .D(n21083), .CLK(clk), .Q(reg_file[4045]) );
  DFFPOSX1 rd1data_reg_77_ ( .D(rd1data1033_77_), .CLK(clk), .Q(rd1data[77])
         );
  DFFPOSX1 rd2data_reg_77_ ( .D(rd2data1040_77_), .CLK(clk), .Q(rd2data[77])
         );
  DFFPOSX1 reg_file_reg_31__78_ ( .D(n21082), .CLK(clk), .Q(reg_file[4046]) );
  DFFPOSX1 rd1data_reg_78_ ( .D(rd1data1033_78_), .CLK(clk), .Q(rd1data[78])
         );
  DFFPOSX1 rd2data_reg_78_ ( .D(rd2data1040_78_), .CLK(clk), .Q(rd2data[78])
         );
  DFFPOSX1 reg_file_reg_31__79_ ( .D(n21081), .CLK(clk), .Q(reg_file[4047]) );
  DFFPOSX1 rd1data_reg_79_ ( .D(rd1data1033_79_), .CLK(clk), .Q(rd1data[79])
         );
  DFFPOSX1 rd2data_reg_79_ ( .D(rd2data1040_79_), .CLK(clk), .Q(rd2data[79])
         );
  DFFPOSX1 reg_file_reg_31__80_ ( .D(n21080), .CLK(clk), .Q(reg_file[4048]) );
  DFFPOSX1 rd1data_reg_80_ ( .D(rd1data1033_80_), .CLK(clk), .Q(rd1data[80])
         );
  DFFPOSX1 rd2data_reg_80_ ( .D(rd2data1040_80_), .CLK(clk), .Q(rd2data[80])
         );
  DFFPOSX1 reg_file_reg_31__81_ ( .D(n21079), .CLK(clk), .Q(reg_file[4049]) );
  DFFPOSX1 rd1data_reg_81_ ( .D(rd1data1033_81_), .CLK(clk), .Q(rd1data[81])
         );
  DFFPOSX1 rd2data_reg_81_ ( .D(rd2data1040_81_), .CLK(clk), .Q(rd2data[81])
         );
  DFFPOSX1 reg_file_reg_31__82_ ( .D(n21078), .CLK(clk), .Q(reg_file[4050]) );
  DFFPOSX1 rd1data_reg_82_ ( .D(rd1data1033_82_), .CLK(clk), .Q(rd1data[82])
         );
  DFFPOSX1 rd2data_reg_82_ ( .D(rd2data1040_82_), .CLK(clk), .Q(rd2data[82])
         );
  DFFPOSX1 reg_file_reg_31__83_ ( .D(n21077), .CLK(clk), .Q(reg_file[4051]) );
  DFFPOSX1 rd1data_reg_83_ ( .D(rd1data1033_83_), .CLK(clk), .Q(rd1data[83])
         );
  DFFPOSX1 rd2data_reg_83_ ( .D(rd2data1040_83_), .CLK(clk), .Q(rd2data[83])
         );
  DFFPOSX1 reg_file_reg_31__84_ ( .D(n21076), .CLK(clk), .Q(reg_file[4052]) );
  DFFPOSX1 rd1data_reg_84_ ( .D(rd1data1033_84_), .CLK(clk), .Q(rd1data[84])
         );
  DFFPOSX1 rd2data_reg_84_ ( .D(rd2data1040_84_), .CLK(clk), .Q(rd2data[84])
         );
  DFFPOSX1 reg_file_reg_31__85_ ( .D(n21075), .CLK(clk), .Q(reg_file[4053]) );
  DFFPOSX1 rd1data_reg_85_ ( .D(rd1data1033_85_), .CLK(clk), .Q(rd1data[85])
         );
  DFFPOSX1 rd2data_reg_85_ ( .D(rd2data1040_85_), .CLK(clk), .Q(rd2data[85])
         );
  DFFPOSX1 reg_file_reg_31__86_ ( .D(n21074), .CLK(clk), .Q(reg_file[4054]) );
  DFFPOSX1 rd1data_reg_86_ ( .D(rd1data1033_86_), .CLK(clk), .Q(rd1data[86])
         );
  DFFPOSX1 rd2data_reg_86_ ( .D(rd2data1040_86_), .CLK(clk), .Q(rd2data[86])
         );
  DFFPOSX1 reg_file_reg_31__87_ ( .D(n21073), .CLK(clk), .Q(reg_file[4055]) );
  DFFPOSX1 rd1data_reg_87_ ( .D(rd1data1033_87_), .CLK(clk), .Q(rd1data[87])
         );
  DFFPOSX1 rd2data_reg_87_ ( .D(rd2data1040_87_), .CLK(clk), .Q(rd2data[87])
         );
  DFFPOSX1 reg_file_reg_31__88_ ( .D(n21072), .CLK(clk), .Q(reg_file[4056]) );
  DFFPOSX1 rd1data_reg_88_ ( .D(rd1data1033_88_), .CLK(clk), .Q(rd1data[88])
         );
  DFFPOSX1 rd2data_reg_88_ ( .D(rd2data1040_88_), .CLK(clk), .Q(rd2data[88])
         );
  DFFPOSX1 reg_file_reg_31__89_ ( .D(n21071), .CLK(clk), .Q(reg_file[4057]) );
  DFFPOSX1 rd1data_reg_89_ ( .D(rd1data1033_89_), .CLK(clk), .Q(rd1data[89])
         );
  DFFPOSX1 rd2data_reg_89_ ( .D(rd2data1040_89_), .CLK(clk), .Q(rd2data[89])
         );
  DFFPOSX1 reg_file_reg_31__90_ ( .D(n21070), .CLK(clk), .Q(reg_file[4058]) );
  DFFPOSX1 rd1data_reg_90_ ( .D(rd1data1033_90_), .CLK(clk), .Q(rd1data[90])
         );
  DFFPOSX1 rd2data_reg_90_ ( .D(rd2data1040_90_), .CLK(clk), .Q(rd2data[90])
         );
  DFFPOSX1 reg_file_reg_31__91_ ( .D(n21069), .CLK(clk), .Q(reg_file[4059]) );
  DFFPOSX1 rd1data_reg_91_ ( .D(rd1data1033_91_), .CLK(clk), .Q(rd1data[91])
         );
  DFFPOSX1 rd2data_reg_91_ ( .D(rd2data1040_91_), .CLK(clk), .Q(rd2data[91])
         );
  DFFPOSX1 reg_file_reg_31__92_ ( .D(n21068), .CLK(clk), .Q(reg_file[4060]) );
  DFFPOSX1 rd1data_reg_92_ ( .D(rd1data1033_92_), .CLK(clk), .Q(rd1data[92])
         );
  DFFPOSX1 rd2data_reg_92_ ( .D(rd2data1040_92_), .CLK(clk), .Q(rd2data[92])
         );
  DFFPOSX1 reg_file_reg_31__93_ ( .D(n21067), .CLK(clk), .Q(reg_file[4061]) );
  DFFPOSX1 rd1data_reg_93_ ( .D(rd1data1033_93_), .CLK(clk), .Q(rd1data[93])
         );
  DFFPOSX1 rd2data_reg_93_ ( .D(rd2data1040_93_), .CLK(clk), .Q(rd2data[93])
         );
  DFFPOSX1 reg_file_reg_31__94_ ( .D(n21066), .CLK(clk), .Q(reg_file[4062]) );
  DFFPOSX1 rd1data_reg_94_ ( .D(rd1data1033_94_), .CLK(clk), .Q(rd1data[94])
         );
  DFFPOSX1 rd2data_reg_94_ ( .D(rd2data1040_94_), .CLK(clk), .Q(rd2data[94])
         );
  DFFPOSX1 reg_file_reg_31__95_ ( .D(n21065), .CLK(clk), .Q(reg_file[4063]) );
  DFFPOSX1 rd1data_reg_95_ ( .D(rd1data1033_95_), .CLK(clk), .Q(rd1data[95])
         );
  DFFPOSX1 rd2data_reg_95_ ( .D(rd2data1040_95_), .CLK(clk), .Q(rd2data[95])
         );
  DFFPOSX1 reg_file_reg_31__96_ ( .D(n21064), .CLK(clk), .Q(reg_file[4064]) );
  DFFPOSX1 rd1data_reg_96_ ( .D(rd1data1033_96_), .CLK(clk), .Q(rd1data[96])
         );
  DFFPOSX1 rd2data_reg_96_ ( .D(rd2data1040_96_), .CLK(clk), .Q(rd2data[96])
         );
  DFFPOSX1 reg_file_reg_31__97_ ( .D(n21063), .CLK(clk), .Q(reg_file[4065]) );
  DFFPOSX1 rd1data_reg_97_ ( .D(rd1data1033_97_), .CLK(clk), .Q(rd1data[97])
         );
  DFFPOSX1 rd2data_reg_97_ ( .D(rd2data1040_97_), .CLK(clk), .Q(rd2data[97])
         );
  DFFPOSX1 reg_file_reg_31__98_ ( .D(n21062), .CLK(clk), .Q(reg_file[4066]) );
  DFFPOSX1 rd1data_reg_98_ ( .D(rd1data1033_98_), .CLK(clk), .Q(rd1data[98])
         );
  DFFPOSX1 rd2data_reg_98_ ( .D(rd2data1040_98_), .CLK(clk), .Q(rd2data[98])
         );
  DFFPOSX1 reg_file_reg_31__99_ ( .D(n21061), .CLK(clk), .Q(reg_file[4067]) );
  DFFPOSX1 rd1data_reg_99_ ( .D(rd1data1033_99_), .CLK(clk), .Q(rd1data[99])
         );
  DFFPOSX1 rd2data_reg_99_ ( .D(rd2data1040_99_), .CLK(clk), .Q(rd2data[99])
         );
  DFFPOSX1 reg_file_reg_31__100_ ( .D(n21060), .CLK(clk), .Q(reg_file[4068])
         );
  DFFPOSX1 rd1data_reg_100_ ( .D(rd1data1033_100_), .CLK(clk), .Q(rd1data[100]) );
  DFFPOSX1 rd2data_reg_100_ ( .D(rd2data1040_100_), .CLK(clk), .Q(rd2data[100]) );
  DFFPOSX1 reg_file_reg_31__101_ ( .D(n21059), .CLK(clk), .Q(reg_file[4069])
         );
  DFFPOSX1 rd1data_reg_101_ ( .D(rd1data1033_101_), .CLK(clk), .Q(rd1data[101]) );
  DFFPOSX1 rd2data_reg_101_ ( .D(rd2data1040_101_), .CLK(clk), .Q(rd2data[101]) );
  DFFPOSX1 reg_file_reg_31__102_ ( .D(n21058), .CLK(clk), .Q(reg_file[4070])
         );
  DFFPOSX1 rd1data_reg_102_ ( .D(rd1data1033_102_), .CLK(clk), .Q(rd1data[102]) );
  DFFPOSX1 rd2data_reg_102_ ( .D(rd2data1040_102_), .CLK(clk), .Q(rd2data[102]) );
  DFFPOSX1 reg_file_reg_31__103_ ( .D(n21057), .CLK(clk), .Q(reg_file[4071])
         );
  DFFPOSX1 rd1data_reg_103_ ( .D(rd1data1033_103_), .CLK(clk), .Q(rd1data[103]) );
  DFFPOSX1 rd2data_reg_103_ ( .D(rd2data1040_103_), .CLK(clk), .Q(rd2data[103]) );
  DFFPOSX1 reg_file_reg_31__104_ ( .D(n21056), .CLK(clk), .Q(reg_file[4072])
         );
  DFFPOSX1 rd1data_reg_104_ ( .D(rd1data1033_104_), .CLK(clk), .Q(rd1data[104]) );
  DFFPOSX1 rd2data_reg_104_ ( .D(rd2data1040_104_), .CLK(clk), .Q(rd2data[104]) );
  DFFPOSX1 reg_file_reg_31__105_ ( .D(n21055), .CLK(clk), .Q(reg_file[4073])
         );
  DFFPOSX1 rd1data_reg_105_ ( .D(rd1data1033_105_), .CLK(clk), .Q(rd1data[105]) );
  DFFPOSX1 rd2data_reg_105_ ( .D(rd2data1040_105_), .CLK(clk), .Q(rd2data[105]) );
  DFFPOSX1 reg_file_reg_31__106_ ( .D(n21054), .CLK(clk), .Q(reg_file[4074])
         );
  DFFPOSX1 rd1data_reg_106_ ( .D(rd1data1033_106_), .CLK(clk), .Q(rd1data[106]) );
  DFFPOSX1 rd2data_reg_106_ ( .D(rd2data1040_106_), .CLK(clk), .Q(rd2data[106]) );
  DFFPOSX1 reg_file_reg_31__107_ ( .D(n21053), .CLK(clk), .Q(reg_file[4075])
         );
  DFFPOSX1 rd1data_reg_107_ ( .D(rd1data1033_107_), .CLK(clk), .Q(rd1data[107]) );
  DFFPOSX1 rd2data_reg_107_ ( .D(rd2data1040_107_), .CLK(clk), .Q(rd2data[107]) );
  DFFPOSX1 reg_file_reg_31__108_ ( .D(n21052), .CLK(clk), .Q(reg_file[4076])
         );
  DFFPOSX1 rd1data_reg_108_ ( .D(rd1data1033_108_), .CLK(clk), .Q(rd1data[108]) );
  DFFPOSX1 rd2data_reg_108_ ( .D(rd2data1040_108_), .CLK(clk), .Q(rd2data[108]) );
  DFFPOSX1 reg_file_reg_31__109_ ( .D(n21051), .CLK(clk), .Q(reg_file[4077])
         );
  DFFPOSX1 rd1data_reg_109_ ( .D(rd1data1033_109_), .CLK(clk), .Q(rd1data[109]) );
  DFFPOSX1 rd2data_reg_109_ ( .D(rd2data1040_109_), .CLK(clk), .Q(rd2data[109]) );
  DFFPOSX1 reg_file_reg_31__110_ ( .D(n21050), .CLK(clk), .Q(reg_file[4078])
         );
  DFFPOSX1 rd1data_reg_110_ ( .D(rd1data1033_110_), .CLK(clk), .Q(rd1data[110]) );
  DFFPOSX1 rd2data_reg_110_ ( .D(rd2data1040_110_), .CLK(clk), .Q(rd2data[110]) );
  DFFPOSX1 reg_file_reg_31__111_ ( .D(n21049), .CLK(clk), .Q(reg_file[4079])
         );
  DFFPOSX1 rd1data_reg_111_ ( .D(rd1data1033_111_), .CLK(clk), .Q(rd1data[111]) );
  DFFPOSX1 rd2data_reg_111_ ( .D(rd2data1040_111_), .CLK(clk), .Q(rd2data[111]) );
  DFFPOSX1 reg_file_reg_31__112_ ( .D(n21048), .CLK(clk), .Q(reg_file[4080])
         );
  DFFPOSX1 rd1data_reg_112_ ( .D(rd1data1033_112_), .CLK(clk), .Q(rd1data[112]) );
  DFFPOSX1 rd2data_reg_112_ ( .D(rd2data1040_112_), .CLK(clk), .Q(rd2data[112]) );
  DFFPOSX1 reg_file_reg_31__113_ ( .D(n21047), .CLK(clk), .Q(reg_file[4081])
         );
  DFFPOSX1 rd1data_reg_113_ ( .D(rd1data1033_113_), .CLK(clk), .Q(rd1data[113]) );
  DFFPOSX1 rd2data_reg_113_ ( .D(rd2data1040_113_), .CLK(clk), .Q(rd2data[113]) );
  DFFPOSX1 reg_file_reg_31__114_ ( .D(n21046), .CLK(clk), .Q(reg_file[4082])
         );
  DFFPOSX1 rd1data_reg_114_ ( .D(rd1data1033_114_), .CLK(clk), .Q(rd1data[114]) );
  DFFPOSX1 rd2data_reg_114_ ( .D(rd2data1040_114_), .CLK(clk), .Q(rd2data[114]) );
  DFFPOSX1 reg_file_reg_31__115_ ( .D(n21045), .CLK(clk), .Q(reg_file[4083])
         );
  DFFPOSX1 rd1data_reg_115_ ( .D(rd1data1033_115_), .CLK(clk), .Q(rd1data[115]) );
  DFFPOSX1 rd2data_reg_115_ ( .D(rd2data1040_115_), .CLK(clk), .Q(rd2data[115]) );
  DFFPOSX1 reg_file_reg_31__116_ ( .D(n21044), .CLK(clk), .Q(reg_file[4084])
         );
  DFFPOSX1 rd1data_reg_116_ ( .D(rd1data1033_116_), .CLK(clk), .Q(rd1data[116]) );
  DFFPOSX1 rd2data_reg_116_ ( .D(rd2data1040_116_), .CLK(clk), .Q(rd2data[116]) );
  DFFPOSX1 reg_file_reg_31__117_ ( .D(n21043), .CLK(clk), .Q(reg_file[4085])
         );
  DFFPOSX1 rd1data_reg_117_ ( .D(rd1data1033_117_), .CLK(clk), .Q(rd1data[117]) );
  DFFPOSX1 rd2data_reg_117_ ( .D(rd2data1040_117_), .CLK(clk), .Q(rd2data[117]) );
  DFFPOSX1 reg_file_reg_31__118_ ( .D(n21042), .CLK(clk), .Q(reg_file[4086])
         );
  DFFPOSX1 rd1data_reg_118_ ( .D(rd1data1033_118_), .CLK(clk), .Q(rd1data[118]) );
  DFFPOSX1 rd2data_reg_118_ ( .D(rd2data1040_118_), .CLK(clk), .Q(rd2data[118]) );
  DFFPOSX1 reg_file_reg_31__119_ ( .D(n21041), .CLK(clk), .Q(reg_file[4087])
         );
  DFFPOSX1 rd1data_reg_119_ ( .D(rd1data1033_119_), .CLK(clk), .Q(rd1data[119]) );
  DFFPOSX1 rd2data_reg_119_ ( .D(rd2data1040_119_), .CLK(clk), .Q(rd2data[119]) );
  DFFPOSX1 reg_file_reg_31__120_ ( .D(n21040), .CLK(clk), .Q(reg_file[4088])
         );
  DFFPOSX1 rd1data_reg_120_ ( .D(rd1data1033_120_), .CLK(clk), .Q(rd1data[120]) );
  DFFPOSX1 rd2data_reg_120_ ( .D(rd2data1040_120_), .CLK(clk), .Q(rd2data[120]) );
  DFFPOSX1 reg_file_reg_31__121_ ( .D(n21039), .CLK(clk), .Q(reg_file[4089])
         );
  DFFPOSX1 rd1data_reg_121_ ( .D(rd1data1033_121_), .CLK(clk), .Q(rd1data[121]) );
  DFFPOSX1 rd2data_reg_121_ ( .D(rd2data1040_121_), .CLK(clk), .Q(rd2data[121]) );
  DFFPOSX1 reg_file_reg_31__122_ ( .D(n21038), .CLK(clk), .Q(reg_file[4090])
         );
  DFFPOSX1 rd1data_reg_122_ ( .D(rd1data1033_122_), .CLK(clk), .Q(rd1data[122]) );
  DFFPOSX1 rd2data_reg_122_ ( .D(rd2data1040_122_), .CLK(clk), .Q(rd2data[122]) );
  DFFPOSX1 reg_file_reg_31__123_ ( .D(n21037), .CLK(clk), .Q(reg_file[4091])
         );
  DFFPOSX1 rd1data_reg_123_ ( .D(rd1data1033_123_), .CLK(clk), .Q(rd1data[123]) );
  DFFPOSX1 rd2data_reg_123_ ( .D(rd2data1040_123_), .CLK(clk), .Q(rd2data[123]) );
  DFFPOSX1 reg_file_reg_31__124_ ( .D(n21036), .CLK(clk), .Q(reg_file[4092])
         );
  DFFPOSX1 rd1data_reg_124_ ( .D(rd1data1033_124_), .CLK(clk), .Q(rd1data[124]) );
  DFFPOSX1 rd2data_reg_124_ ( .D(rd2data1040_124_), .CLK(clk), .Q(rd2data[124]) );
  DFFPOSX1 reg_file_reg_31__125_ ( .D(n21035), .CLK(clk), .Q(reg_file[4093])
         );
  DFFPOSX1 rd1data_reg_125_ ( .D(rd1data1033_125_), .CLK(clk), .Q(rd1data[125]) );
  DFFPOSX1 rd2data_reg_125_ ( .D(rd2data1040_125_), .CLK(clk), .Q(rd2data[125]) );
  DFFPOSX1 reg_file_reg_31__126_ ( .D(n21034), .CLK(clk), .Q(reg_file[4094])
         );
  DFFPOSX1 rd1data_reg_126_ ( .D(rd1data1033_126_), .CLK(clk), .Q(rd1data[126]) );
  DFFPOSX1 rd2data_reg_126_ ( .D(rd2data1040_126_), .CLK(clk), .Q(rd2data[126]) );
  DFFPOSX1 reg_file_reg_31__127_ ( .D(n21033), .CLK(clk), .Q(reg_file[4095])
         );
  DFFPOSX1 rd1data_reg_127_ ( .D(rd1data1033_127_), .CLK(clk), .Q(rd1data[127]) );
  DFFPOSX1 rd2data_reg_127_ ( .D(rd2data1040_127_), .CLK(clk), .Q(rd2data[127]) );
  BUFX2 U14324 ( .A(n34913), .Y(n25129) );
  BUFX2 U14325 ( .A(n34915), .Y(n25130) );
  BUFX2 U14326 ( .A(n34916), .Y(n25131) );
  BUFX2 U14327 ( .A(n34917), .Y(n25132) );
  BUFX2 U14328 ( .A(n34918), .Y(n25133) );
  BUFX2 U14329 ( .A(n34919), .Y(n25134) );
  BUFX2 U14330 ( .A(n34920), .Y(n25135) );
  BUFX2 U14331 ( .A(n34921), .Y(n25136) );
  BUFX2 U14332 ( .A(n34914), .Y(n25839) );
  BUFX2 U14333 ( .A(n34914), .Y(n25845) );
  BUFX2 U14334 ( .A(n34914), .Y(n25844) );
  BUFX2 U14335 ( .A(n34914), .Y(n25843) );
  BUFX2 U14336 ( .A(n34914), .Y(n25842) );
  BUFX2 U14337 ( .A(n34914), .Y(n25841) );
  BUFX2 U14338 ( .A(n34914), .Y(n25840) );
  BUFX2 U14339 ( .A(n34914), .Y(n25846) );
  BUFX2 U14340 ( .A(n36625), .Y(n26039) );
  BUFX2 U14341 ( .A(n36495), .Y(n26031) );
  BUFX2 U14342 ( .A(n36103), .Y(n25975) );
  BUFX2 U14343 ( .A(n35973), .Y(n25967) );
  BUFX2 U14344 ( .A(n35581), .Y(n25911) );
  BUFX2 U14345 ( .A(n35451), .Y(n25903) );
  BUFX2 U14346 ( .A(n34924), .Y(n25847) );
  BUFX2 U14347 ( .A(n37018), .Y(n26087) );
  BUFX2 U14348 ( .A(n37017), .Y(n26079) );
  BUFX2 U14349 ( .A(n36493), .Y(n26023) );
  BUFX2 U14350 ( .A(n36492), .Y(n26015) );
  BUFX2 U14351 ( .A(n35971), .Y(n25959) );
  BUFX2 U14352 ( .A(n35970), .Y(n25951) );
  BUFX2 U14353 ( .A(n37016), .Y(n26071) );
  BUFX2 U14354 ( .A(n37015), .Y(n26063) );
  BUFX2 U14355 ( .A(n36887), .Y(n26055) );
  BUFX2 U14356 ( .A(n36758), .Y(n26047) );
  BUFX2 U14357 ( .A(n36491), .Y(n26007) );
  BUFX2 U14358 ( .A(n36490), .Y(n25999) );
  BUFX2 U14359 ( .A(n36362), .Y(n25991) );
  BUFX2 U14360 ( .A(n36233), .Y(n25983) );
  BUFX2 U14361 ( .A(n35969), .Y(n25943) );
  BUFX2 U14362 ( .A(n35968), .Y(n25935) );
  BUFX2 U14363 ( .A(n35840), .Y(n25927) );
  BUFX2 U14364 ( .A(n35711), .Y(n25919) );
  BUFX2 U14365 ( .A(n35322), .Y(n25895) );
  BUFX2 U14366 ( .A(n35189), .Y(n25887) );
  BUFX2 U14367 ( .A(n35060), .Y(n25879) );
  BUFX2 U14368 ( .A(n34930), .Y(n25871) );
  BUFX2 U14369 ( .A(n34928), .Y(n25863) );
  BUFX2 U14370 ( .A(n34926), .Y(n25855) );
  BUFX2 U14371 ( .A(n31552), .Y(n25594) );
  BUFX2 U14372 ( .A(n31554), .Y(n25615) );
  BUFX2 U14373 ( .A(n31552), .Y(n25593) );
  BUFX2 U14374 ( .A(n31554), .Y(n25614) );
  BUFX2 U14375 ( .A(n31552), .Y(n25600) );
  BUFX2 U14376 ( .A(n31554), .Y(n25621) );
  BUFX2 U14377 ( .A(n31552), .Y(n25599) );
  BUFX2 U14378 ( .A(n31554), .Y(n25620) );
  BUFX2 U14379 ( .A(n31552), .Y(n25598) );
  BUFX2 U14380 ( .A(n31554), .Y(n25619) );
  BUFX2 U14381 ( .A(n31552), .Y(n25597) );
  BUFX2 U14382 ( .A(n31554), .Y(n25618) );
  BUFX2 U14383 ( .A(n31552), .Y(n25596) );
  BUFX2 U14384 ( .A(n31554), .Y(n25617) );
  BUFX2 U14385 ( .A(n31552), .Y(n25595) );
  BUFX2 U14386 ( .A(n31554), .Y(n25616) );
  BUFX2 U14387 ( .A(n31552), .Y(n25592) );
  BUFX2 U14388 ( .A(n31554), .Y(n25613) );
  BUFX2 U14389 ( .A(n36625), .Y(n26045) );
  BUFX2 U14390 ( .A(n36625), .Y(n26044) );
  BUFX2 U14391 ( .A(n36625), .Y(n26043) );
  BUFX2 U14392 ( .A(n36625), .Y(n26042) );
  BUFX2 U14393 ( .A(n36625), .Y(n26041) );
  BUFX2 U14394 ( .A(n36625), .Y(n26040) );
  BUFX2 U14395 ( .A(n36495), .Y(n26037) );
  BUFX2 U14396 ( .A(n36495), .Y(n26036) );
  BUFX2 U14397 ( .A(n36495), .Y(n26035) );
  BUFX2 U14398 ( .A(n36495), .Y(n26034) );
  BUFX2 U14399 ( .A(n36495), .Y(n26033) );
  BUFX2 U14400 ( .A(n36495), .Y(n26032) );
  BUFX2 U14401 ( .A(n36103), .Y(n25981) );
  BUFX2 U14402 ( .A(n36103), .Y(n25980) );
  BUFX2 U14403 ( .A(n36103), .Y(n25979) );
  BUFX2 U14404 ( .A(n36103), .Y(n25978) );
  BUFX2 U14405 ( .A(n36103), .Y(n25977) );
  BUFX2 U14406 ( .A(n36103), .Y(n25976) );
  BUFX2 U14407 ( .A(n35973), .Y(n25973) );
  BUFX2 U14408 ( .A(n35973), .Y(n25972) );
  BUFX2 U14409 ( .A(n35973), .Y(n25971) );
  BUFX2 U14410 ( .A(n35973), .Y(n25970) );
  BUFX2 U14411 ( .A(n35973), .Y(n25969) );
  BUFX2 U14412 ( .A(n35973), .Y(n25968) );
  BUFX2 U14413 ( .A(n35581), .Y(n25917) );
  BUFX2 U14414 ( .A(n35581), .Y(n25916) );
  BUFX2 U14415 ( .A(n35581), .Y(n25915) );
  BUFX2 U14416 ( .A(n35581), .Y(n25914) );
  BUFX2 U14417 ( .A(n35581), .Y(n25913) );
  BUFX2 U14418 ( .A(n35581), .Y(n25912) );
  BUFX2 U14419 ( .A(n35451), .Y(n25909) );
  BUFX2 U14420 ( .A(n35451), .Y(n25908) );
  BUFX2 U14421 ( .A(n35451), .Y(n25907) );
  BUFX2 U14422 ( .A(n35451), .Y(n25906) );
  BUFX2 U14423 ( .A(n35451), .Y(n25905) );
  BUFX2 U14424 ( .A(n35451), .Y(n25904) );
  BUFX2 U14425 ( .A(n34924), .Y(n25853) );
  BUFX2 U14426 ( .A(n34924), .Y(n25852) );
  BUFX2 U14427 ( .A(n34924), .Y(n25851) );
  BUFX2 U14428 ( .A(n34924), .Y(n25850) );
  BUFX2 U14429 ( .A(n34924), .Y(n25849) );
  BUFX2 U14430 ( .A(n34924), .Y(n25848) );
  BUFX2 U14431 ( .A(n37018), .Y(n26093) );
  BUFX2 U14432 ( .A(n37018), .Y(n26092) );
  BUFX2 U14433 ( .A(n37018), .Y(n26091) );
  BUFX2 U14434 ( .A(n37018), .Y(n26090) );
  BUFX2 U14435 ( .A(n37018), .Y(n26089) );
  BUFX2 U14436 ( .A(n37018), .Y(n26088) );
  BUFX2 U14437 ( .A(n37017), .Y(n26085) );
  BUFX2 U14438 ( .A(n37017), .Y(n26084) );
  BUFX2 U14439 ( .A(n37017), .Y(n26083) );
  BUFX2 U14440 ( .A(n37017), .Y(n26082) );
  BUFX2 U14441 ( .A(n37017), .Y(n26081) );
  BUFX2 U14442 ( .A(n37017), .Y(n26080) );
  BUFX2 U14443 ( .A(n36493), .Y(n26029) );
  BUFX2 U14444 ( .A(n36493), .Y(n26028) );
  BUFX2 U14445 ( .A(n36493), .Y(n26027) );
  BUFX2 U14446 ( .A(n36493), .Y(n26026) );
  BUFX2 U14447 ( .A(n36493), .Y(n26025) );
  BUFX2 U14448 ( .A(n36493), .Y(n26024) );
  BUFX2 U14449 ( .A(n36492), .Y(n26021) );
  BUFX2 U14450 ( .A(n36492), .Y(n26020) );
  BUFX2 U14451 ( .A(n36492), .Y(n26019) );
  BUFX2 U14452 ( .A(n36492), .Y(n26018) );
  BUFX2 U14453 ( .A(n36492), .Y(n26017) );
  BUFX2 U14454 ( .A(n36492), .Y(n26016) );
  BUFX2 U14455 ( .A(n35971), .Y(n25965) );
  BUFX2 U14456 ( .A(n35971), .Y(n25964) );
  BUFX2 U14457 ( .A(n35971), .Y(n25963) );
  BUFX2 U14458 ( .A(n35971), .Y(n25962) );
  BUFX2 U14459 ( .A(n35971), .Y(n25961) );
  BUFX2 U14460 ( .A(n35971), .Y(n25960) );
  BUFX2 U14461 ( .A(n35970), .Y(n25957) );
  BUFX2 U14462 ( .A(n35970), .Y(n25956) );
  BUFX2 U14463 ( .A(n35970), .Y(n25955) );
  BUFX2 U14464 ( .A(n35970), .Y(n25954) );
  BUFX2 U14465 ( .A(n35970), .Y(n25953) );
  BUFX2 U14466 ( .A(n35970), .Y(n25952) );
  BUFX2 U14467 ( .A(n37016), .Y(n26077) );
  BUFX2 U14468 ( .A(n37016), .Y(n26076) );
  BUFX2 U14469 ( .A(n37016), .Y(n26075) );
  BUFX2 U14470 ( .A(n37016), .Y(n26074) );
  BUFX2 U14471 ( .A(n37016), .Y(n26073) );
  BUFX2 U14472 ( .A(n37016), .Y(n26072) );
  BUFX2 U14473 ( .A(n37015), .Y(n26069) );
  BUFX2 U14474 ( .A(n37015), .Y(n26068) );
  BUFX2 U14475 ( .A(n37015), .Y(n26067) );
  BUFX2 U14476 ( .A(n37015), .Y(n26066) );
  BUFX2 U14477 ( .A(n37015), .Y(n26065) );
  BUFX2 U14478 ( .A(n37015), .Y(n26064) );
  BUFX2 U14479 ( .A(n36887), .Y(n26061) );
  BUFX2 U14480 ( .A(n36887), .Y(n26060) );
  BUFX2 U14481 ( .A(n36887), .Y(n26059) );
  BUFX2 U14482 ( .A(n36887), .Y(n26058) );
  BUFX2 U14483 ( .A(n36887), .Y(n26057) );
  BUFX2 U14484 ( .A(n36887), .Y(n26056) );
  BUFX2 U14485 ( .A(n36758), .Y(n26053) );
  BUFX2 U14486 ( .A(n36758), .Y(n26052) );
  BUFX2 U14487 ( .A(n36758), .Y(n26051) );
  BUFX2 U14488 ( .A(n36758), .Y(n26050) );
  BUFX2 U14489 ( .A(n36758), .Y(n26049) );
  BUFX2 U14490 ( .A(n36758), .Y(n26048) );
  BUFX2 U14491 ( .A(n36491), .Y(n26013) );
  BUFX2 U14492 ( .A(n36491), .Y(n26012) );
  BUFX2 U14493 ( .A(n36491), .Y(n26011) );
  BUFX2 U14494 ( .A(n36491), .Y(n26010) );
  BUFX2 U14495 ( .A(n36491), .Y(n26009) );
  BUFX2 U14496 ( .A(n36491), .Y(n26008) );
  BUFX2 U14497 ( .A(n36490), .Y(n26005) );
  BUFX2 U14498 ( .A(n36490), .Y(n26004) );
  BUFX2 U14499 ( .A(n36490), .Y(n26003) );
  BUFX2 U14500 ( .A(n36490), .Y(n26002) );
  BUFX2 U14501 ( .A(n36490), .Y(n26001) );
  BUFX2 U14502 ( .A(n36490), .Y(n26000) );
  BUFX2 U14503 ( .A(n36362), .Y(n25997) );
  BUFX2 U14504 ( .A(n36362), .Y(n25996) );
  BUFX2 U14505 ( .A(n36362), .Y(n25995) );
  BUFX2 U14506 ( .A(n36362), .Y(n25994) );
  BUFX2 U14507 ( .A(n36362), .Y(n25993) );
  BUFX2 U14508 ( .A(n36362), .Y(n25992) );
  BUFX2 U14509 ( .A(n36233), .Y(n25989) );
  BUFX2 U14510 ( .A(n36233), .Y(n25988) );
  BUFX2 U14511 ( .A(n36233), .Y(n25987) );
  BUFX2 U14512 ( .A(n36233), .Y(n25986) );
  BUFX2 U14513 ( .A(n36233), .Y(n25985) );
  BUFX2 U14514 ( .A(n36233), .Y(n25984) );
  BUFX2 U14515 ( .A(n35969), .Y(n25949) );
  BUFX2 U14516 ( .A(n35969), .Y(n25948) );
  BUFX2 U14517 ( .A(n35969), .Y(n25947) );
  BUFX2 U14518 ( .A(n35969), .Y(n25946) );
  BUFX2 U14519 ( .A(n35969), .Y(n25945) );
  BUFX2 U14520 ( .A(n35969), .Y(n25944) );
  BUFX2 U14521 ( .A(n35968), .Y(n25941) );
  BUFX2 U14522 ( .A(n35968), .Y(n25940) );
  BUFX2 U14523 ( .A(n35968), .Y(n25939) );
  BUFX2 U14524 ( .A(n35968), .Y(n25938) );
  BUFX2 U14525 ( .A(n35968), .Y(n25937) );
  BUFX2 U14526 ( .A(n35968), .Y(n25936) );
  BUFX2 U14527 ( .A(n35840), .Y(n25933) );
  BUFX2 U14528 ( .A(n35840), .Y(n25932) );
  BUFX2 U14529 ( .A(n35840), .Y(n25931) );
  BUFX2 U14530 ( .A(n35840), .Y(n25930) );
  BUFX2 U14531 ( .A(n35840), .Y(n25929) );
  BUFX2 U14532 ( .A(n35840), .Y(n25928) );
  BUFX2 U14533 ( .A(n35711), .Y(n25925) );
  BUFX2 U14534 ( .A(n35711), .Y(n25924) );
  BUFX2 U14535 ( .A(n35711), .Y(n25923) );
  BUFX2 U14536 ( .A(n35711), .Y(n25922) );
  BUFX2 U14537 ( .A(n35711), .Y(n25921) );
  BUFX2 U14538 ( .A(n35711), .Y(n25920) );
  BUFX2 U14539 ( .A(n31539), .Y(n25508) );
  BUFX2 U14540 ( .A(n31541), .Y(n25529) );
  BUFX2 U14541 ( .A(n31567), .Y(n25680) );
  BUFX2 U14542 ( .A(n31569), .Y(n25701) );
  BUFX2 U14543 ( .A(n31580), .Y(n25766) );
  BUFX2 U14544 ( .A(n31582), .Y(n25787) );
  BUFX2 U14545 ( .A(n31539), .Y(n25507) );
  BUFX2 U14546 ( .A(n31541), .Y(n25528) );
  BUFX2 U14547 ( .A(n31567), .Y(n25679) );
  BUFX2 U14548 ( .A(n31569), .Y(n25700) );
  BUFX2 U14549 ( .A(n31580), .Y(n25765) );
  BUFX2 U14550 ( .A(n31582), .Y(n25786) );
  BUFX2 U14551 ( .A(n31539), .Y(n25514) );
  BUFX2 U14552 ( .A(n31541), .Y(n25535) );
  BUFX2 U14553 ( .A(n31567), .Y(n25686) );
  BUFX2 U14554 ( .A(n31569), .Y(n25707) );
  BUFX2 U14555 ( .A(n31580), .Y(n25772) );
  BUFX2 U14556 ( .A(n31582), .Y(n25793) );
  BUFX2 U14557 ( .A(n31539), .Y(n25513) );
  BUFX2 U14558 ( .A(n31541), .Y(n25534) );
  BUFX2 U14559 ( .A(n31567), .Y(n25685) );
  BUFX2 U14560 ( .A(n31569), .Y(n25706) );
  BUFX2 U14561 ( .A(n31580), .Y(n25771) );
  BUFX2 U14562 ( .A(n31582), .Y(n25792) );
  BUFX2 U14563 ( .A(n31539), .Y(n25512) );
  BUFX2 U14564 ( .A(n31541), .Y(n25533) );
  BUFX2 U14565 ( .A(n31567), .Y(n25684) );
  BUFX2 U14566 ( .A(n31569), .Y(n25705) );
  BUFX2 U14567 ( .A(n31580), .Y(n25770) );
  BUFX2 U14568 ( .A(n31582), .Y(n25791) );
  BUFX2 U14569 ( .A(n31539), .Y(n25511) );
  BUFX2 U14570 ( .A(n31541), .Y(n25532) );
  BUFX2 U14571 ( .A(n31567), .Y(n25683) );
  BUFX2 U14572 ( .A(n31569), .Y(n25704) );
  BUFX2 U14573 ( .A(n31580), .Y(n25769) );
  BUFX2 U14574 ( .A(n31582), .Y(n25790) );
  BUFX2 U14575 ( .A(n31539), .Y(n25510) );
  BUFX2 U14576 ( .A(n31541), .Y(n25531) );
  BUFX2 U14577 ( .A(n31567), .Y(n25682) );
  BUFX2 U14578 ( .A(n31569), .Y(n25703) );
  BUFX2 U14579 ( .A(n31580), .Y(n25768) );
  BUFX2 U14580 ( .A(n31582), .Y(n25789) );
  BUFX2 U14581 ( .A(n31539), .Y(n25509) );
  BUFX2 U14582 ( .A(n31541), .Y(n25530) );
  BUFX2 U14583 ( .A(n31567), .Y(n25681) );
  BUFX2 U14584 ( .A(n31569), .Y(n25702) );
  BUFX2 U14585 ( .A(n31580), .Y(n25767) );
  BUFX2 U14586 ( .A(n31582), .Y(n25788) );
  BUFX2 U14587 ( .A(n31539), .Y(n25506) );
  BUFX2 U14588 ( .A(n31541), .Y(n25527) );
  BUFX2 U14589 ( .A(n31567), .Y(n25678) );
  BUFX2 U14590 ( .A(n31569), .Y(n25699) );
  BUFX2 U14591 ( .A(n31580), .Y(n25764) );
  BUFX2 U14592 ( .A(n31582), .Y(n25785) );
  BUFX2 U14593 ( .A(n35322), .Y(n25901) );
  BUFX2 U14594 ( .A(n35322), .Y(n25900) );
  BUFX2 U14595 ( .A(n35322), .Y(n25899) );
  BUFX2 U14596 ( .A(n35322), .Y(n25898) );
  BUFX2 U14597 ( .A(n35322), .Y(n25897) );
  BUFX2 U14598 ( .A(n35322), .Y(n25896) );
  BUFX2 U14599 ( .A(n35189), .Y(n25893) );
  BUFX2 U14600 ( .A(n35189), .Y(n25892) );
  BUFX2 U14601 ( .A(n35189), .Y(n25891) );
  BUFX2 U14602 ( .A(n35189), .Y(n25890) );
  BUFX2 U14603 ( .A(n35189), .Y(n25889) );
  BUFX2 U14604 ( .A(n35189), .Y(n25888) );
  BUFX2 U14605 ( .A(n35060), .Y(n25885) );
  BUFX2 U14606 ( .A(n35060), .Y(n25884) );
  BUFX2 U14607 ( .A(n35060), .Y(n25883) );
  BUFX2 U14608 ( .A(n35060), .Y(n25882) );
  BUFX2 U14609 ( .A(n35060), .Y(n25881) );
  BUFX2 U14610 ( .A(n35060), .Y(n25880) );
  BUFX2 U14611 ( .A(n34930), .Y(n25877) );
  BUFX2 U14612 ( .A(n34930), .Y(n25876) );
  BUFX2 U14613 ( .A(n34930), .Y(n25875) );
  BUFX2 U14614 ( .A(n34930), .Y(n25874) );
  BUFX2 U14615 ( .A(n34930), .Y(n25873) );
  BUFX2 U14616 ( .A(n34930), .Y(n25872) );
  BUFX2 U14617 ( .A(n34928), .Y(n25869) );
  BUFX2 U14618 ( .A(n34928), .Y(n25868) );
  BUFX2 U14619 ( .A(n34928), .Y(n25867) );
  BUFX2 U14620 ( .A(n34928), .Y(n25866) );
  BUFX2 U14621 ( .A(n34928), .Y(n25865) );
  BUFX2 U14622 ( .A(n34928), .Y(n25864) );
  BUFX2 U14623 ( .A(n34926), .Y(n25861) );
  BUFX2 U14624 ( .A(n34926), .Y(n25860) );
  BUFX2 U14625 ( .A(n34926), .Y(n25859) );
  BUFX2 U14626 ( .A(n34926), .Y(n25858) );
  BUFX2 U14627 ( .A(n34926), .Y(n25857) );
  BUFX2 U14628 ( .A(n34926), .Y(n25856) );
  BUFX2 U14629 ( .A(n26131), .Y(n25287) );
  BUFX2 U14630 ( .A(n26133), .Y(n25308) );
  BUFX2 U14631 ( .A(n26131), .Y(n25286) );
  BUFX2 U14632 ( .A(n26133), .Y(n25307) );
  BUFX2 U14633 ( .A(n26131), .Y(n25293) );
  BUFX2 U14634 ( .A(n26133), .Y(n25314) );
  BUFX2 U14635 ( .A(n26131), .Y(n25292) );
  BUFX2 U14636 ( .A(n26133), .Y(n25313) );
  BUFX2 U14637 ( .A(n26131), .Y(n25291) );
  BUFX2 U14638 ( .A(n26133), .Y(n25312) );
  BUFX2 U14639 ( .A(n26131), .Y(n25290) );
  BUFX2 U14640 ( .A(n26133), .Y(n25311) );
  BUFX2 U14641 ( .A(n26131), .Y(n25289) );
  BUFX2 U14642 ( .A(n26133), .Y(n25310) );
  BUFX2 U14643 ( .A(n26131), .Y(n25288) );
  BUFX2 U14644 ( .A(n26133), .Y(n25309) );
  BUFX2 U14645 ( .A(n26131), .Y(n25285) );
  BUFX2 U14646 ( .A(n26133), .Y(n25306) );
  BUFX2 U14647 ( .A(n26114), .Y(n25203) );
  BUFX2 U14648 ( .A(n26116), .Y(n25224) );
  BUFX2 U14649 ( .A(n26150), .Y(n25371) );
  BUFX2 U14650 ( .A(n26152), .Y(n25392) );
  BUFX2 U14651 ( .A(n26167), .Y(n25455) );
  BUFX2 U14652 ( .A(n26169), .Y(n25476) );
  BUFX2 U14653 ( .A(n26114), .Y(n25202) );
  BUFX2 U14654 ( .A(n26116), .Y(n25223) );
  BUFX2 U14655 ( .A(n26150), .Y(n25370) );
  BUFX2 U14656 ( .A(n26152), .Y(n25391) );
  BUFX2 U14657 ( .A(n26167), .Y(n25454) );
  BUFX2 U14658 ( .A(n26169), .Y(n25475) );
  BUFX2 U14659 ( .A(n26114), .Y(n25209) );
  BUFX2 U14660 ( .A(n26116), .Y(n25230) );
  BUFX2 U14661 ( .A(n26150), .Y(n25377) );
  BUFX2 U14662 ( .A(n26152), .Y(n25398) );
  BUFX2 U14663 ( .A(n26167), .Y(n25461) );
  BUFX2 U14664 ( .A(n26169), .Y(n25482) );
  BUFX2 U14665 ( .A(n26114), .Y(n25208) );
  BUFX2 U14666 ( .A(n26116), .Y(n25229) );
  BUFX2 U14667 ( .A(n26150), .Y(n25376) );
  BUFX2 U14668 ( .A(n26152), .Y(n25397) );
  BUFX2 U14669 ( .A(n26167), .Y(n25460) );
  BUFX2 U14670 ( .A(n26169), .Y(n25481) );
  BUFX2 U14671 ( .A(n26114), .Y(n25207) );
  BUFX2 U14672 ( .A(n26116), .Y(n25228) );
  BUFX2 U14673 ( .A(n26150), .Y(n25375) );
  BUFX2 U14674 ( .A(n26152), .Y(n25396) );
  BUFX2 U14675 ( .A(n26167), .Y(n25459) );
  BUFX2 U14676 ( .A(n26169), .Y(n25480) );
  BUFX2 U14677 ( .A(n26114), .Y(n25206) );
  BUFX2 U14678 ( .A(n26116), .Y(n25227) );
  BUFX2 U14679 ( .A(n26150), .Y(n25374) );
  BUFX2 U14680 ( .A(n26152), .Y(n25395) );
  BUFX2 U14681 ( .A(n26167), .Y(n25458) );
  BUFX2 U14682 ( .A(n26169), .Y(n25479) );
  BUFX2 U14683 ( .A(n26114), .Y(n25205) );
  BUFX2 U14684 ( .A(n26116), .Y(n25226) );
  BUFX2 U14685 ( .A(n26150), .Y(n25373) );
  BUFX2 U14686 ( .A(n26152), .Y(n25394) );
  BUFX2 U14687 ( .A(n26167), .Y(n25457) );
  BUFX2 U14688 ( .A(n26169), .Y(n25478) );
  BUFX2 U14689 ( .A(n26114), .Y(n25204) );
  BUFX2 U14690 ( .A(n26116), .Y(n25225) );
  BUFX2 U14691 ( .A(n26150), .Y(n25372) );
  BUFX2 U14692 ( .A(n26152), .Y(n25393) );
  BUFX2 U14693 ( .A(n26167), .Y(n25456) );
  BUFX2 U14694 ( .A(n26169), .Y(n25477) );
  BUFX2 U14695 ( .A(n26114), .Y(n25201) );
  BUFX2 U14696 ( .A(n26116), .Y(n25222) );
  BUFX2 U14697 ( .A(n26150), .Y(n25369) );
  BUFX2 U14698 ( .A(n26152), .Y(n25390) );
  BUFX2 U14699 ( .A(n26167), .Y(n25453) );
  BUFX2 U14700 ( .A(n26169), .Y(n25474) );
  BUFX2 U14701 ( .A(n26122), .Y(n25234) );
  BUFX2 U14702 ( .A(n26122), .Y(n25233) );
  BUFX2 U14703 ( .A(n26122), .Y(n25240) );
  BUFX2 U14704 ( .A(n26122), .Y(n25239) );
  BUFX2 U14705 ( .A(n26122), .Y(n25238) );
  BUFX2 U14706 ( .A(n26122), .Y(n25237) );
  BUFX2 U14707 ( .A(n26122), .Y(n25236) );
  BUFX2 U14708 ( .A(n26122), .Y(n25235) );
  BUFX2 U14709 ( .A(n26122), .Y(n25232) );
  BUFX2 U14710 ( .A(n26105), .Y(n25150) );
  BUFX2 U14711 ( .A(n26109), .Y(n25171) );
  BUFX2 U14712 ( .A(n26126), .Y(n25255) );
  BUFX2 U14713 ( .A(n26141), .Y(n25318) );
  BUFX2 U14714 ( .A(n26145), .Y(n25339) );
  BUFX2 U14715 ( .A(n26158), .Y(n25402) );
  BUFX2 U14716 ( .A(n26162), .Y(n25423) );
  BUFX2 U14717 ( .A(n26105), .Y(n25149) );
  BUFX2 U14718 ( .A(n26109), .Y(n25170) );
  BUFX2 U14719 ( .A(n26126), .Y(n25254) );
  BUFX2 U14720 ( .A(n26141), .Y(n25317) );
  BUFX2 U14721 ( .A(n26145), .Y(n25338) );
  BUFX2 U14722 ( .A(n26158), .Y(n25401) );
  BUFX2 U14723 ( .A(n26162), .Y(n25422) );
  BUFX2 U14724 ( .A(n26105), .Y(n25156) );
  BUFX2 U14725 ( .A(n26109), .Y(n25177) );
  BUFX2 U14726 ( .A(n26126), .Y(n25261) );
  BUFX2 U14727 ( .A(n26141), .Y(n25324) );
  BUFX2 U14728 ( .A(n26145), .Y(n25345) );
  BUFX2 U14729 ( .A(n26158), .Y(n25408) );
  BUFX2 U14730 ( .A(n26162), .Y(n25429) );
  BUFX2 U14731 ( .A(n26105), .Y(n25155) );
  BUFX2 U14732 ( .A(n26109), .Y(n25176) );
  BUFX2 U14733 ( .A(n26126), .Y(n25260) );
  BUFX2 U14734 ( .A(n26141), .Y(n25323) );
  BUFX2 U14735 ( .A(n26145), .Y(n25344) );
  BUFX2 U14736 ( .A(n26158), .Y(n25407) );
  BUFX2 U14737 ( .A(n26162), .Y(n25428) );
  BUFX2 U14738 ( .A(n26105), .Y(n25154) );
  BUFX2 U14739 ( .A(n26109), .Y(n25175) );
  BUFX2 U14740 ( .A(n26126), .Y(n25259) );
  BUFX2 U14741 ( .A(n26141), .Y(n25322) );
  BUFX2 U14742 ( .A(n26145), .Y(n25343) );
  BUFX2 U14743 ( .A(n26158), .Y(n25406) );
  BUFX2 U14744 ( .A(n26162), .Y(n25427) );
  BUFX2 U14745 ( .A(n26105), .Y(n25153) );
  BUFX2 U14746 ( .A(n26109), .Y(n25174) );
  BUFX2 U14747 ( .A(n26126), .Y(n25258) );
  BUFX2 U14748 ( .A(n26141), .Y(n25321) );
  BUFX2 U14749 ( .A(n26145), .Y(n25342) );
  BUFX2 U14750 ( .A(n26158), .Y(n25405) );
  BUFX2 U14751 ( .A(n26162), .Y(n25426) );
  BUFX2 U14752 ( .A(n26105), .Y(n25152) );
  BUFX2 U14753 ( .A(n26109), .Y(n25173) );
  BUFX2 U14754 ( .A(n26126), .Y(n25257) );
  BUFX2 U14755 ( .A(n26141), .Y(n25320) );
  BUFX2 U14756 ( .A(n26145), .Y(n25341) );
  BUFX2 U14757 ( .A(n26158), .Y(n25404) );
  BUFX2 U14758 ( .A(n26162), .Y(n25425) );
  BUFX2 U14759 ( .A(n26105), .Y(n25151) );
  BUFX2 U14760 ( .A(n26109), .Y(n25172) );
  BUFX2 U14761 ( .A(n26126), .Y(n25256) );
  BUFX2 U14762 ( .A(n26141), .Y(n25319) );
  BUFX2 U14763 ( .A(n26145), .Y(n25340) );
  BUFX2 U14764 ( .A(n26158), .Y(n25403) );
  BUFX2 U14765 ( .A(n26162), .Y(n25424) );
  BUFX2 U14766 ( .A(n26105), .Y(n25148) );
  BUFX2 U14767 ( .A(n26109), .Y(n25169) );
  BUFX2 U14768 ( .A(n26126), .Y(n25253) );
  BUFX2 U14769 ( .A(n26141), .Y(n25316) );
  BUFX2 U14770 ( .A(n26145), .Y(n25337) );
  BUFX2 U14771 ( .A(n26158), .Y(n25400) );
  BUFX2 U14772 ( .A(n26162), .Y(n25421) );
  BUFX2 U14773 ( .A(n31551), .Y(n25583) );
  BUFX2 U14774 ( .A(n31551), .Y(n25582) );
  BUFX2 U14775 ( .A(n31551), .Y(n25590) );
  BUFX2 U14776 ( .A(n31551), .Y(n25589) );
  BUFX2 U14777 ( .A(n31551), .Y(n25588) );
  BUFX2 U14778 ( .A(n31551), .Y(n25587) );
  BUFX2 U14779 ( .A(n31551), .Y(n25586) );
  BUFX2 U14780 ( .A(n31551), .Y(n25585) );
  BUFX2 U14781 ( .A(n31551), .Y(n25584) );
  BUFX2 U14782 ( .A(n31551), .Y(n25581) );
  BUFX2 U14783 ( .A(n31538), .Y(n25497) );
  BUFX2 U14784 ( .A(n31540), .Y(n25518) );
  BUFX2 U14785 ( .A(n31553), .Y(n25604) );
  BUFX2 U14786 ( .A(n31566), .Y(n25669) );
  BUFX2 U14787 ( .A(n31568), .Y(n25690) );
  BUFX2 U14788 ( .A(n31579), .Y(n25755) );
  BUFX2 U14789 ( .A(n31581), .Y(n25776) );
  BUFX2 U14790 ( .A(n31538), .Y(n25496) );
  BUFX2 U14791 ( .A(n31540), .Y(n25517) );
  BUFX2 U14792 ( .A(n31553), .Y(n25603) );
  BUFX2 U14793 ( .A(n31566), .Y(n25668) );
  BUFX2 U14794 ( .A(n31568), .Y(n25689) );
  BUFX2 U14795 ( .A(n31579), .Y(n25754) );
  BUFX2 U14796 ( .A(n31581), .Y(n25775) );
  BUFX2 U14797 ( .A(n31538), .Y(n25504) );
  BUFX2 U14798 ( .A(n31540), .Y(n25525) );
  BUFX2 U14799 ( .A(n31553), .Y(n25611) );
  BUFX2 U14800 ( .A(n31566), .Y(n25676) );
  BUFX2 U14801 ( .A(n31568), .Y(n25697) );
  BUFX2 U14802 ( .A(n31579), .Y(n25762) );
  BUFX2 U14803 ( .A(n31581), .Y(n25783) );
  BUFX2 U14804 ( .A(n31538), .Y(n25503) );
  BUFX2 U14805 ( .A(n31540), .Y(n25524) );
  BUFX2 U14806 ( .A(n31553), .Y(n25610) );
  BUFX2 U14807 ( .A(n31566), .Y(n25675) );
  BUFX2 U14808 ( .A(n31568), .Y(n25696) );
  BUFX2 U14809 ( .A(n31579), .Y(n25761) );
  BUFX2 U14810 ( .A(n31581), .Y(n25782) );
  BUFX2 U14811 ( .A(n31538), .Y(n25502) );
  BUFX2 U14812 ( .A(n31540), .Y(n25523) );
  BUFX2 U14813 ( .A(n31553), .Y(n25609) );
  BUFX2 U14814 ( .A(n31566), .Y(n25674) );
  BUFX2 U14815 ( .A(n31568), .Y(n25695) );
  BUFX2 U14816 ( .A(n31579), .Y(n25760) );
  BUFX2 U14817 ( .A(n31581), .Y(n25781) );
  BUFX2 U14818 ( .A(n31538), .Y(n25501) );
  BUFX2 U14819 ( .A(n31540), .Y(n25522) );
  BUFX2 U14820 ( .A(n31553), .Y(n25608) );
  BUFX2 U14821 ( .A(n31566), .Y(n25673) );
  BUFX2 U14822 ( .A(n31568), .Y(n25694) );
  BUFX2 U14823 ( .A(n31579), .Y(n25759) );
  BUFX2 U14824 ( .A(n31581), .Y(n25780) );
  BUFX2 U14825 ( .A(n31538), .Y(n25500) );
  BUFX2 U14826 ( .A(n31540), .Y(n25521) );
  BUFX2 U14827 ( .A(n31553), .Y(n25607) );
  BUFX2 U14828 ( .A(n31566), .Y(n25672) );
  BUFX2 U14829 ( .A(n31568), .Y(n25693) );
  BUFX2 U14830 ( .A(n31579), .Y(n25758) );
  BUFX2 U14831 ( .A(n31581), .Y(n25779) );
  BUFX2 U14832 ( .A(n31538), .Y(n25499) );
  BUFX2 U14833 ( .A(n31540), .Y(n25520) );
  BUFX2 U14834 ( .A(n31553), .Y(n25606) );
  BUFX2 U14835 ( .A(n31566), .Y(n25671) );
  BUFX2 U14836 ( .A(n31568), .Y(n25692) );
  BUFX2 U14837 ( .A(n31579), .Y(n25757) );
  BUFX2 U14838 ( .A(n31581), .Y(n25778) );
  BUFX2 U14839 ( .A(n31538), .Y(n25498) );
  BUFX2 U14840 ( .A(n31540), .Y(n25519) );
  BUFX2 U14841 ( .A(n31553), .Y(n25605) );
  BUFX2 U14842 ( .A(n31566), .Y(n25670) );
  BUFX2 U14843 ( .A(n31568), .Y(n25691) );
  BUFX2 U14844 ( .A(n31579), .Y(n25756) );
  BUFX2 U14845 ( .A(n31581), .Y(n25777) );
  BUFX2 U14846 ( .A(n31538), .Y(n25495) );
  BUFX2 U14847 ( .A(n31540), .Y(n25516) );
  BUFX2 U14848 ( .A(n31553), .Y(n25602) );
  BUFX2 U14849 ( .A(n31566), .Y(n25667) );
  BUFX2 U14850 ( .A(n31568), .Y(n25688) );
  BUFX2 U14851 ( .A(n31579), .Y(n25753) );
  BUFX2 U14852 ( .A(n31581), .Y(n25774) );
  BUFX2 U14853 ( .A(n31556), .Y(n25636) );
  BUFX2 U14854 ( .A(n31558), .Y(n25658) );
  BUFX2 U14855 ( .A(n31556), .Y(n25635) );
  BUFX2 U14856 ( .A(n31558), .Y(n25657) );
  BUFX2 U14857 ( .A(n31556), .Y(n25643) );
  BUFX2 U14858 ( .A(n31558), .Y(n25665) );
  BUFX2 U14859 ( .A(n31556), .Y(n25642) );
  BUFX2 U14860 ( .A(n31558), .Y(n25664) );
  BUFX2 U14861 ( .A(n31556), .Y(n25641) );
  BUFX2 U14862 ( .A(n31558), .Y(n25663) );
  BUFX2 U14863 ( .A(n31556), .Y(n25640) );
  BUFX2 U14864 ( .A(n31558), .Y(n25662) );
  BUFX2 U14865 ( .A(n31556), .Y(n25639) );
  BUFX2 U14866 ( .A(n31558), .Y(n25661) );
  BUFX2 U14867 ( .A(n31556), .Y(n25638) );
  BUFX2 U14868 ( .A(n31558), .Y(n25660) );
  BUFX2 U14869 ( .A(n31556), .Y(n25637) );
  BUFX2 U14870 ( .A(n31558), .Y(n25659) );
  BUFX2 U14871 ( .A(n31556), .Y(n25634) );
  BUFX2 U14872 ( .A(n31558), .Y(n25656) );
  BUFX2 U14873 ( .A(n31543), .Y(n25550) );
  BUFX2 U14874 ( .A(n31545), .Y(n25572) );
  BUFX2 U14875 ( .A(n31571), .Y(n25722) );
  BUFX2 U14876 ( .A(n31573), .Y(n25744) );
  BUFX2 U14877 ( .A(n31584), .Y(n25808) );
  BUFX2 U14878 ( .A(n31586), .Y(n25830) );
  BUFX2 U14879 ( .A(n31543), .Y(n25549) );
  BUFX2 U14880 ( .A(n31545), .Y(n25571) );
  BUFX2 U14881 ( .A(n31571), .Y(n25721) );
  BUFX2 U14882 ( .A(n31573), .Y(n25743) );
  BUFX2 U14883 ( .A(n31584), .Y(n25807) );
  BUFX2 U14884 ( .A(n31586), .Y(n25829) );
  BUFX2 U14885 ( .A(n31543), .Y(n25557) );
  BUFX2 U14886 ( .A(n31545), .Y(n25579) );
  BUFX2 U14887 ( .A(n31571), .Y(n25729) );
  BUFX2 U14888 ( .A(n31573), .Y(n25751) );
  BUFX2 U14889 ( .A(n31584), .Y(n25815) );
  BUFX2 U14890 ( .A(n31586), .Y(n25837) );
  BUFX2 U14891 ( .A(n31543), .Y(n25556) );
  BUFX2 U14892 ( .A(n31545), .Y(n25578) );
  BUFX2 U14893 ( .A(n31571), .Y(n25728) );
  BUFX2 U14894 ( .A(n31573), .Y(n25750) );
  BUFX2 U14895 ( .A(n31584), .Y(n25814) );
  BUFX2 U14896 ( .A(n31586), .Y(n25836) );
  BUFX2 U14897 ( .A(n31543), .Y(n25555) );
  BUFX2 U14898 ( .A(n31545), .Y(n25577) );
  BUFX2 U14899 ( .A(n31571), .Y(n25727) );
  BUFX2 U14900 ( .A(n31573), .Y(n25749) );
  BUFX2 U14901 ( .A(n31584), .Y(n25813) );
  BUFX2 U14902 ( .A(n31586), .Y(n25835) );
  BUFX2 U14903 ( .A(n31543), .Y(n25554) );
  BUFX2 U14904 ( .A(n31545), .Y(n25576) );
  BUFX2 U14905 ( .A(n31571), .Y(n25726) );
  BUFX2 U14906 ( .A(n31573), .Y(n25748) );
  BUFX2 U14907 ( .A(n31584), .Y(n25812) );
  BUFX2 U14908 ( .A(n31586), .Y(n25834) );
  BUFX2 U14909 ( .A(n31543), .Y(n25553) );
  BUFX2 U14910 ( .A(n31545), .Y(n25575) );
  BUFX2 U14911 ( .A(n31571), .Y(n25725) );
  BUFX2 U14912 ( .A(n31573), .Y(n25747) );
  BUFX2 U14913 ( .A(n31584), .Y(n25811) );
  BUFX2 U14914 ( .A(n31586), .Y(n25833) );
  BUFX2 U14915 ( .A(n31543), .Y(n25552) );
  BUFX2 U14916 ( .A(n31545), .Y(n25574) );
  BUFX2 U14917 ( .A(n31571), .Y(n25724) );
  BUFX2 U14918 ( .A(n31573), .Y(n25746) );
  BUFX2 U14919 ( .A(n31584), .Y(n25810) );
  BUFX2 U14920 ( .A(n31586), .Y(n25832) );
  BUFX2 U14921 ( .A(n31543), .Y(n25551) );
  BUFX2 U14922 ( .A(n31545), .Y(n25573) );
  BUFX2 U14923 ( .A(n31571), .Y(n25723) );
  BUFX2 U14924 ( .A(n31573), .Y(n25745) );
  BUFX2 U14925 ( .A(n31584), .Y(n25809) );
  BUFX2 U14926 ( .A(n31586), .Y(n25831) );
  BUFX2 U14927 ( .A(n31543), .Y(n25548) );
  BUFX2 U14928 ( .A(n31545), .Y(n25570) );
  BUFX2 U14929 ( .A(n31571), .Y(n25720) );
  BUFX2 U14930 ( .A(n31573), .Y(n25742) );
  BUFX2 U14931 ( .A(n31584), .Y(n25806) );
  BUFX2 U14932 ( .A(n31586), .Y(n25828) );
  BUFX2 U14933 ( .A(n26124), .Y(n25244) );
  BUFX2 U14934 ( .A(n26128), .Y(n25265) );
  BUFX2 U14935 ( .A(n26124), .Y(n25243) );
  BUFX2 U14936 ( .A(n26128), .Y(n25264) );
  BUFX2 U14937 ( .A(n26124), .Y(n25251) );
  BUFX2 U14938 ( .A(n26128), .Y(n25272) );
  BUFX2 U14939 ( .A(n26124), .Y(n25250) );
  BUFX2 U14940 ( .A(n26128), .Y(n25271) );
  BUFX2 U14941 ( .A(n26124), .Y(n25249) );
  BUFX2 U14942 ( .A(n26128), .Y(n25270) );
  BUFX2 U14943 ( .A(n26124), .Y(n25248) );
  BUFX2 U14944 ( .A(n26128), .Y(n25269) );
  BUFX2 U14945 ( .A(n26124), .Y(n25247) );
  BUFX2 U14946 ( .A(n26128), .Y(n25268) );
  BUFX2 U14947 ( .A(n26124), .Y(n25246) );
  BUFX2 U14948 ( .A(n26128), .Y(n25267) );
  BUFX2 U14949 ( .A(n26124), .Y(n25245) );
  BUFX2 U14950 ( .A(n26128), .Y(n25266) );
  BUFX2 U14951 ( .A(n26124), .Y(n25242) );
  BUFX2 U14952 ( .A(n26128), .Y(n25263) );
  BUFX2 U14953 ( .A(n26107), .Y(n25160) );
  BUFX2 U14954 ( .A(n26111), .Y(n25181) );
  BUFX2 U14955 ( .A(n26143), .Y(n25328) );
  BUFX2 U14956 ( .A(n26147), .Y(n25349) );
  BUFX2 U14957 ( .A(n26160), .Y(n25412) );
  BUFX2 U14958 ( .A(n26164), .Y(n25433) );
  BUFX2 U14959 ( .A(n26107), .Y(n25159) );
  BUFX2 U14960 ( .A(n26111), .Y(n25180) );
  BUFX2 U14961 ( .A(n26143), .Y(n25327) );
  BUFX2 U14962 ( .A(n26147), .Y(n25348) );
  BUFX2 U14963 ( .A(n26160), .Y(n25411) );
  BUFX2 U14964 ( .A(n26164), .Y(n25432) );
  BUFX2 U14965 ( .A(n26107), .Y(n25167) );
  BUFX2 U14966 ( .A(n26111), .Y(n25188) );
  BUFX2 U14967 ( .A(n26143), .Y(n25335) );
  BUFX2 U14968 ( .A(n26147), .Y(n25356) );
  BUFX2 U14969 ( .A(n26160), .Y(n25419) );
  BUFX2 U14970 ( .A(n26164), .Y(n25440) );
  BUFX2 U14971 ( .A(n26107), .Y(n25166) );
  BUFX2 U14972 ( .A(n26111), .Y(n25187) );
  BUFX2 U14973 ( .A(n26143), .Y(n25334) );
  BUFX2 U14974 ( .A(n26147), .Y(n25355) );
  BUFX2 U14975 ( .A(n26160), .Y(n25418) );
  BUFX2 U14976 ( .A(n26164), .Y(n25439) );
  BUFX2 U14977 ( .A(n26107), .Y(n25165) );
  BUFX2 U14978 ( .A(n26111), .Y(n25186) );
  BUFX2 U14979 ( .A(n26143), .Y(n25333) );
  BUFX2 U14980 ( .A(n26147), .Y(n25354) );
  BUFX2 U14981 ( .A(n26160), .Y(n25417) );
  BUFX2 U14982 ( .A(n26164), .Y(n25438) );
  BUFX2 U14983 ( .A(n26107), .Y(n25164) );
  BUFX2 U14984 ( .A(n26111), .Y(n25185) );
  BUFX2 U14985 ( .A(n26143), .Y(n25332) );
  BUFX2 U14986 ( .A(n26147), .Y(n25353) );
  BUFX2 U14987 ( .A(n26160), .Y(n25416) );
  BUFX2 U14988 ( .A(n26164), .Y(n25437) );
  BUFX2 U14989 ( .A(n26107), .Y(n25163) );
  BUFX2 U14990 ( .A(n26111), .Y(n25184) );
  BUFX2 U14991 ( .A(n26143), .Y(n25331) );
  BUFX2 U14992 ( .A(n26147), .Y(n25352) );
  BUFX2 U14993 ( .A(n26160), .Y(n25415) );
  BUFX2 U14994 ( .A(n26164), .Y(n25436) );
  BUFX2 U14995 ( .A(n26107), .Y(n25162) );
  BUFX2 U14996 ( .A(n26111), .Y(n25183) );
  BUFX2 U14997 ( .A(n26143), .Y(n25330) );
  BUFX2 U14998 ( .A(n26147), .Y(n25351) );
  BUFX2 U14999 ( .A(n26160), .Y(n25414) );
  BUFX2 U15000 ( .A(n26164), .Y(n25435) );
  BUFX2 U15001 ( .A(n26107), .Y(n25161) );
  BUFX2 U15002 ( .A(n26111), .Y(n25182) );
  BUFX2 U15003 ( .A(n26143), .Y(n25329) );
  BUFX2 U15004 ( .A(n26147), .Y(n25350) );
  BUFX2 U15005 ( .A(n26160), .Y(n25413) );
  BUFX2 U15006 ( .A(n26164), .Y(n25434) );
  BUFX2 U15007 ( .A(n26107), .Y(n25158) );
  BUFX2 U15008 ( .A(n26111), .Y(n25179) );
  BUFX2 U15009 ( .A(n26143), .Y(n25326) );
  BUFX2 U15010 ( .A(n26147), .Y(n25347) );
  BUFX2 U15011 ( .A(n26160), .Y(n25410) );
  BUFX2 U15012 ( .A(n26164), .Y(n25431) );
  BUFX2 U15013 ( .A(n26130), .Y(n25276) );
  BUFX2 U15014 ( .A(n26132), .Y(n25297) );
  BUFX2 U15015 ( .A(n26130), .Y(n25275) );
  BUFX2 U15016 ( .A(n26132), .Y(n25296) );
  BUFX2 U15017 ( .A(n26130), .Y(n25283) );
  BUFX2 U15018 ( .A(n26132), .Y(n25304) );
  BUFX2 U15019 ( .A(n26130), .Y(n25282) );
  BUFX2 U15020 ( .A(n26132), .Y(n25303) );
  BUFX2 U15021 ( .A(n26130), .Y(n25281) );
  BUFX2 U15022 ( .A(n26132), .Y(n25302) );
  BUFX2 U15023 ( .A(n26130), .Y(n25280) );
  BUFX2 U15024 ( .A(n26132), .Y(n25301) );
  BUFX2 U15025 ( .A(n26130), .Y(n25279) );
  BUFX2 U15026 ( .A(n26132), .Y(n25300) );
  BUFX2 U15027 ( .A(n26130), .Y(n25278) );
  BUFX2 U15028 ( .A(n26132), .Y(n25299) );
  BUFX2 U15029 ( .A(n26130), .Y(n25277) );
  BUFX2 U15030 ( .A(n26132), .Y(n25298) );
  BUFX2 U15031 ( .A(n26130), .Y(n25274) );
  BUFX2 U15032 ( .A(n26132), .Y(n25295) );
  BUFX2 U15033 ( .A(n26113), .Y(n25192) );
  BUFX2 U15034 ( .A(n26115), .Y(n25213) );
  BUFX2 U15035 ( .A(n26149), .Y(n25360) );
  BUFX2 U15036 ( .A(n26151), .Y(n25381) );
  BUFX2 U15037 ( .A(n26166), .Y(n25444) );
  BUFX2 U15038 ( .A(n26168), .Y(n25465) );
  BUFX2 U15039 ( .A(n26113), .Y(n25191) );
  BUFX2 U15040 ( .A(n26115), .Y(n25212) );
  BUFX2 U15041 ( .A(n26149), .Y(n25359) );
  BUFX2 U15042 ( .A(n26151), .Y(n25380) );
  BUFX2 U15043 ( .A(n26166), .Y(n25443) );
  BUFX2 U15044 ( .A(n26168), .Y(n25464) );
  BUFX2 U15045 ( .A(n26113), .Y(n25199) );
  BUFX2 U15046 ( .A(n26115), .Y(n25220) );
  BUFX2 U15047 ( .A(n26149), .Y(n25367) );
  BUFX2 U15048 ( .A(n26151), .Y(n25388) );
  BUFX2 U15049 ( .A(n26166), .Y(n25451) );
  BUFX2 U15050 ( .A(n26168), .Y(n25472) );
  BUFX2 U15051 ( .A(n26113), .Y(n25198) );
  BUFX2 U15052 ( .A(n26115), .Y(n25219) );
  BUFX2 U15053 ( .A(n26149), .Y(n25366) );
  BUFX2 U15054 ( .A(n26151), .Y(n25387) );
  BUFX2 U15055 ( .A(n26166), .Y(n25450) );
  BUFX2 U15056 ( .A(n26168), .Y(n25471) );
  BUFX2 U15057 ( .A(n26113), .Y(n25197) );
  BUFX2 U15058 ( .A(n26115), .Y(n25218) );
  BUFX2 U15059 ( .A(n26149), .Y(n25365) );
  BUFX2 U15060 ( .A(n26151), .Y(n25386) );
  BUFX2 U15061 ( .A(n26166), .Y(n25449) );
  BUFX2 U15062 ( .A(n26168), .Y(n25470) );
  BUFX2 U15063 ( .A(n26113), .Y(n25196) );
  BUFX2 U15064 ( .A(n26115), .Y(n25217) );
  BUFX2 U15065 ( .A(n26149), .Y(n25364) );
  BUFX2 U15066 ( .A(n26151), .Y(n25385) );
  BUFX2 U15067 ( .A(n26166), .Y(n25448) );
  BUFX2 U15068 ( .A(n26168), .Y(n25469) );
  BUFX2 U15069 ( .A(n26113), .Y(n25195) );
  BUFX2 U15070 ( .A(n26115), .Y(n25216) );
  BUFX2 U15071 ( .A(n26149), .Y(n25363) );
  BUFX2 U15072 ( .A(n26151), .Y(n25384) );
  BUFX2 U15073 ( .A(n26166), .Y(n25447) );
  BUFX2 U15074 ( .A(n26168), .Y(n25468) );
  BUFX2 U15075 ( .A(n26113), .Y(n25194) );
  BUFX2 U15076 ( .A(n26115), .Y(n25215) );
  BUFX2 U15077 ( .A(n26149), .Y(n25362) );
  BUFX2 U15078 ( .A(n26151), .Y(n25383) );
  BUFX2 U15079 ( .A(n26166), .Y(n25446) );
  BUFX2 U15080 ( .A(n26168), .Y(n25467) );
  BUFX2 U15081 ( .A(n26113), .Y(n25193) );
  BUFX2 U15082 ( .A(n26115), .Y(n25214) );
  BUFX2 U15083 ( .A(n26149), .Y(n25361) );
  BUFX2 U15084 ( .A(n26151), .Y(n25382) );
  BUFX2 U15085 ( .A(n26166), .Y(n25445) );
  BUFX2 U15086 ( .A(n26168), .Y(n25466) );
  BUFX2 U15087 ( .A(n26113), .Y(n25190) );
  BUFX2 U15088 ( .A(n26115), .Y(n25211) );
  BUFX2 U15089 ( .A(n26149), .Y(n25358) );
  BUFX2 U15090 ( .A(n26151), .Y(n25379) );
  BUFX2 U15091 ( .A(n26166), .Y(n25442) );
  BUFX2 U15092 ( .A(n26168), .Y(n25463) );
  BUFX2 U15093 ( .A(n31555), .Y(n25625) );
  BUFX2 U15094 ( .A(n31557), .Y(n25647) );
  BUFX2 U15095 ( .A(n31555), .Y(n25624) );
  BUFX2 U15096 ( .A(n31557), .Y(n25646) );
  BUFX2 U15097 ( .A(n31555), .Y(n25632) );
  BUFX2 U15098 ( .A(n31557), .Y(n25654) );
  BUFX2 U15099 ( .A(n31555), .Y(n25631) );
  BUFX2 U15100 ( .A(n31557), .Y(n25653) );
  BUFX2 U15101 ( .A(n31555), .Y(n25630) );
  BUFX2 U15102 ( .A(n31557), .Y(n25652) );
  BUFX2 U15103 ( .A(n31555), .Y(n25629) );
  BUFX2 U15104 ( .A(n31557), .Y(n25651) );
  BUFX2 U15105 ( .A(n31555), .Y(n25628) );
  BUFX2 U15106 ( .A(n31557), .Y(n25650) );
  BUFX2 U15107 ( .A(n31555), .Y(n25627) );
  BUFX2 U15108 ( .A(n31557), .Y(n25649) );
  BUFX2 U15109 ( .A(n31555), .Y(n25626) );
  BUFX2 U15110 ( .A(n31557), .Y(n25648) );
  BUFX2 U15111 ( .A(n31555), .Y(n25623) );
  BUFX2 U15112 ( .A(n31557), .Y(n25645) );
  BUFX2 U15113 ( .A(n31542), .Y(n25539) );
  BUFX2 U15114 ( .A(n31544), .Y(n25561) );
  BUFX2 U15115 ( .A(n31570), .Y(n25711) );
  BUFX2 U15116 ( .A(n31572), .Y(n25733) );
  BUFX2 U15117 ( .A(n31583), .Y(n25797) );
  BUFX2 U15118 ( .A(n31585), .Y(n25819) );
  BUFX2 U15119 ( .A(n31542), .Y(n25538) );
  BUFX2 U15120 ( .A(n31544), .Y(n25560) );
  BUFX2 U15121 ( .A(n31570), .Y(n25710) );
  BUFX2 U15122 ( .A(n31572), .Y(n25732) );
  BUFX2 U15123 ( .A(n31583), .Y(n25796) );
  BUFX2 U15124 ( .A(n31585), .Y(n25818) );
  BUFX2 U15125 ( .A(n31542), .Y(n25546) );
  BUFX2 U15126 ( .A(n31544), .Y(n25568) );
  BUFX2 U15127 ( .A(n31570), .Y(n25718) );
  BUFX2 U15128 ( .A(n31572), .Y(n25740) );
  BUFX2 U15129 ( .A(n31583), .Y(n25804) );
  BUFX2 U15130 ( .A(n31585), .Y(n25826) );
  BUFX2 U15131 ( .A(n31542), .Y(n25545) );
  BUFX2 U15132 ( .A(n31544), .Y(n25567) );
  BUFX2 U15133 ( .A(n31570), .Y(n25717) );
  BUFX2 U15134 ( .A(n31572), .Y(n25739) );
  BUFX2 U15135 ( .A(n31583), .Y(n25803) );
  BUFX2 U15136 ( .A(n31585), .Y(n25825) );
  BUFX2 U15137 ( .A(n31542), .Y(n25544) );
  BUFX2 U15138 ( .A(n31544), .Y(n25566) );
  BUFX2 U15139 ( .A(n31570), .Y(n25716) );
  BUFX2 U15140 ( .A(n31572), .Y(n25738) );
  BUFX2 U15141 ( .A(n31583), .Y(n25802) );
  BUFX2 U15142 ( .A(n31585), .Y(n25824) );
  BUFX2 U15143 ( .A(n31542), .Y(n25543) );
  BUFX2 U15144 ( .A(n31544), .Y(n25565) );
  BUFX2 U15145 ( .A(n31570), .Y(n25715) );
  BUFX2 U15146 ( .A(n31572), .Y(n25737) );
  BUFX2 U15147 ( .A(n31583), .Y(n25801) );
  BUFX2 U15148 ( .A(n31585), .Y(n25823) );
  BUFX2 U15149 ( .A(n31542), .Y(n25542) );
  BUFX2 U15150 ( .A(n31544), .Y(n25564) );
  BUFX2 U15151 ( .A(n31570), .Y(n25714) );
  BUFX2 U15152 ( .A(n31572), .Y(n25736) );
  BUFX2 U15153 ( .A(n31583), .Y(n25800) );
  BUFX2 U15154 ( .A(n31585), .Y(n25822) );
  BUFX2 U15155 ( .A(n31542), .Y(n25541) );
  BUFX2 U15156 ( .A(n31544), .Y(n25563) );
  BUFX2 U15157 ( .A(n31570), .Y(n25713) );
  BUFX2 U15158 ( .A(n31572), .Y(n25735) );
  BUFX2 U15159 ( .A(n31583), .Y(n25799) );
  BUFX2 U15160 ( .A(n31585), .Y(n25821) );
  BUFX2 U15161 ( .A(n31542), .Y(n25540) );
  BUFX2 U15162 ( .A(n31544), .Y(n25562) );
  BUFX2 U15163 ( .A(n31570), .Y(n25712) );
  BUFX2 U15164 ( .A(n31572), .Y(n25734) );
  BUFX2 U15165 ( .A(n31583), .Y(n25798) );
  BUFX2 U15166 ( .A(n31585), .Y(n25820) );
  BUFX2 U15167 ( .A(n31542), .Y(n25537) );
  BUFX2 U15168 ( .A(n31544), .Y(n25559) );
  BUFX2 U15169 ( .A(n31570), .Y(n25709) );
  BUFX2 U15170 ( .A(n31572), .Y(n25731) );
  BUFX2 U15171 ( .A(n31583), .Y(n25795) );
  BUFX2 U15172 ( .A(n31585), .Y(n25817) );
  BUFX2 U15173 ( .A(n31552), .Y(n25601) );
  BUFX2 U15174 ( .A(n31554), .Y(n25622) );
  BUFX2 U15175 ( .A(n31539), .Y(n25515) );
  BUFX2 U15176 ( .A(n31541), .Y(n25536) );
  BUFX2 U15177 ( .A(n31567), .Y(n25687) );
  BUFX2 U15178 ( .A(n31569), .Y(n25708) );
  BUFX2 U15179 ( .A(n31580), .Y(n25773) );
  BUFX2 U15180 ( .A(n31582), .Y(n25794) );
  BUFX2 U15181 ( .A(n26131), .Y(n25294) );
  BUFX2 U15182 ( .A(n26133), .Y(n25315) );
  BUFX2 U15183 ( .A(n26114), .Y(n25210) );
  BUFX2 U15184 ( .A(n26116), .Y(n25231) );
  BUFX2 U15185 ( .A(n26150), .Y(n25378) );
  BUFX2 U15186 ( .A(n26152), .Y(n25399) );
  BUFX2 U15187 ( .A(n26167), .Y(n25462) );
  BUFX2 U15188 ( .A(n26169), .Y(n25483) );
  BUFX2 U15189 ( .A(n26122), .Y(n25241) );
  BUFX2 U15190 ( .A(n26105), .Y(n25157) );
  BUFX2 U15191 ( .A(n26109), .Y(n25178) );
  BUFX2 U15192 ( .A(n26126), .Y(n25262) );
  BUFX2 U15193 ( .A(n26141), .Y(n25325) );
  BUFX2 U15194 ( .A(n26145), .Y(n25346) );
  BUFX2 U15195 ( .A(n26158), .Y(n25409) );
  BUFX2 U15196 ( .A(n26162), .Y(n25430) );
  BUFX2 U15197 ( .A(n36625), .Y(n26046) );
  BUFX2 U15198 ( .A(n36495), .Y(n26038) );
  BUFX2 U15199 ( .A(n36103), .Y(n25982) );
  BUFX2 U15200 ( .A(n35973), .Y(n25974) );
  BUFX2 U15201 ( .A(n35581), .Y(n25918) );
  BUFX2 U15202 ( .A(n35451), .Y(n25910) );
  BUFX2 U15203 ( .A(n34924), .Y(n25854) );
  BUFX2 U15204 ( .A(n37018), .Y(n26094) );
  BUFX2 U15205 ( .A(n37017), .Y(n26086) );
  BUFX2 U15206 ( .A(n36493), .Y(n26030) );
  BUFX2 U15207 ( .A(n36492), .Y(n26022) );
  BUFX2 U15208 ( .A(n35971), .Y(n25966) );
  BUFX2 U15209 ( .A(n35970), .Y(n25958) );
  BUFX2 U15210 ( .A(n37016), .Y(n26078) );
  BUFX2 U15211 ( .A(n37015), .Y(n26070) );
  BUFX2 U15212 ( .A(n36887), .Y(n26062) );
  BUFX2 U15213 ( .A(n36758), .Y(n26054) );
  BUFX2 U15214 ( .A(n36491), .Y(n26014) );
  BUFX2 U15215 ( .A(n36490), .Y(n26006) );
  BUFX2 U15216 ( .A(n36362), .Y(n25998) );
  BUFX2 U15217 ( .A(n36233), .Y(n25990) );
  BUFX2 U15218 ( .A(n35969), .Y(n25950) );
  BUFX2 U15219 ( .A(n35968), .Y(n25942) );
  BUFX2 U15220 ( .A(n35840), .Y(n25934) );
  BUFX2 U15221 ( .A(n35711), .Y(n25926) );
  BUFX2 U15222 ( .A(n35322), .Y(n25902) );
  BUFX2 U15223 ( .A(n35189), .Y(n25894) );
  BUFX2 U15224 ( .A(n35060), .Y(n25886) );
  BUFX2 U15225 ( .A(n34930), .Y(n25878) );
  BUFX2 U15226 ( .A(n34928), .Y(n25870) );
  BUFX2 U15227 ( .A(n34926), .Y(n25862) );
  BUFX2 U15228 ( .A(n31551), .Y(n25591) );
  BUFX2 U15229 ( .A(n31538), .Y(n25505) );
  BUFX2 U15230 ( .A(n31540), .Y(n25526) );
  BUFX2 U15231 ( .A(n31553), .Y(n25612) );
  BUFX2 U15232 ( .A(n31566), .Y(n25677) );
  BUFX2 U15233 ( .A(n31568), .Y(n25698) );
  BUFX2 U15234 ( .A(n31579), .Y(n25763) );
  BUFX2 U15235 ( .A(n31581), .Y(n25784) );
  BUFX2 U15236 ( .A(n31556), .Y(n25644) );
  BUFX2 U15237 ( .A(n31558), .Y(n25666) );
  BUFX2 U15238 ( .A(n31543), .Y(n25558) );
  BUFX2 U15239 ( .A(n31545), .Y(n25580) );
  BUFX2 U15240 ( .A(n31571), .Y(n25730) );
  BUFX2 U15241 ( .A(n31573), .Y(n25752) );
  BUFX2 U15242 ( .A(n31584), .Y(n25816) );
  BUFX2 U15243 ( .A(n31586), .Y(n25838) );
  BUFX2 U15244 ( .A(n26124), .Y(n25252) );
  BUFX2 U15245 ( .A(n26128), .Y(n25273) );
  BUFX2 U15246 ( .A(n26107), .Y(n25168) );
  BUFX2 U15247 ( .A(n26111), .Y(n25189) );
  BUFX2 U15248 ( .A(n26143), .Y(n25336) );
  BUFX2 U15249 ( .A(n26147), .Y(n25357) );
  BUFX2 U15250 ( .A(n26160), .Y(n25420) );
  BUFX2 U15251 ( .A(n26164), .Y(n25441) );
  BUFX2 U15252 ( .A(n26130), .Y(n25284) );
  BUFX2 U15253 ( .A(n26132), .Y(n25305) );
  BUFX2 U15254 ( .A(n26113), .Y(n25200) );
  BUFX2 U15255 ( .A(n26115), .Y(n25221) );
  BUFX2 U15256 ( .A(n26149), .Y(n25368) );
  BUFX2 U15257 ( .A(n26151), .Y(n25389) );
  BUFX2 U15258 ( .A(n26166), .Y(n25452) );
  BUFX2 U15259 ( .A(n26168), .Y(n25473) );
  BUFX2 U15260 ( .A(n31555), .Y(n25633) );
  BUFX2 U15261 ( .A(n31557), .Y(n25655) );
  BUFX2 U15262 ( .A(n31542), .Y(n25547) );
  BUFX2 U15263 ( .A(n31544), .Y(n25569) );
  BUFX2 U15264 ( .A(n31570), .Y(n25719) );
  BUFX2 U15265 ( .A(n31572), .Y(n25741) );
  BUFX2 U15266 ( .A(n31583), .Y(n25805) );
  BUFX2 U15267 ( .A(n31585), .Y(n25827) );
  BUFX2 U15268 ( .A(n26097), .Y(n25139) );
  BUFX2 U15269 ( .A(n31530), .Y(n25486) );
  BUFX2 U15270 ( .A(n26097), .Y(n25138) );
  BUFX2 U15271 ( .A(n31530), .Y(n25485) );
  BUFX2 U15272 ( .A(n26097), .Y(n25146) );
  BUFX2 U15273 ( .A(n31530), .Y(n25493) );
  BUFX2 U15274 ( .A(n26097), .Y(n25145) );
  BUFX2 U15275 ( .A(n31530), .Y(n25492) );
  BUFX2 U15276 ( .A(n26097), .Y(n25144) );
  BUFX2 U15277 ( .A(n31530), .Y(n25491) );
  BUFX2 U15278 ( .A(n26097), .Y(n25143) );
  BUFX2 U15279 ( .A(n31530), .Y(n25490) );
  BUFX2 U15280 ( .A(n26097), .Y(n25142) );
  BUFX2 U15281 ( .A(n31530), .Y(n25489) );
  BUFX2 U15282 ( .A(n26097), .Y(n25141) );
  BUFX2 U15283 ( .A(n31530), .Y(n25488) );
  BUFX2 U15284 ( .A(n26097), .Y(n25140) );
  BUFX2 U15285 ( .A(n31530), .Y(n25487) );
  BUFX2 U15286 ( .A(n26097), .Y(n25137) );
  BUFX2 U15287 ( .A(n31530), .Y(n25484) );
  BUFX2 U15288 ( .A(n26097), .Y(n25147) );
  BUFX2 U15289 ( .A(n31530), .Y(n25494) );
  AOI21X1 U15290 ( .A(n26095), .B(n26096), .C(n25147), .Y(rd2data1040_9_) );
  NOR2X1 U15291 ( .A(n26098), .B(n26099), .Y(n26096) );
  NAND3X1 U15292 ( .A(n26100), .B(n26101), .C(n26102), .Y(n26099) );
  NOR2X1 U15293 ( .A(n26103), .B(n26104), .Y(n26102) );
  OAI22X1 U15294 ( .A(n25157), .B(n26106), .C(n25168), .D(n26108), .Y(n26104)
         );
  OAI22X1 U15295 ( .A(n25178), .B(n26110), .C(n25189), .D(n26112), .Y(n26103)
         );
  AOI22X1 U15296 ( .A(reg_file[1417]), .B(n25200), .C(reg_file[1289]), .D(
        n25210), .Y(n26101) );
  AOI22X1 U15297 ( .A(reg_file[1161]), .B(n25221), .C(reg_file[1033]), .D(
        n25231), .Y(n26100) );
  NAND3X1 U15298 ( .A(n26117), .B(n26118), .C(n26119), .Y(n26098) );
  NOR2X1 U15299 ( .A(n26120), .B(n26121), .Y(n26119) );
  OAI22X1 U15300 ( .A(n25241), .B(n26123), .C(n25252), .D(n26125), .Y(n26121)
         );
  OAI22X1 U15301 ( .A(n25262), .B(n26127), .C(n25273), .D(n26129), .Y(n26120)
         );
  AOI22X1 U15302 ( .A(reg_file[521]), .B(n25284), .C(reg_file[649]), .D(n25294), .Y(n26118) );
  AOI22X1 U15303 ( .A(reg_file[777]), .B(n25305), .C(reg_file[905]), .D(n25315), .Y(n26117) );
  NOR2X1 U15304 ( .A(n26134), .B(n26135), .Y(n26095) );
  NAND3X1 U15305 ( .A(n26136), .B(n26137), .C(n26138), .Y(n26135) );
  NOR2X1 U15306 ( .A(n26139), .B(n26140), .Y(n26138) );
  OAI22X1 U15307 ( .A(n25325), .B(n26142), .C(n25336), .D(n26144), .Y(n26140)
         );
  OAI22X1 U15308 ( .A(n25346), .B(n26146), .C(n25357), .D(n26148), .Y(n26139)
         );
  AOI22X1 U15309 ( .A(reg_file[3465]), .B(n25368), .C(reg_file[3337]), .D(
        n25378), .Y(n26137) );
  AOI22X1 U15310 ( .A(reg_file[3209]), .B(n25389), .C(reg_file[3081]), .D(
        n25399), .Y(n26136) );
  NAND3X1 U15311 ( .A(n26153), .B(n26154), .C(n26155), .Y(n26134) );
  NOR2X1 U15312 ( .A(n26156), .B(n26157), .Y(n26155) );
  OAI22X1 U15313 ( .A(n25409), .B(n26159), .C(n25420), .D(n26161), .Y(n26157)
         );
  OAI22X1 U15314 ( .A(n25430), .B(n26163), .C(n25441), .D(n26165), .Y(n26156)
         );
  AOI22X1 U15315 ( .A(reg_file[2441]), .B(n25452), .C(reg_file[2313]), .D(
        n25462), .Y(n26154) );
  AOI22X1 U15316 ( .A(reg_file[2185]), .B(n25473), .C(reg_file[2057]), .D(
        n25483), .Y(n26153) );
  AOI21X1 U15317 ( .A(n26170), .B(n26171), .C(n25147), .Y(rd2data1040_99_) );
  NOR2X1 U15318 ( .A(n26172), .B(n26173), .Y(n26171) );
  NAND3X1 U15319 ( .A(n26174), .B(n26175), .C(n26176), .Y(n26173) );
  NOR2X1 U15320 ( .A(n26177), .B(n26178), .Y(n26176) );
  OAI22X1 U15321 ( .A(n25157), .B(n26179), .C(n25168), .D(n26180), .Y(n26178)
         );
  OAI22X1 U15322 ( .A(n25178), .B(n26181), .C(n25189), .D(n26182), .Y(n26177)
         );
  AOI22X1 U15323 ( .A(reg_file[1507]), .B(n25200), .C(reg_file[1379]), .D(
        n25210), .Y(n26175) );
  AOI22X1 U15324 ( .A(reg_file[1251]), .B(n25221), .C(reg_file[1123]), .D(
        n25231), .Y(n26174) );
  NAND3X1 U15325 ( .A(n26183), .B(n26184), .C(n26185), .Y(n26172) );
  NOR2X1 U15326 ( .A(n26186), .B(n26187), .Y(n26185) );
  OAI22X1 U15327 ( .A(n25241), .B(n26188), .C(n25252), .D(n26189), .Y(n26187)
         );
  OAI22X1 U15328 ( .A(n25262), .B(n26190), .C(n25273), .D(n26191), .Y(n26186)
         );
  AOI22X1 U15329 ( .A(reg_file[611]), .B(n25284), .C(reg_file[739]), .D(n25294), .Y(n26184) );
  AOI22X1 U15330 ( .A(reg_file[867]), .B(n25305), .C(reg_file[995]), .D(n25315), .Y(n26183) );
  NOR2X1 U15331 ( .A(n26192), .B(n26193), .Y(n26170) );
  NAND3X1 U15332 ( .A(n26194), .B(n26195), .C(n26196), .Y(n26193) );
  NOR2X1 U15333 ( .A(n26197), .B(n26198), .Y(n26196) );
  OAI22X1 U15334 ( .A(n25325), .B(n26199), .C(n25336), .D(n26200), .Y(n26198)
         );
  OAI22X1 U15335 ( .A(n25346), .B(n26201), .C(n25357), .D(n26202), .Y(n26197)
         );
  AOI22X1 U15336 ( .A(reg_file[3555]), .B(n25368), .C(reg_file[3427]), .D(
        n25378), .Y(n26195) );
  AOI22X1 U15337 ( .A(reg_file[3299]), .B(n25389), .C(reg_file[3171]), .D(
        n25399), .Y(n26194) );
  NAND3X1 U15338 ( .A(n26203), .B(n26204), .C(n26205), .Y(n26192) );
  NOR2X1 U15339 ( .A(n26206), .B(n26207), .Y(n26205) );
  OAI22X1 U15340 ( .A(n25409), .B(n26208), .C(n25420), .D(n26209), .Y(n26207)
         );
  OAI22X1 U15341 ( .A(n25430), .B(n26210), .C(n25441), .D(n26211), .Y(n26206)
         );
  AOI22X1 U15342 ( .A(reg_file[2531]), .B(n25452), .C(reg_file[2403]), .D(
        n25462), .Y(n26204) );
  AOI22X1 U15343 ( .A(reg_file[2275]), .B(n25473), .C(reg_file[2147]), .D(
        n25483), .Y(n26203) );
  AOI21X1 U15344 ( .A(n26212), .B(n26213), .C(n25147), .Y(rd2data1040_98_) );
  NOR2X1 U15345 ( .A(n26214), .B(n26215), .Y(n26213) );
  NAND3X1 U15346 ( .A(n26216), .B(n26217), .C(n26218), .Y(n26215) );
  NOR2X1 U15347 ( .A(n26219), .B(n26220), .Y(n26218) );
  OAI22X1 U15348 ( .A(n25157), .B(n26221), .C(n25168), .D(n26222), .Y(n26220)
         );
  OAI22X1 U15349 ( .A(n25178), .B(n26223), .C(n25189), .D(n26224), .Y(n26219)
         );
  AOI22X1 U15350 ( .A(reg_file[1506]), .B(n25200), .C(reg_file[1378]), .D(
        n25210), .Y(n26217) );
  AOI22X1 U15351 ( .A(reg_file[1250]), .B(n25221), .C(reg_file[1122]), .D(
        n25231), .Y(n26216) );
  NAND3X1 U15352 ( .A(n26225), .B(n26226), .C(n26227), .Y(n26214) );
  NOR2X1 U15353 ( .A(n26228), .B(n26229), .Y(n26227) );
  OAI22X1 U15354 ( .A(n25241), .B(n26230), .C(n25252), .D(n26231), .Y(n26229)
         );
  OAI22X1 U15355 ( .A(n25262), .B(n26232), .C(n25273), .D(n26233), .Y(n26228)
         );
  AOI22X1 U15356 ( .A(reg_file[610]), .B(n25284), .C(reg_file[738]), .D(n25294), .Y(n26226) );
  AOI22X1 U15357 ( .A(reg_file[866]), .B(n25305), .C(reg_file[994]), .D(n25315), .Y(n26225) );
  NOR2X1 U15358 ( .A(n26234), .B(n26235), .Y(n26212) );
  NAND3X1 U15359 ( .A(n26236), .B(n26237), .C(n26238), .Y(n26235) );
  NOR2X1 U15360 ( .A(n26239), .B(n26240), .Y(n26238) );
  OAI22X1 U15361 ( .A(n25325), .B(n26241), .C(n25336), .D(n26242), .Y(n26240)
         );
  OAI22X1 U15362 ( .A(n25346), .B(n26243), .C(n25357), .D(n26244), .Y(n26239)
         );
  AOI22X1 U15363 ( .A(reg_file[3554]), .B(n25368), .C(reg_file[3426]), .D(
        n25378), .Y(n26237) );
  AOI22X1 U15364 ( .A(reg_file[3298]), .B(n25389), .C(reg_file[3170]), .D(
        n25399), .Y(n26236) );
  NAND3X1 U15365 ( .A(n26245), .B(n26246), .C(n26247), .Y(n26234) );
  NOR2X1 U15366 ( .A(n26248), .B(n26249), .Y(n26247) );
  OAI22X1 U15367 ( .A(n25409), .B(n26250), .C(n25420), .D(n26251), .Y(n26249)
         );
  OAI22X1 U15368 ( .A(n25430), .B(n26252), .C(n25441), .D(n26253), .Y(n26248)
         );
  AOI22X1 U15369 ( .A(reg_file[2530]), .B(n25452), .C(reg_file[2402]), .D(
        n25462), .Y(n26246) );
  AOI22X1 U15370 ( .A(reg_file[2274]), .B(n25473), .C(reg_file[2146]), .D(
        n25483), .Y(n26245) );
  AOI21X1 U15371 ( .A(n26254), .B(n26255), .C(n25147), .Y(rd2data1040_97_) );
  NOR2X1 U15372 ( .A(n26256), .B(n26257), .Y(n26255) );
  NAND3X1 U15373 ( .A(n26258), .B(n26259), .C(n26260), .Y(n26257) );
  NOR2X1 U15374 ( .A(n26261), .B(n26262), .Y(n26260) );
  OAI22X1 U15375 ( .A(n25157), .B(n26263), .C(n25168), .D(n26264), .Y(n26262)
         );
  OAI22X1 U15376 ( .A(n25178), .B(n26265), .C(n25189), .D(n26266), .Y(n26261)
         );
  AOI22X1 U15377 ( .A(reg_file[1505]), .B(n25200), .C(reg_file[1377]), .D(
        n25210), .Y(n26259) );
  AOI22X1 U15378 ( .A(reg_file[1249]), .B(n25221), .C(reg_file[1121]), .D(
        n25231), .Y(n26258) );
  NAND3X1 U15379 ( .A(n26267), .B(n26268), .C(n26269), .Y(n26256) );
  NOR2X1 U15380 ( .A(n26270), .B(n26271), .Y(n26269) );
  OAI22X1 U15381 ( .A(n25241), .B(n26272), .C(n25252), .D(n26273), .Y(n26271)
         );
  OAI22X1 U15382 ( .A(n25262), .B(n26274), .C(n25273), .D(n26275), .Y(n26270)
         );
  AOI22X1 U15383 ( .A(reg_file[609]), .B(n25284), .C(reg_file[737]), .D(n25294), .Y(n26268) );
  AOI22X1 U15384 ( .A(reg_file[865]), .B(n25305), .C(reg_file[993]), .D(n25315), .Y(n26267) );
  NOR2X1 U15385 ( .A(n26276), .B(n26277), .Y(n26254) );
  NAND3X1 U15386 ( .A(n26278), .B(n26279), .C(n26280), .Y(n26277) );
  NOR2X1 U15387 ( .A(n26281), .B(n26282), .Y(n26280) );
  OAI22X1 U15388 ( .A(n25325), .B(n26283), .C(n25336), .D(n26284), .Y(n26282)
         );
  OAI22X1 U15389 ( .A(n25346), .B(n26285), .C(n25357), .D(n26286), .Y(n26281)
         );
  AOI22X1 U15390 ( .A(reg_file[3553]), .B(n25368), .C(reg_file[3425]), .D(
        n25378), .Y(n26279) );
  AOI22X1 U15391 ( .A(reg_file[3297]), .B(n25389), .C(reg_file[3169]), .D(
        n25399), .Y(n26278) );
  NAND3X1 U15392 ( .A(n26287), .B(n26288), .C(n26289), .Y(n26276) );
  NOR2X1 U15393 ( .A(n26290), .B(n26291), .Y(n26289) );
  OAI22X1 U15394 ( .A(n25409), .B(n26292), .C(n25420), .D(n26293), .Y(n26291)
         );
  OAI22X1 U15395 ( .A(n25430), .B(n26294), .C(n25441), .D(n26295), .Y(n26290)
         );
  AOI22X1 U15396 ( .A(reg_file[2529]), .B(n25452), .C(reg_file[2401]), .D(
        n25462), .Y(n26288) );
  AOI22X1 U15397 ( .A(reg_file[2273]), .B(n25473), .C(reg_file[2145]), .D(
        n25483), .Y(n26287) );
  AOI21X1 U15398 ( .A(n26296), .B(n26297), .C(n25147), .Y(rd2data1040_96_) );
  NOR2X1 U15399 ( .A(n26298), .B(n26299), .Y(n26297) );
  NAND3X1 U15400 ( .A(n26300), .B(n26301), .C(n26302), .Y(n26299) );
  NOR2X1 U15401 ( .A(n26303), .B(n26304), .Y(n26302) );
  OAI22X1 U15402 ( .A(n25157), .B(n26305), .C(n25168), .D(n26306), .Y(n26304)
         );
  OAI22X1 U15403 ( .A(n25178), .B(n26307), .C(n25189), .D(n26308), .Y(n26303)
         );
  AOI22X1 U15404 ( .A(reg_file[1504]), .B(n25200), .C(reg_file[1376]), .D(
        n25210), .Y(n26301) );
  AOI22X1 U15405 ( .A(reg_file[1248]), .B(n25221), .C(reg_file[1120]), .D(
        n25231), .Y(n26300) );
  NAND3X1 U15406 ( .A(n26309), .B(n26310), .C(n26311), .Y(n26298) );
  NOR2X1 U15407 ( .A(n26312), .B(n26313), .Y(n26311) );
  OAI22X1 U15408 ( .A(n25241), .B(n26314), .C(n25252), .D(n26315), .Y(n26313)
         );
  OAI22X1 U15409 ( .A(n25262), .B(n26316), .C(n25273), .D(n26317), .Y(n26312)
         );
  AOI22X1 U15410 ( .A(reg_file[608]), .B(n25284), .C(reg_file[736]), .D(n25294), .Y(n26310) );
  AOI22X1 U15411 ( .A(reg_file[864]), .B(n25305), .C(reg_file[992]), .D(n25315), .Y(n26309) );
  NOR2X1 U15412 ( .A(n26318), .B(n26319), .Y(n26296) );
  NAND3X1 U15413 ( .A(n26320), .B(n26321), .C(n26322), .Y(n26319) );
  NOR2X1 U15414 ( .A(n26323), .B(n26324), .Y(n26322) );
  OAI22X1 U15415 ( .A(n25325), .B(n26325), .C(n25336), .D(n26326), .Y(n26324)
         );
  OAI22X1 U15416 ( .A(n25346), .B(n26327), .C(n25357), .D(n26328), .Y(n26323)
         );
  AOI22X1 U15417 ( .A(reg_file[3552]), .B(n25368), .C(reg_file[3424]), .D(
        n25378), .Y(n26321) );
  AOI22X1 U15418 ( .A(reg_file[3296]), .B(n25389), .C(reg_file[3168]), .D(
        n25399), .Y(n26320) );
  NAND3X1 U15419 ( .A(n26329), .B(n26330), .C(n26331), .Y(n26318) );
  NOR2X1 U15420 ( .A(n26332), .B(n26333), .Y(n26331) );
  OAI22X1 U15421 ( .A(n25409), .B(n26334), .C(n25420), .D(n26335), .Y(n26333)
         );
  OAI22X1 U15422 ( .A(n25430), .B(n26336), .C(n25441), .D(n26337), .Y(n26332)
         );
  AOI22X1 U15423 ( .A(reg_file[2528]), .B(n25452), .C(reg_file[2400]), .D(
        n25462), .Y(n26330) );
  AOI22X1 U15424 ( .A(reg_file[2272]), .B(n25473), .C(reg_file[2144]), .D(
        n25483), .Y(n26329) );
  AOI21X1 U15425 ( .A(n26338), .B(n26339), .C(n25147), .Y(rd2data1040_95_) );
  NOR2X1 U15426 ( .A(n26340), .B(n26341), .Y(n26339) );
  NAND3X1 U15427 ( .A(n26342), .B(n26343), .C(n26344), .Y(n26341) );
  NOR2X1 U15428 ( .A(n26345), .B(n26346), .Y(n26344) );
  OAI22X1 U15429 ( .A(n25157), .B(n26347), .C(n25168), .D(n26348), .Y(n26346)
         );
  OAI22X1 U15430 ( .A(n25178), .B(n26349), .C(n25189), .D(n26350), .Y(n26345)
         );
  AOI22X1 U15431 ( .A(reg_file[1503]), .B(n25200), .C(reg_file[1375]), .D(
        n25210), .Y(n26343) );
  AOI22X1 U15432 ( .A(reg_file[1247]), .B(n25221), .C(reg_file[1119]), .D(
        n25231), .Y(n26342) );
  NAND3X1 U15433 ( .A(n26351), .B(n26352), .C(n26353), .Y(n26340) );
  NOR2X1 U15434 ( .A(n26354), .B(n26355), .Y(n26353) );
  OAI22X1 U15435 ( .A(n25241), .B(n26356), .C(n25252), .D(n26357), .Y(n26355)
         );
  OAI22X1 U15436 ( .A(n25262), .B(n26358), .C(n25273), .D(n26359), .Y(n26354)
         );
  AOI22X1 U15437 ( .A(reg_file[607]), .B(n25284), .C(reg_file[735]), .D(n25294), .Y(n26352) );
  AOI22X1 U15438 ( .A(reg_file[863]), .B(n25305), .C(reg_file[991]), .D(n25315), .Y(n26351) );
  NOR2X1 U15439 ( .A(n26360), .B(n26361), .Y(n26338) );
  NAND3X1 U15440 ( .A(n26362), .B(n26363), .C(n26364), .Y(n26361) );
  NOR2X1 U15441 ( .A(n26365), .B(n26366), .Y(n26364) );
  OAI22X1 U15442 ( .A(n25325), .B(n26367), .C(n25336), .D(n26368), .Y(n26366)
         );
  OAI22X1 U15443 ( .A(n25346), .B(n26369), .C(n25357), .D(n26370), .Y(n26365)
         );
  AOI22X1 U15444 ( .A(reg_file[3551]), .B(n25368), .C(reg_file[3423]), .D(
        n25378), .Y(n26363) );
  AOI22X1 U15445 ( .A(reg_file[3295]), .B(n25389), .C(reg_file[3167]), .D(
        n25399), .Y(n26362) );
  NAND3X1 U15446 ( .A(n26371), .B(n26372), .C(n26373), .Y(n26360) );
  NOR2X1 U15447 ( .A(n26374), .B(n26375), .Y(n26373) );
  OAI22X1 U15448 ( .A(n25409), .B(n26376), .C(n25420), .D(n26377), .Y(n26375)
         );
  OAI22X1 U15449 ( .A(n25430), .B(n26378), .C(n25441), .D(n26379), .Y(n26374)
         );
  AOI22X1 U15450 ( .A(reg_file[2527]), .B(n25452), .C(reg_file[2399]), .D(
        n25462), .Y(n26372) );
  AOI22X1 U15451 ( .A(reg_file[2271]), .B(n25473), .C(reg_file[2143]), .D(
        n25483), .Y(n26371) );
  AOI21X1 U15452 ( .A(n26380), .B(n26381), .C(n25147), .Y(rd2data1040_94_) );
  NOR2X1 U15453 ( .A(n26382), .B(n26383), .Y(n26381) );
  NAND3X1 U15454 ( .A(n26384), .B(n26385), .C(n26386), .Y(n26383) );
  NOR2X1 U15455 ( .A(n26387), .B(n26388), .Y(n26386) );
  OAI22X1 U15456 ( .A(n25157), .B(n26389), .C(n25168), .D(n26390), .Y(n26388)
         );
  OAI22X1 U15457 ( .A(n25178), .B(n26391), .C(n25189), .D(n26392), .Y(n26387)
         );
  AOI22X1 U15458 ( .A(reg_file[1502]), .B(n25200), .C(reg_file[1374]), .D(
        n25210), .Y(n26385) );
  AOI22X1 U15459 ( .A(reg_file[1246]), .B(n25221), .C(reg_file[1118]), .D(
        n25231), .Y(n26384) );
  NAND3X1 U15460 ( .A(n26393), .B(n26394), .C(n26395), .Y(n26382) );
  NOR2X1 U15461 ( .A(n26396), .B(n26397), .Y(n26395) );
  OAI22X1 U15462 ( .A(n25241), .B(n26398), .C(n25252), .D(n26399), .Y(n26397)
         );
  OAI22X1 U15463 ( .A(n25262), .B(n26400), .C(n25273), .D(n26401), .Y(n26396)
         );
  AOI22X1 U15464 ( .A(reg_file[606]), .B(n25284), .C(reg_file[734]), .D(n25294), .Y(n26394) );
  AOI22X1 U15465 ( .A(reg_file[862]), .B(n25305), .C(reg_file[990]), .D(n25315), .Y(n26393) );
  NOR2X1 U15466 ( .A(n26402), .B(n26403), .Y(n26380) );
  NAND3X1 U15467 ( .A(n26404), .B(n26405), .C(n26406), .Y(n26403) );
  NOR2X1 U15468 ( .A(n26407), .B(n26408), .Y(n26406) );
  OAI22X1 U15469 ( .A(n25325), .B(n26409), .C(n25336), .D(n26410), .Y(n26408)
         );
  OAI22X1 U15470 ( .A(n25346), .B(n26411), .C(n25357), .D(n26412), .Y(n26407)
         );
  AOI22X1 U15471 ( .A(reg_file[3550]), .B(n25368), .C(reg_file[3422]), .D(
        n25378), .Y(n26405) );
  AOI22X1 U15472 ( .A(reg_file[3294]), .B(n25389), .C(reg_file[3166]), .D(
        n25399), .Y(n26404) );
  NAND3X1 U15473 ( .A(n26413), .B(n26414), .C(n26415), .Y(n26402) );
  NOR2X1 U15474 ( .A(n26416), .B(n26417), .Y(n26415) );
  OAI22X1 U15475 ( .A(n25409), .B(n26418), .C(n25420), .D(n26419), .Y(n26417)
         );
  OAI22X1 U15476 ( .A(n25430), .B(n26420), .C(n25441), .D(n26421), .Y(n26416)
         );
  AOI22X1 U15477 ( .A(reg_file[2526]), .B(n25452), .C(reg_file[2398]), .D(
        n25462), .Y(n26414) );
  AOI22X1 U15478 ( .A(reg_file[2270]), .B(n25473), .C(reg_file[2142]), .D(
        n25483), .Y(n26413) );
  AOI21X1 U15479 ( .A(n26422), .B(n26423), .C(n25147), .Y(rd2data1040_93_) );
  NOR2X1 U15480 ( .A(n26424), .B(n26425), .Y(n26423) );
  NAND3X1 U15481 ( .A(n26426), .B(n26427), .C(n26428), .Y(n26425) );
  NOR2X1 U15482 ( .A(n26429), .B(n26430), .Y(n26428) );
  OAI22X1 U15483 ( .A(n25157), .B(n26431), .C(n25168), .D(n26432), .Y(n26430)
         );
  OAI22X1 U15484 ( .A(n25178), .B(n26433), .C(n25189), .D(n26434), .Y(n26429)
         );
  AOI22X1 U15485 ( .A(reg_file[1501]), .B(n25200), .C(reg_file[1373]), .D(
        n25210), .Y(n26427) );
  AOI22X1 U15486 ( .A(reg_file[1245]), .B(n25221), .C(reg_file[1117]), .D(
        n25231), .Y(n26426) );
  NAND3X1 U15487 ( .A(n26435), .B(n26436), .C(n26437), .Y(n26424) );
  NOR2X1 U15488 ( .A(n26438), .B(n26439), .Y(n26437) );
  OAI22X1 U15489 ( .A(n25241), .B(n26440), .C(n25252), .D(n26441), .Y(n26439)
         );
  OAI22X1 U15490 ( .A(n25262), .B(n26442), .C(n25273), .D(n26443), .Y(n26438)
         );
  AOI22X1 U15491 ( .A(reg_file[605]), .B(n25284), .C(reg_file[733]), .D(n25294), .Y(n26436) );
  AOI22X1 U15492 ( .A(reg_file[861]), .B(n25305), .C(reg_file[989]), .D(n25315), .Y(n26435) );
  NOR2X1 U15493 ( .A(n26444), .B(n26445), .Y(n26422) );
  NAND3X1 U15494 ( .A(n26446), .B(n26447), .C(n26448), .Y(n26445) );
  NOR2X1 U15495 ( .A(n26449), .B(n26450), .Y(n26448) );
  OAI22X1 U15496 ( .A(n25325), .B(n26451), .C(n25336), .D(n26452), .Y(n26450)
         );
  OAI22X1 U15497 ( .A(n25346), .B(n26453), .C(n25357), .D(n26454), .Y(n26449)
         );
  AOI22X1 U15498 ( .A(reg_file[3549]), .B(n25368), .C(reg_file[3421]), .D(
        n25378), .Y(n26447) );
  AOI22X1 U15499 ( .A(reg_file[3293]), .B(n25389), .C(reg_file[3165]), .D(
        n25399), .Y(n26446) );
  NAND3X1 U15500 ( .A(n26455), .B(n26456), .C(n26457), .Y(n26444) );
  NOR2X1 U15501 ( .A(n26458), .B(n26459), .Y(n26457) );
  OAI22X1 U15502 ( .A(n25409), .B(n26460), .C(n25420), .D(n26461), .Y(n26459)
         );
  OAI22X1 U15503 ( .A(n25430), .B(n26462), .C(n25441), .D(n26463), .Y(n26458)
         );
  AOI22X1 U15504 ( .A(reg_file[2525]), .B(n25452), .C(reg_file[2397]), .D(
        n25462), .Y(n26456) );
  AOI22X1 U15505 ( .A(reg_file[2269]), .B(n25473), .C(reg_file[2141]), .D(
        n25483), .Y(n26455) );
  AOI21X1 U15506 ( .A(n26464), .B(n26465), .C(n25146), .Y(rd2data1040_92_) );
  NOR2X1 U15507 ( .A(n26466), .B(n26467), .Y(n26465) );
  NAND3X1 U15508 ( .A(n26468), .B(n26469), .C(n26470), .Y(n26467) );
  NOR2X1 U15509 ( .A(n26471), .B(n26472), .Y(n26470) );
  OAI22X1 U15510 ( .A(n25157), .B(n26473), .C(n25167), .D(n26474), .Y(n26472)
         );
  OAI22X1 U15511 ( .A(n25178), .B(n26475), .C(n25188), .D(n26476), .Y(n26471)
         );
  AOI22X1 U15512 ( .A(reg_file[1500]), .B(n25199), .C(reg_file[1372]), .D(
        n25210), .Y(n26469) );
  AOI22X1 U15513 ( .A(reg_file[1244]), .B(n25220), .C(reg_file[1116]), .D(
        n25231), .Y(n26468) );
  NAND3X1 U15514 ( .A(n26477), .B(n26478), .C(n26479), .Y(n26466) );
  NOR2X1 U15515 ( .A(n26480), .B(n26481), .Y(n26479) );
  OAI22X1 U15516 ( .A(n25241), .B(n26482), .C(n25251), .D(n26483), .Y(n26481)
         );
  OAI22X1 U15517 ( .A(n25262), .B(n26484), .C(n25272), .D(n26485), .Y(n26480)
         );
  AOI22X1 U15518 ( .A(reg_file[604]), .B(n25283), .C(reg_file[732]), .D(n25294), .Y(n26478) );
  AOI22X1 U15519 ( .A(reg_file[860]), .B(n25304), .C(reg_file[988]), .D(n25315), .Y(n26477) );
  NOR2X1 U15520 ( .A(n26486), .B(n26487), .Y(n26464) );
  NAND3X1 U15521 ( .A(n26488), .B(n26489), .C(n26490), .Y(n26487) );
  NOR2X1 U15522 ( .A(n26491), .B(n26492), .Y(n26490) );
  OAI22X1 U15523 ( .A(n25325), .B(n26493), .C(n25335), .D(n26494), .Y(n26492)
         );
  OAI22X1 U15524 ( .A(n25346), .B(n26495), .C(n25356), .D(n26496), .Y(n26491)
         );
  AOI22X1 U15525 ( .A(reg_file[3548]), .B(n25367), .C(reg_file[3420]), .D(
        n25378), .Y(n26489) );
  AOI22X1 U15526 ( .A(reg_file[3292]), .B(n25388), .C(reg_file[3164]), .D(
        n25399), .Y(n26488) );
  NAND3X1 U15527 ( .A(n26497), .B(n26498), .C(n26499), .Y(n26486) );
  NOR2X1 U15528 ( .A(n26500), .B(n26501), .Y(n26499) );
  OAI22X1 U15529 ( .A(n25409), .B(n26502), .C(n25419), .D(n26503), .Y(n26501)
         );
  OAI22X1 U15530 ( .A(n25430), .B(n26504), .C(n25440), .D(n26505), .Y(n26500)
         );
  AOI22X1 U15531 ( .A(reg_file[2524]), .B(n25451), .C(reg_file[2396]), .D(
        n25462), .Y(n26498) );
  AOI22X1 U15532 ( .A(reg_file[2268]), .B(n25472), .C(reg_file[2140]), .D(
        n25483), .Y(n26497) );
  AOI21X1 U15533 ( .A(n26506), .B(n26507), .C(n25146), .Y(rd2data1040_91_) );
  NOR2X1 U15534 ( .A(n26508), .B(n26509), .Y(n26507) );
  NAND3X1 U15535 ( .A(n26510), .B(n26511), .C(n26512), .Y(n26509) );
  NOR2X1 U15536 ( .A(n26513), .B(n26514), .Y(n26512) );
  OAI22X1 U15537 ( .A(n25157), .B(n26515), .C(n25167), .D(n26516), .Y(n26514)
         );
  OAI22X1 U15538 ( .A(n25178), .B(n26517), .C(n25188), .D(n26518), .Y(n26513)
         );
  AOI22X1 U15539 ( .A(reg_file[1499]), .B(n25199), .C(reg_file[1371]), .D(
        n25210), .Y(n26511) );
  AOI22X1 U15540 ( .A(reg_file[1243]), .B(n25220), .C(reg_file[1115]), .D(
        n25231), .Y(n26510) );
  NAND3X1 U15541 ( .A(n26519), .B(n26520), .C(n26521), .Y(n26508) );
  NOR2X1 U15542 ( .A(n26522), .B(n26523), .Y(n26521) );
  OAI22X1 U15543 ( .A(n25241), .B(n26524), .C(n25251), .D(n26525), .Y(n26523)
         );
  OAI22X1 U15544 ( .A(n25262), .B(n26526), .C(n25272), .D(n26527), .Y(n26522)
         );
  AOI22X1 U15545 ( .A(reg_file[603]), .B(n25283), .C(reg_file[731]), .D(n25294), .Y(n26520) );
  AOI22X1 U15546 ( .A(reg_file[859]), .B(n25304), .C(reg_file[987]), .D(n25315), .Y(n26519) );
  NOR2X1 U15547 ( .A(n26528), .B(n26529), .Y(n26506) );
  NAND3X1 U15548 ( .A(n26530), .B(n26531), .C(n26532), .Y(n26529) );
  NOR2X1 U15549 ( .A(n26533), .B(n26534), .Y(n26532) );
  OAI22X1 U15550 ( .A(n25325), .B(n26535), .C(n25335), .D(n26536), .Y(n26534)
         );
  OAI22X1 U15551 ( .A(n25346), .B(n26537), .C(n25356), .D(n26538), .Y(n26533)
         );
  AOI22X1 U15552 ( .A(reg_file[3547]), .B(n25367), .C(reg_file[3419]), .D(
        n25378), .Y(n26531) );
  AOI22X1 U15553 ( .A(reg_file[3291]), .B(n25388), .C(reg_file[3163]), .D(
        n25399), .Y(n26530) );
  NAND3X1 U15554 ( .A(n26539), .B(n26540), .C(n26541), .Y(n26528) );
  NOR2X1 U15555 ( .A(n26542), .B(n26543), .Y(n26541) );
  OAI22X1 U15556 ( .A(n25409), .B(n26544), .C(n25419), .D(n26545), .Y(n26543)
         );
  OAI22X1 U15557 ( .A(n25430), .B(n26546), .C(n25440), .D(n26547), .Y(n26542)
         );
  AOI22X1 U15558 ( .A(reg_file[2523]), .B(n25451), .C(reg_file[2395]), .D(
        n25462), .Y(n26540) );
  AOI22X1 U15559 ( .A(reg_file[2267]), .B(n25472), .C(reg_file[2139]), .D(
        n25483), .Y(n26539) );
  AOI21X1 U15560 ( .A(n26548), .B(n26549), .C(n25146), .Y(rd2data1040_90_) );
  NOR2X1 U15561 ( .A(n26550), .B(n26551), .Y(n26549) );
  NAND3X1 U15562 ( .A(n26552), .B(n26553), .C(n26554), .Y(n26551) );
  NOR2X1 U15563 ( .A(n26555), .B(n26556), .Y(n26554) );
  OAI22X1 U15564 ( .A(n25157), .B(n26557), .C(n25167), .D(n26558), .Y(n26556)
         );
  OAI22X1 U15565 ( .A(n25178), .B(n26559), .C(n25188), .D(n26560), .Y(n26555)
         );
  AOI22X1 U15566 ( .A(reg_file[1498]), .B(n25199), .C(reg_file[1370]), .D(
        n25210), .Y(n26553) );
  AOI22X1 U15567 ( .A(reg_file[1242]), .B(n25220), .C(reg_file[1114]), .D(
        n25231), .Y(n26552) );
  NAND3X1 U15568 ( .A(n26561), .B(n26562), .C(n26563), .Y(n26550) );
  NOR2X1 U15569 ( .A(n26564), .B(n26565), .Y(n26563) );
  OAI22X1 U15570 ( .A(n25241), .B(n26566), .C(n25251), .D(n26567), .Y(n26565)
         );
  OAI22X1 U15571 ( .A(n25262), .B(n26568), .C(n25272), .D(n26569), .Y(n26564)
         );
  AOI22X1 U15572 ( .A(reg_file[602]), .B(n25283), .C(reg_file[730]), .D(n25294), .Y(n26562) );
  AOI22X1 U15573 ( .A(reg_file[858]), .B(n25304), .C(reg_file[986]), .D(n25315), .Y(n26561) );
  NOR2X1 U15574 ( .A(n26570), .B(n26571), .Y(n26548) );
  NAND3X1 U15575 ( .A(n26572), .B(n26573), .C(n26574), .Y(n26571) );
  NOR2X1 U15576 ( .A(n26575), .B(n26576), .Y(n26574) );
  OAI22X1 U15577 ( .A(n25325), .B(n26577), .C(n25335), .D(n26578), .Y(n26576)
         );
  OAI22X1 U15578 ( .A(n25346), .B(n26579), .C(n25356), .D(n26580), .Y(n26575)
         );
  AOI22X1 U15579 ( .A(reg_file[3546]), .B(n25367), .C(reg_file[3418]), .D(
        n25378), .Y(n26573) );
  AOI22X1 U15580 ( .A(reg_file[3290]), .B(n25388), .C(reg_file[3162]), .D(
        n25399), .Y(n26572) );
  NAND3X1 U15581 ( .A(n26581), .B(n26582), .C(n26583), .Y(n26570) );
  NOR2X1 U15582 ( .A(n26584), .B(n26585), .Y(n26583) );
  OAI22X1 U15583 ( .A(n25409), .B(n26586), .C(n25419), .D(n26587), .Y(n26585)
         );
  OAI22X1 U15584 ( .A(n25430), .B(n26588), .C(n25440), .D(n26589), .Y(n26584)
         );
  AOI22X1 U15585 ( .A(reg_file[2522]), .B(n25451), .C(reg_file[2394]), .D(
        n25462), .Y(n26582) );
  AOI22X1 U15586 ( .A(reg_file[2266]), .B(n25472), .C(reg_file[2138]), .D(
        n25483), .Y(n26581) );
  AOI21X1 U15587 ( .A(n26590), .B(n26591), .C(n25146), .Y(rd2data1040_8_) );
  NOR2X1 U15588 ( .A(n26592), .B(n26593), .Y(n26591) );
  NAND3X1 U15589 ( .A(n26594), .B(n26595), .C(n26596), .Y(n26593) );
  NOR2X1 U15590 ( .A(n26597), .B(n26598), .Y(n26596) );
  OAI22X1 U15591 ( .A(n25156), .B(n26599), .C(n25167), .D(n26600), .Y(n26598)
         );
  OAI22X1 U15592 ( .A(n25177), .B(n26601), .C(n25188), .D(n26602), .Y(n26597)
         );
  AOI22X1 U15593 ( .A(reg_file[1416]), .B(n25199), .C(reg_file[1288]), .D(
        n25209), .Y(n26595) );
  AOI22X1 U15594 ( .A(reg_file[1160]), .B(n25220), .C(reg_file[1032]), .D(
        n25230), .Y(n26594) );
  NAND3X1 U15595 ( .A(n26603), .B(n26604), .C(n26605), .Y(n26592) );
  NOR2X1 U15596 ( .A(n26606), .B(n26607), .Y(n26605) );
  OAI22X1 U15597 ( .A(n25240), .B(n26608), .C(n25251), .D(n26609), .Y(n26607)
         );
  OAI22X1 U15598 ( .A(n25261), .B(n26610), .C(n25272), .D(n26611), .Y(n26606)
         );
  AOI22X1 U15599 ( .A(reg_file[520]), .B(n25283), .C(reg_file[648]), .D(n25293), .Y(n26604) );
  AOI22X1 U15600 ( .A(reg_file[776]), .B(n25304), .C(reg_file[904]), .D(n25314), .Y(n26603) );
  NOR2X1 U15601 ( .A(n26612), .B(n26613), .Y(n26590) );
  NAND3X1 U15602 ( .A(n26614), .B(n26615), .C(n26616), .Y(n26613) );
  NOR2X1 U15603 ( .A(n26617), .B(n26618), .Y(n26616) );
  OAI22X1 U15604 ( .A(n25324), .B(n26619), .C(n25335), .D(n26620), .Y(n26618)
         );
  OAI22X1 U15605 ( .A(n25345), .B(n26621), .C(n25356), .D(n26622), .Y(n26617)
         );
  AOI22X1 U15606 ( .A(reg_file[3464]), .B(n25367), .C(reg_file[3336]), .D(
        n25377), .Y(n26615) );
  AOI22X1 U15607 ( .A(reg_file[3208]), .B(n25388), .C(reg_file[3080]), .D(
        n25398), .Y(n26614) );
  NAND3X1 U15608 ( .A(n26623), .B(n26624), .C(n26625), .Y(n26612) );
  NOR2X1 U15609 ( .A(n26626), .B(n26627), .Y(n26625) );
  OAI22X1 U15610 ( .A(n25408), .B(n26628), .C(n25419), .D(n26629), .Y(n26627)
         );
  OAI22X1 U15611 ( .A(n25429), .B(n26630), .C(n25440), .D(n26631), .Y(n26626)
         );
  AOI22X1 U15612 ( .A(reg_file[2440]), .B(n25451), .C(reg_file[2312]), .D(
        n25461), .Y(n26624) );
  AOI22X1 U15613 ( .A(reg_file[2184]), .B(n25472), .C(reg_file[2056]), .D(
        n25482), .Y(n26623) );
  AOI21X1 U15614 ( .A(n26632), .B(n26633), .C(n25146), .Y(rd2data1040_89_) );
  NOR2X1 U15615 ( .A(n26634), .B(n26635), .Y(n26633) );
  NAND3X1 U15616 ( .A(n26636), .B(n26637), .C(n26638), .Y(n26635) );
  NOR2X1 U15617 ( .A(n26639), .B(n26640), .Y(n26638) );
  OAI22X1 U15618 ( .A(n25156), .B(n26641), .C(n25167), .D(n26642), .Y(n26640)
         );
  OAI22X1 U15619 ( .A(n25177), .B(n26643), .C(n25188), .D(n26644), .Y(n26639)
         );
  AOI22X1 U15620 ( .A(reg_file[1497]), .B(n25199), .C(reg_file[1369]), .D(
        n25209), .Y(n26637) );
  AOI22X1 U15621 ( .A(reg_file[1241]), .B(n25220), .C(reg_file[1113]), .D(
        n25230), .Y(n26636) );
  NAND3X1 U15622 ( .A(n26645), .B(n26646), .C(n26647), .Y(n26634) );
  NOR2X1 U15623 ( .A(n26648), .B(n26649), .Y(n26647) );
  OAI22X1 U15624 ( .A(n25240), .B(n26650), .C(n25251), .D(n26651), .Y(n26649)
         );
  OAI22X1 U15625 ( .A(n25261), .B(n26652), .C(n25272), .D(n26653), .Y(n26648)
         );
  AOI22X1 U15626 ( .A(reg_file[601]), .B(n25283), .C(reg_file[729]), .D(n25293), .Y(n26646) );
  AOI22X1 U15627 ( .A(reg_file[857]), .B(n25304), .C(reg_file[985]), .D(n25314), .Y(n26645) );
  NOR2X1 U15628 ( .A(n26654), .B(n26655), .Y(n26632) );
  NAND3X1 U15629 ( .A(n26656), .B(n26657), .C(n26658), .Y(n26655) );
  NOR2X1 U15630 ( .A(n26659), .B(n26660), .Y(n26658) );
  OAI22X1 U15631 ( .A(n25324), .B(n26661), .C(n25335), .D(n26662), .Y(n26660)
         );
  OAI22X1 U15632 ( .A(n25345), .B(n26663), .C(n25356), .D(n26664), .Y(n26659)
         );
  AOI22X1 U15633 ( .A(reg_file[3545]), .B(n25367), .C(reg_file[3417]), .D(
        n25377), .Y(n26657) );
  AOI22X1 U15634 ( .A(reg_file[3289]), .B(n25388), .C(reg_file[3161]), .D(
        n25398), .Y(n26656) );
  NAND3X1 U15635 ( .A(n26665), .B(n26666), .C(n26667), .Y(n26654) );
  NOR2X1 U15636 ( .A(n26668), .B(n26669), .Y(n26667) );
  OAI22X1 U15637 ( .A(n25408), .B(n26670), .C(n25419), .D(n26671), .Y(n26669)
         );
  OAI22X1 U15638 ( .A(n25429), .B(n26672), .C(n25440), .D(n26673), .Y(n26668)
         );
  AOI22X1 U15639 ( .A(reg_file[2521]), .B(n25451), .C(reg_file[2393]), .D(
        n25461), .Y(n26666) );
  AOI22X1 U15640 ( .A(reg_file[2265]), .B(n25472), .C(reg_file[2137]), .D(
        n25482), .Y(n26665) );
  AOI21X1 U15641 ( .A(n26674), .B(n26675), .C(n25146), .Y(rd2data1040_88_) );
  NOR2X1 U15642 ( .A(n26676), .B(n26677), .Y(n26675) );
  NAND3X1 U15643 ( .A(n26678), .B(n26679), .C(n26680), .Y(n26677) );
  NOR2X1 U15644 ( .A(n26681), .B(n26682), .Y(n26680) );
  OAI22X1 U15645 ( .A(n25156), .B(n26683), .C(n25167), .D(n26684), .Y(n26682)
         );
  OAI22X1 U15646 ( .A(n25177), .B(n26685), .C(n25188), .D(n26686), .Y(n26681)
         );
  AOI22X1 U15647 ( .A(reg_file[1496]), .B(n25199), .C(reg_file[1368]), .D(
        n25209), .Y(n26679) );
  AOI22X1 U15648 ( .A(reg_file[1240]), .B(n25220), .C(reg_file[1112]), .D(
        n25230), .Y(n26678) );
  NAND3X1 U15649 ( .A(n26687), .B(n26688), .C(n26689), .Y(n26676) );
  NOR2X1 U15650 ( .A(n26690), .B(n26691), .Y(n26689) );
  OAI22X1 U15651 ( .A(n25240), .B(n26692), .C(n25251), .D(n26693), .Y(n26691)
         );
  OAI22X1 U15652 ( .A(n25261), .B(n26694), .C(n25272), .D(n26695), .Y(n26690)
         );
  AOI22X1 U15653 ( .A(reg_file[600]), .B(n25283), .C(reg_file[728]), .D(n25293), .Y(n26688) );
  AOI22X1 U15654 ( .A(reg_file[856]), .B(n25304), .C(reg_file[984]), .D(n25314), .Y(n26687) );
  NOR2X1 U15655 ( .A(n26696), .B(n26697), .Y(n26674) );
  NAND3X1 U15656 ( .A(n26698), .B(n26699), .C(n26700), .Y(n26697) );
  NOR2X1 U15657 ( .A(n26701), .B(n26702), .Y(n26700) );
  OAI22X1 U15658 ( .A(n25324), .B(n26703), .C(n25335), .D(n26704), .Y(n26702)
         );
  OAI22X1 U15659 ( .A(n25345), .B(n26705), .C(n25356), .D(n26706), .Y(n26701)
         );
  AOI22X1 U15660 ( .A(reg_file[3544]), .B(n25367), .C(reg_file[3416]), .D(
        n25377), .Y(n26699) );
  AOI22X1 U15661 ( .A(reg_file[3288]), .B(n25388), .C(reg_file[3160]), .D(
        n25398), .Y(n26698) );
  NAND3X1 U15662 ( .A(n26707), .B(n26708), .C(n26709), .Y(n26696) );
  NOR2X1 U15663 ( .A(n26710), .B(n26711), .Y(n26709) );
  OAI22X1 U15664 ( .A(n25408), .B(n26712), .C(n25419), .D(n26713), .Y(n26711)
         );
  OAI22X1 U15665 ( .A(n25429), .B(n26714), .C(n25440), .D(n26715), .Y(n26710)
         );
  AOI22X1 U15666 ( .A(reg_file[2520]), .B(n25451), .C(reg_file[2392]), .D(
        n25461), .Y(n26708) );
  AOI22X1 U15667 ( .A(reg_file[2264]), .B(n25472), .C(reg_file[2136]), .D(
        n25482), .Y(n26707) );
  AOI21X1 U15668 ( .A(n26716), .B(n26717), .C(n25146), .Y(rd2data1040_87_) );
  NOR2X1 U15669 ( .A(n26718), .B(n26719), .Y(n26717) );
  NAND3X1 U15670 ( .A(n26720), .B(n26721), .C(n26722), .Y(n26719) );
  NOR2X1 U15671 ( .A(n26723), .B(n26724), .Y(n26722) );
  OAI22X1 U15672 ( .A(n25156), .B(n26725), .C(n25167), .D(n26726), .Y(n26724)
         );
  OAI22X1 U15673 ( .A(n25177), .B(n26727), .C(n25188), .D(n26728), .Y(n26723)
         );
  AOI22X1 U15674 ( .A(reg_file[1495]), .B(n25199), .C(reg_file[1367]), .D(
        n25209), .Y(n26721) );
  AOI22X1 U15675 ( .A(reg_file[1239]), .B(n25220), .C(reg_file[1111]), .D(
        n25230), .Y(n26720) );
  NAND3X1 U15676 ( .A(n26729), .B(n26730), .C(n26731), .Y(n26718) );
  NOR2X1 U15677 ( .A(n26732), .B(n26733), .Y(n26731) );
  OAI22X1 U15678 ( .A(n25240), .B(n26734), .C(n25251), .D(n26735), .Y(n26733)
         );
  OAI22X1 U15679 ( .A(n25261), .B(n26736), .C(n25272), .D(n26737), .Y(n26732)
         );
  AOI22X1 U15680 ( .A(reg_file[599]), .B(n25283), .C(reg_file[727]), .D(n25293), .Y(n26730) );
  AOI22X1 U15681 ( .A(reg_file[855]), .B(n25304), .C(reg_file[983]), .D(n25314), .Y(n26729) );
  NOR2X1 U15682 ( .A(n26738), .B(n26739), .Y(n26716) );
  NAND3X1 U15683 ( .A(n26740), .B(n26741), .C(n26742), .Y(n26739) );
  NOR2X1 U15684 ( .A(n26743), .B(n26744), .Y(n26742) );
  OAI22X1 U15685 ( .A(n25324), .B(n26745), .C(n25335), .D(n26746), .Y(n26744)
         );
  OAI22X1 U15686 ( .A(n25345), .B(n26747), .C(n25356), .D(n26748), .Y(n26743)
         );
  AOI22X1 U15687 ( .A(reg_file[3543]), .B(n25367), .C(reg_file[3415]), .D(
        n25377), .Y(n26741) );
  AOI22X1 U15688 ( .A(reg_file[3287]), .B(n25388), .C(reg_file[3159]), .D(
        n25398), .Y(n26740) );
  NAND3X1 U15689 ( .A(n26749), .B(n26750), .C(n26751), .Y(n26738) );
  NOR2X1 U15690 ( .A(n26752), .B(n26753), .Y(n26751) );
  OAI22X1 U15691 ( .A(n25408), .B(n26754), .C(n25419), .D(n26755), .Y(n26753)
         );
  OAI22X1 U15692 ( .A(n25429), .B(n26756), .C(n25440), .D(n26757), .Y(n26752)
         );
  AOI22X1 U15693 ( .A(reg_file[2519]), .B(n25451), .C(reg_file[2391]), .D(
        n25461), .Y(n26750) );
  AOI22X1 U15694 ( .A(reg_file[2263]), .B(n25472), .C(reg_file[2135]), .D(
        n25482), .Y(n26749) );
  AOI21X1 U15695 ( .A(n26758), .B(n26759), .C(n25146), .Y(rd2data1040_86_) );
  NOR2X1 U15696 ( .A(n26760), .B(n26761), .Y(n26759) );
  NAND3X1 U15697 ( .A(n26762), .B(n26763), .C(n26764), .Y(n26761) );
  NOR2X1 U15698 ( .A(n26765), .B(n26766), .Y(n26764) );
  OAI22X1 U15699 ( .A(n25156), .B(n26767), .C(n25167), .D(n26768), .Y(n26766)
         );
  OAI22X1 U15700 ( .A(n25177), .B(n26769), .C(n25188), .D(n26770), .Y(n26765)
         );
  AOI22X1 U15701 ( .A(reg_file[1494]), .B(n25199), .C(reg_file[1366]), .D(
        n25209), .Y(n26763) );
  AOI22X1 U15702 ( .A(reg_file[1238]), .B(n25220), .C(reg_file[1110]), .D(
        n25230), .Y(n26762) );
  NAND3X1 U15703 ( .A(n26771), .B(n26772), .C(n26773), .Y(n26760) );
  NOR2X1 U15704 ( .A(n26774), .B(n26775), .Y(n26773) );
  OAI22X1 U15705 ( .A(n25240), .B(n26776), .C(n25251), .D(n26777), .Y(n26775)
         );
  OAI22X1 U15706 ( .A(n25261), .B(n26778), .C(n25272), .D(n26779), .Y(n26774)
         );
  AOI22X1 U15707 ( .A(reg_file[598]), .B(n25283), .C(reg_file[726]), .D(n25293), .Y(n26772) );
  AOI22X1 U15708 ( .A(reg_file[854]), .B(n25304), .C(reg_file[982]), .D(n25314), .Y(n26771) );
  NOR2X1 U15709 ( .A(n26780), .B(n26781), .Y(n26758) );
  NAND3X1 U15710 ( .A(n26782), .B(n26783), .C(n26784), .Y(n26781) );
  NOR2X1 U15711 ( .A(n26785), .B(n26786), .Y(n26784) );
  OAI22X1 U15712 ( .A(n25324), .B(n26787), .C(n25335), .D(n26788), .Y(n26786)
         );
  OAI22X1 U15713 ( .A(n25345), .B(n26789), .C(n25356), .D(n26790), .Y(n26785)
         );
  AOI22X1 U15714 ( .A(reg_file[3542]), .B(n25367), .C(reg_file[3414]), .D(
        n25377), .Y(n26783) );
  AOI22X1 U15715 ( .A(reg_file[3286]), .B(n25388), .C(reg_file[3158]), .D(
        n25398), .Y(n26782) );
  NAND3X1 U15716 ( .A(n26791), .B(n26792), .C(n26793), .Y(n26780) );
  NOR2X1 U15717 ( .A(n26794), .B(n26795), .Y(n26793) );
  OAI22X1 U15718 ( .A(n25408), .B(n26796), .C(n25419), .D(n26797), .Y(n26795)
         );
  OAI22X1 U15719 ( .A(n25429), .B(n26798), .C(n25440), .D(n26799), .Y(n26794)
         );
  AOI22X1 U15720 ( .A(reg_file[2518]), .B(n25451), .C(reg_file[2390]), .D(
        n25461), .Y(n26792) );
  AOI22X1 U15721 ( .A(reg_file[2262]), .B(n25472), .C(reg_file[2134]), .D(
        n25482), .Y(n26791) );
  AOI21X1 U15722 ( .A(n26800), .B(n26801), .C(n25146), .Y(rd2data1040_85_) );
  NOR2X1 U15723 ( .A(n26802), .B(n26803), .Y(n26801) );
  NAND3X1 U15724 ( .A(n26804), .B(n26805), .C(n26806), .Y(n26803) );
  NOR2X1 U15725 ( .A(n26807), .B(n26808), .Y(n26806) );
  OAI22X1 U15726 ( .A(n25156), .B(n26809), .C(n25167), .D(n26810), .Y(n26808)
         );
  OAI22X1 U15727 ( .A(n25177), .B(n26811), .C(n25188), .D(n26812), .Y(n26807)
         );
  AOI22X1 U15728 ( .A(reg_file[1493]), .B(n25199), .C(reg_file[1365]), .D(
        n25209), .Y(n26805) );
  AOI22X1 U15729 ( .A(reg_file[1237]), .B(n25220), .C(reg_file[1109]), .D(
        n25230), .Y(n26804) );
  NAND3X1 U15730 ( .A(n26813), .B(n26814), .C(n26815), .Y(n26802) );
  NOR2X1 U15731 ( .A(n26816), .B(n26817), .Y(n26815) );
  OAI22X1 U15732 ( .A(n25240), .B(n26818), .C(n25251), .D(n26819), .Y(n26817)
         );
  OAI22X1 U15733 ( .A(n25261), .B(n26820), .C(n25272), .D(n26821), .Y(n26816)
         );
  AOI22X1 U15734 ( .A(reg_file[597]), .B(n25283), .C(reg_file[725]), .D(n25293), .Y(n26814) );
  AOI22X1 U15735 ( .A(reg_file[853]), .B(n25304), .C(reg_file[981]), .D(n25314), .Y(n26813) );
  NOR2X1 U15736 ( .A(n26822), .B(n26823), .Y(n26800) );
  NAND3X1 U15737 ( .A(n26824), .B(n26825), .C(n26826), .Y(n26823) );
  NOR2X1 U15738 ( .A(n26827), .B(n26828), .Y(n26826) );
  OAI22X1 U15739 ( .A(n25324), .B(n26829), .C(n25335), .D(n26830), .Y(n26828)
         );
  OAI22X1 U15740 ( .A(n25345), .B(n26831), .C(n25356), .D(n26832), .Y(n26827)
         );
  AOI22X1 U15741 ( .A(reg_file[3541]), .B(n25367), .C(reg_file[3413]), .D(
        n25377), .Y(n26825) );
  AOI22X1 U15742 ( .A(reg_file[3285]), .B(n25388), .C(reg_file[3157]), .D(
        n25398), .Y(n26824) );
  NAND3X1 U15743 ( .A(n26833), .B(n26834), .C(n26835), .Y(n26822) );
  NOR2X1 U15744 ( .A(n26836), .B(n26837), .Y(n26835) );
  OAI22X1 U15745 ( .A(n25408), .B(n26838), .C(n25419), .D(n26839), .Y(n26837)
         );
  OAI22X1 U15746 ( .A(n25429), .B(n26840), .C(n25440), .D(n26841), .Y(n26836)
         );
  AOI22X1 U15747 ( .A(reg_file[2517]), .B(n25451), .C(reg_file[2389]), .D(
        n25461), .Y(n26834) );
  AOI22X1 U15748 ( .A(reg_file[2261]), .B(n25472), .C(reg_file[2133]), .D(
        n25482), .Y(n26833) );
  AOI21X1 U15749 ( .A(n26842), .B(n26843), .C(n25146), .Y(rd2data1040_84_) );
  NOR2X1 U15750 ( .A(n26844), .B(n26845), .Y(n26843) );
  NAND3X1 U15751 ( .A(n26846), .B(n26847), .C(n26848), .Y(n26845) );
  NOR2X1 U15752 ( .A(n26849), .B(n26850), .Y(n26848) );
  OAI22X1 U15753 ( .A(n25156), .B(n26851), .C(n25167), .D(n26852), .Y(n26850)
         );
  OAI22X1 U15754 ( .A(n25177), .B(n26853), .C(n25188), .D(n26854), .Y(n26849)
         );
  AOI22X1 U15755 ( .A(reg_file[1492]), .B(n25199), .C(reg_file[1364]), .D(
        n25209), .Y(n26847) );
  AOI22X1 U15756 ( .A(reg_file[1236]), .B(n25220), .C(reg_file[1108]), .D(
        n25230), .Y(n26846) );
  NAND3X1 U15757 ( .A(n26855), .B(n26856), .C(n26857), .Y(n26844) );
  NOR2X1 U15758 ( .A(n26858), .B(n26859), .Y(n26857) );
  OAI22X1 U15759 ( .A(n25240), .B(n26860), .C(n25251), .D(n26861), .Y(n26859)
         );
  OAI22X1 U15760 ( .A(n25261), .B(n26862), .C(n25272), .D(n26863), .Y(n26858)
         );
  AOI22X1 U15761 ( .A(reg_file[596]), .B(n25283), .C(reg_file[724]), .D(n25293), .Y(n26856) );
  AOI22X1 U15762 ( .A(reg_file[852]), .B(n25304), .C(reg_file[980]), .D(n25314), .Y(n26855) );
  NOR2X1 U15763 ( .A(n26864), .B(n26865), .Y(n26842) );
  NAND3X1 U15764 ( .A(n26866), .B(n26867), .C(n26868), .Y(n26865) );
  NOR2X1 U15765 ( .A(n26869), .B(n26870), .Y(n26868) );
  OAI22X1 U15766 ( .A(n25324), .B(n26871), .C(n25335), .D(n26872), .Y(n26870)
         );
  OAI22X1 U15767 ( .A(n25345), .B(n26873), .C(n25356), .D(n26874), .Y(n26869)
         );
  AOI22X1 U15768 ( .A(reg_file[3540]), .B(n25367), .C(reg_file[3412]), .D(
        n25377), .Y(n26867) );
  AOI22X1 U15769 ( .A(reg_file[3284]), .B(n25388), .C(reg_file[3156]), .D(
        n25398), .Y(n26866) );
  NAND3X1 U15770 ( .A(n26875), .B(n26876), .C(n26877), .Y(n26864) );
  NOR2X1 U15771 ( .A(n26878), .B(n26879), .Y(n26877) );
  OAI22X1 U15772 ( .A(n25408), .B(n26880), .C(n25419), .D(n26881), .Y(n26879)
         );
  OAI22X1 U15773 ( .A(n25429), .B(n26882), .C(n25440), .D(n26883), .Y(n26878)
         );
  AOI22X1 U15774 ( .A(reg_file[2516]), .B(n25451), .C(reg_file[2388]), .D(
        n25461), .Y(n26876) );
  AOI22X1 U15775 ( .A(reg_file[2260]), .B(n25472), .C(reg_file[2132]), .D(
        n25482), .Y(n26875) );
  AOI21X1 U15776 ( .A(n26884), .B(n26885), .C(n25146), .Y(rd2data1040_83_) );
  NOR2X1 U15777 ( .A(n26886), .B(n26887), .Y(n26885) );
  NAND3X1 U15778 ( .A(n26888), .B(n26889), .C(n26890), .Y(n26887) );
  NOR2X1 U15779 ( .A(n26891), .B(n26892), .Y(n26890) );
  OAI22X1 U15780 ( .A(n25156), .B(n26893), .C(n25167), .D(n26894), .Y(n26892)
         );
  OAI22X1 U15781 ( .A(n25177), .B(n26895), .C(n25188), .D(n26896), .Y(n26891)
         );
  AOI22X1 U15782 ( .A(reg_file[1491]), .B(n25199), .C(reg_file[1363]), .D(
        n25209), .Y(n26889) );
  AOI22X1 U15783 ( .A(reg_file[1235]), .B(n25220), .C(reg_file[1107]), .D(
        n25230), .Y(n26888) );
  NAND3X1 U15784 ( .A(n26897), .B(n26898), .C(n26899), .Y(n26886) );
  NOR2X1 U15785 ( .A(n26900), .B(n26901), .Y(n26899) );
  OAI22X1 U15786 ( .A(n25240), .B(n26902), .C(n25251), .D(n26903), .Y(n26901)
         );
  OAI22X1 U15787 ( .A(n25261), .B(n26904), .C(n25272), .D(n26905), .Y(n26900)
         );
  AOI22X1 U15788 ( .A(reg_file[595]), .B(n25283), .C(reg_file[723]), .D(n25293), .Y(n26898) );
  AOI22X1 U15789 ( .A(reg_file[851]), .B(n25304), .C(reg_file[979]), .D(n25314), .Y(n26897) );
  NOR2X1 U15790 ( .A(n26906), .B(n26907), .Y(n26884) );
  NAND3X1 U15791 ( .A(n26908), .B(n26909), .C(n26910), .Y(n26907) );
  NOR2X1 U15792 ( .A(n26911), .B(n26912), .Y(n26910) );
  OAI22X1 U15793 ( .A(n25324), .B(n26913), .C(n25335), .D(n26914), .Y(n26912)
         );
  OAI22X1 U15794 ( .A(n25345), .B(n26915), .C(n25356), .D(n26916), .Y(n26911)
         );
  AOI22X1 U15795 ( .A(reg_file[3539]), .B(n25367), .C(reg_file[3411]), .D(
        n25377), .Y(n26909) );
  AOI22X1 U15796 ( .A(reg_file[3283]), .B(n25388), .C(reg_file[3155]), .D(
        n25398), .Y(n26908) );
  NAND3X1 U15797 ( .A(n26917), .B(n26918), .C(n26919), .Y(n26906) );
  NOR2X1 U15798 ( .A(n26920), .B(n26921), .Y(n26919) );
  OAI22X1 U15799 ( .A(n25408), .B(n26922), .C(n25419), .D(n26923), .Y(n26921)
         );
  OAI22X1 U15800 ( .A(n25429), .B(n26924), .C(n25440), .D(n26925), .Y(n26920)
         );
  AOI22X1 U15801 ( .A(reg_file[2515]), .B(n25451), .C(reg_file[2387]), .D(
        n25461), .Y(n26918) );
  AOI22X1 U15802 ( .A(reg_file[2259]), .B(n25472), .C(reg_file[2131]), .D(
        n25482), .Y(n26917) );
  AOI21X1 U15803 ( .A(n26926), .B(n26927), .C(n25146), .Y(rd2data1040_82_) );
  NOR2X1 U15804 ( .A(n26928), .B(n26929), .Y(n26927) );
  NAND3X1 U15805 ( .A(n26930), .B(n26931), .C(n26932), .Y(n26929) );
  NOR2X1 U15806 ( .A(n26933), .B(n26934), .Y(n26932) );
  OAI22X1 U15807 ( .A(n25156), .B(n26935), .C(n25167), .D(n26936), .Y(n26934)
         );
  OAI22X1 U15808 ( .A(n25177), .B(n26937), .C(n25188), .D(n26938), .Y(n26933)
         );
  AOI22X1 U15809 ( .A(reg_file[1490]), .B(n25199), .C(reg_file[1362]), .D(
        n25209), .Y(n26931) );
  AOI22X1 U15810 ( .A(reg_file[1234]), .B(n25220), .C(reg_file[1106]), .D(
        n25230), .Y(n26930) );
  NAND3X1 U15811 ( .A(n26939), .B(n26940), .C(n26941), .Y(n26928) );
  NOR2X1 U15812 ( .A(n26942), .B(n26943), .Y(n26941) );
  OAI22X1 U15813 ( .A(n25240), .B(n26944), .C(n25251), .D(n26945), .Y(n26943)
         );
  OAI22X1 U15814 ( .A(n25261), .B(n26946), .C(n25272), .D(n26947), .Y(n26942)
         );
  AOI22X1 U15815 ( .A(reg_file[594]), .B(n25283), .C(reg_file[722]), .D(n25293), .Y(n26940) );
  AOI22X1 U15816 ( .A(reg_file[850]), .B(n25304), .C(reg_file[978]), .D(n25314), .Y(n26939) );
  NOR2X1 U15817 ( .A(n26948), .B(n26949), .Y(n26926) );
  NAND3X1 U15818 ( .A(n26950), .B(n26951), .C(n26952), .Y(n26949) );
  NOR2X1 U15819 ( .A(n26953), .B(n26954), .Y(n26952) );
  OAI22X1 U15820 ( .A(n25324), .B(n26955), .C(n25335), .D(n26956), .Y(n26954)
         );
  OAI22X1 U15821 ( .A(n25345), .B(n26957), .C(n25356), .D(n26958), .Y(n26953)
         );
  AOI22X1 U15822 ( .A(reg_file[3538]), .B(n25367), .C(reg_file[3410]), .D(
        n25377), .Y(n26951) );
  AOI22X1 U15823 ( .A(reg_file[3282]), .B(n25388), .C(reg_file[3154]), .D(
        n25398), .Y(n26950) );
  NAND3X1 U15824 ( .A(n26959), .B(n26960), .C(n26961), .Y(n26948) );
  NOR2X1 U15825 ( .A(n26962), .B(n26963), .Y(n26961) );
  OAI22X1 U15826 ( .A(n25408), .B(n26964), .C(n25419), .D(n26965), .Y(n26963)
         );
  OAI22X1 U15827 ( .A(n25429), .B(n26966), .C(n25440), .D(n26967), .Y(n26962)
         );
  AOI22X1 U15828 ( .A(reg_file[2514]), .B(n25451), .C(reg_file[2386]), .D(
        n25461), .Y(n26960) );
  AOI22X1 U15829 ( .A(reg_file[2258]), .B(n25472), .C(reg_file[2130]), .D(
        n25482), .Y(n26959) );
  AOI21X1 U15830 ( .A(n26968), .B(n26969), .C(n25145), .Y(rd2data1040_81_) );
  NOR2X1 U15831 ( .A(n26970), .B(n26971), .Y(n26969) );
  NAND3X1 U15832 ( .A(n26972), .B(n26973), .C(n26974), .Y(n26971) );
  NOR2X1 U15833 ( .A(n26975), .B(n26976), .Y(n26974) );
  OAI22X1 U15834 ( .A(n25156), .B(n26977), .C(n25166), .D(n26978), .Y(n26976)
         );
  OAI22X1 U15835 ( .A(n25177), .B(n26979), .C(n25187), .D(n26980), .Y(n26975)
         );
  AOI22X1 U15836 ( .A(reg_file[1489]), .B(n25198), .C(reg_file[1361]), .D(
        n25209), .Y(n26973) );
  AOI22X1 U15837 ( .A(reg_file[1233]), .B(n25219), .C(reg_file[1105]), .D(
        n25230), .Y(n26972) );
  NAND3X1 U15838 ( .A(n26981), .B(n26982), .C(n26983), .Y(n26970) );
  NOR2X1 U15839 ( .A(n26984), .B(n26985), .Y(n26983) );
  OAI22X1 U15840 ( .A(n25240), .B(n26986), .C(n25250), .D(n26987), .Y(n26985)
         );
  OAI22X1 U15841 ( .A(n25261), .B(n26988), .C(n25271), .D(n26989), .Y(n26984)
         );
  AOI22X1 U15842 ( .A(reg_file[593]), .B(n25282), .C(reg_file[721]), .D(n25293), .Y(n26982) );
  AOI22X1 U15843 ( .A(reg_file[849]), .B(n25303), .C(reg_file[977]), .D(n25314), .Y(n26981) );
  NOR2X1 U15844 ( .A(n26990), .B(n26991), .Y(n26968) );
  NAND3X1 U15845 ( .A(n26992), .B(n26993), .C(n26994), .Y(n26991) );
  NOR2X1 U15846 ( .A(n26995), .B(n26996), .Y(n26994) );
  OAI22X1 U15847 ( .A(n25324), .B(n26997), .C(n25334), .D(n26998), .Y(n26996)
         );
  OAI22X1 U15848 ( .A(n25345), .B(n26999), .C(n25355), .D(n27000), .Y(n26995)
         );
  AOI22X1 U15849 ( .A(reg_file[3537]), .B(n25366), .C(reg_file[3409]), .D(
        n25377), .Y(n26993) );
  AOI22X1 U15850 ( .A(reg_file[3281]), .B(n25387), .C(reg_file[3153]), .D(
        n25398), .Y(n26992) );
  NAND3X1 U15851 ( .A(n27001), .B(n27002), .C(n27003), .Y(n26990) );
  NOR2X1 U15852 ( .A(n27004), .B(n27005), .Y(n27003) );
  OAI22X1 U15853 ( .A(n25408), .B(n27006), .C(n25418), .D(n27007), .Y(n27005)
         );
  OAI22X1 U15854 ( .A(n25429), .B(n27008), .C(n25439), .D(n27009), .Y(n27004)
         );
  AOI22X1 U15855 ( .A(reg_file[2513]), .B(n25450), .C(reg_file[2385]), .D(
        n25461), .Y(n27002) );
  AOI22X1 U15856 ( .A(reg_file[2257]), .B(n25471), .C(reg_file[2129]), .D(
        n25482), .Y(n27001) );
  AOI21X1 U15857 ( .A(n27010), .B(n27011), .C(n25145), .Y(rd2data1040_80_) );
  NOR2X1 U15858 ( .A(n27012), .B(n27013), .Y(n27011) );
  NAND3X1 U15859 ( .A(n27014), .B(n27015), .C(n27016), .Y(n27013) );
  NOR2X1 U15860 ( .A(n27017), .B(n27018), .Y(n27016) );
  OAI22X1 U15861 ( .A(n25156), .B(n27019), .C(n25166), .D(n27020), .Y(n27018)
         );
  OAI22X1 U15862 ( .A(n25177), .B(n27021), .C(n25187), .D(n27022), .Y(n27017)
         );
  AOI22X1 U15863 ( .A(reg_file[1488]), .B(n25198), .C(reg_file[1360]), .D(
        n25209), .Y(n27015) );
  AOI22X1 U15864 ( .A(reg_file[1232]), .B(n25219), .C(reg_file[1104]), .D(
        n25230), .Y(n27014) );
  NAND3X1 U15865 ( .A(n27023), .B(n27024), .C(n27025), .Y(n27012) );
  NOR2X1 U15866 ( .A(n27026), .B(n27027), .Y(n27025) );
  OAI22X1 U15867 ( .A(n25240), .B(n27028), .C(n25250), .D(n27029), .Y(n27027)
         );
  OAI22X1 U15868 ( .A(n25261), .B(n27030), .C(n25271), .D(n27031), .Y(n27026)
         );
  AOI22X1 U15869 ( .A(reg_file[592]), .B(n25282), .C(reg_file[720]), .D(n25293), .Y(n27024) );
  AOI22X1 U15870 ( .A(reg_file[848]), .B(n25303), .C(reg_file[976]), .D(n25314), .Y(n27023) );
  NOR2X1 U15871 ( .A(n27032), .B(n27033), .Y(n27010) );
  NAND3X1 U15872 ( .A(n27034), .B(n27035), .C(n27036), .Y(n27033) );
  NOR2X1 U15873 ( .A(n27037), .B(n27038), .Y(n27036) );
  OAI22X1 U15874 ( .A(n25324), .B(n27039), .C(n25334), .D(n27040), .Y(n27038)
         );
  OAI22X1 U15875 ( .A(n25345), .B(n27041), .C(n25355), .D(n27042), .Y(n27037)
         );
  AOI22X1 U15876 ( .A(reg_file[3536]), .B(n25366), .C(reg_file[3408]), .D(
        n25377), .Y(n27035) );
  AOI22X1 U15877 ( .A(reg_file[3280]), .B(n25387), .C(reg_file[3152]), .D(
        n25398), .Y(n27034) );
  NAND3X1 U15878 ( .A(n27043), .B(n27044), .C(n27045), .Y(n27032) );
  NOR2X1 U15879 ( .A(n27046), .B(n27047), .Y(n27045) );
  OAI22X1 U15880 ( .A(n25408), .B(n27048), .C(n25418), .D(n27049), .Y(n27047)
         );
  OAI22X1 U15881 ( .A(n25429), .B(n27050), .C(n25439), .D(n27051), .Y(n27046)
         );
  AOI22X1 U15882 ( .A(reg_file[2512]), .B(n25450), .C(reg_file[2384]), .D(
        n25461), .Y(n27044) );
  AOI22X1 U15883 ( .A(reg_file[2256]), .B(n25471), .C(reg_file[2128]), .D(
        n25482), .Y(n27043) );
  AOI21X1 U15884 ( .A(n27052), .B(n27053), .C(n25145), .Y(rd2data1040_7_) );
  NOR2X1 U15885 ( .A(n27054), .B(n27055), .Y(n27053) );
  NAND3X1 U15886 ( .A(n27056), .B(n27057), .C(n27058), .Y(n27055) );
  NOR2X1 U15887 ( .A(n27059), .B(n27060), .Y(n27058) );
  OAI22X1 U15888 ( .A(n25156), .B(n27061), .C(n25166), .D(n27062), .Y(n27060)
         );
  OAI22X1 U15889 ( .A(n25177), .B(n27063), .C(n25187), .D(n27064), .Y(n27059)
         );
  AOI22X1 U15890 ( .A(reg_file[1415]), .B(n25198), .C(reg_file[1287]), .D(
        n25209), .Y(n27057) );
  AOI22X1 U15891 ( .A(reg_file[1159]), .B(n25219), .C(reg_file[1031]), .D(
        n25230), .Y(n27056) );
  NAND3X1 U15892 ( .A(n27065), .B(n27066), .C(n27067), .Y(n27054) );
  NOR2X1 U15893 ( .A(n27068), .B(n27069), .Y(n27067) );
  OAI22X1 U15894 ( .A(n25240), .B(n27070), .C(n25250), .D(n27071), .Y(n27069)
         );
  OAI22X1 U15895 ( .A(n25261), .B(n27072), .C(n25271), .D(n27073), .Y(n27068)
         );
  AOI22X1 U15896 ( .A(reg_file[519]), .B(n25282), .C(reg_file[647]), .D(n25293), .Y(n27066) );
  AOI22X1 U15897 ( .A(reg_file[775]), .B(n25303), .C(reg_file[903]), .D(n25314), .Y(n27065) );
  NOR2X1 U15898 ( .A(n27074), .B(n27075), .Y(n27052) );
  NAND3X1 U15899 ( .A(n27076), .B(n27077), .C(n27078), .Y(n27075) );
  NOR2X1 U15900 ( .A(n27079), .B(n27080), .Y(n27078) );
  OAI22X1 U15901 ( .A(n25324), .B(n27081), .C(n25334), .D(n27082), .Y(n27080)
         );
  OAI22X1 U15902 ( .A(n25345), .B(n27083), .C(n25355), .D(n27084), .Y(n27079)
         );
  AOI22X1 U15903 ( .A(reg_file[3463]), .B(n25366), .C(reg_file[3335]), .D(
        n25377), .Y(n27077) );
  AOI22X1 U15904 ( .A(reg_file[3207]), .B(n25387), .C(reg_file[3079]), .D(
        n25398), .Y(n27076) );
  NAND3X1 U15905 ( .A(n27085), .B(n27086), .C(n27087), .Y(n27074) );
  NOR2X1 U15906 ( .A(n27088), .B(n27089), .Y(n27087) );
  OAI22X1 U15907 ( .A(n25408), .B(n27090), .C(n25418), .D(n27091), .Y(n27089)
         );
  OAI22X1 U15908 ( .A(n25429), .B(n27092), .C(n25439), .D(n27093), .Y(n27088)
         );
  AOI22X1 U15909 ( .A(reg_file[2439]), .B(n25450), .C(reg_file[2311]), .D(
        n25461), .Y(n27086) );
  AOI22X1 U15910 ( .A(reg_file[2183]), .B(n25471), .C(reg_file[2055]), .D(
        n25482), .Y(n27085) );
  AOI21X1 U15911 ( .A(n27094), .B(n27095), .C(n25145), .Y(rd2data1040_79_) );
  NOR2X1 U15912 ( .A(n27096), .B(n27097), .Y(n27095) );
  NAND3X1 U15913 ( .A(n27098), .B(n27099), .C(n27100), .Y(n27097) );
  NOR2X1 U15914 ( .A(n27101), .B(n27102), .Y(n27100) );
  OAI22X1 U15915 ( .A(n25156), .B(n27103), .C(n25166), .D(n27104), .Y(n27102)
         );
  OAI22X1 U15916 ( .A(n25177), .B(n27105), .C(n25187), .D(n27106), .Y(n27101)
         );
  AOI22X1 U15917 ( .A(reg_file[1487]), .B(n25198), .C(reg_file[1359]), .D(
        n25209), .Y(n27099) );
  AOI22X1 U15918 ( .A(reg_file[1231]), .B(n25219), .C(reg_file[1103]), .D(
        n25230), .Y(n27098) );
  NAND3X1 U15919 ( .A(n27107), .B(n27108), .C(n27109), .Y(n27096) );
  NOR2X1 U15920 ( .A(n27110), .B(n27111), .Y(n27109) );
  OAI22X1 U15921 ( .A(n25240), .B(n27112), .C(n25250), .D(n27113), .Y(n27111)
         );
  OAI22X1 U15922 ( .A(n25261), .B(n27114), .C(n25271), .D(n27115), .Y(n27110)
         );
  AOI22X1 U15923 ( .A(reg_file[591]), .B(n25282), .C(reg_file[719]), .D(n25293), .Y(n27108) );
  AOI22X1 U15924 ( .A(reg_file[847]), .B(n25303), .C(reg_file[975]), .D(n25314), .Y(n27107) );
  NOR2X1 U15925 ( .A(n27116), .B(n27117), .Y(n27094) );
  NAND3X1 U15926 ( .A(n27118), .B(n27119), .C(n27120), .Y(n27117) );
  NOR2X1 U15927 ( .A(n27121), .B(n27122), .Y(n27120) );
  OAI22X1 U15928 ( .A(n25324), .B(n27123), .C(n25334), .D(n27124), .Y(n27122)
         );
  OAI22X1 U15929 ( .A(n25345), .B(n27125), .C(n25355), .D(n27126), .Y(n27121)
         );
  AOI22X1 U15930 ( .A(reg_file[3535]), .B(n25366), .C(reg_file[3407]), .D(
        n25377), .Y(n27119) );
  AOI22X1 U15931 ( .A(reg_file[3279]), .B(n25387), .C(reg_file[3151]), .D(
        n25398), .Y(n27118) );
  NAND3X1 U15932 ( .A(n27127), .B(n27128), .C(n27129), .Y(n27116) );
  NOR2X1 U15933 ( .A(n27130), .B(n27131), .Y(n27129) );
  OAI22X1 U15934 ( .A(n25408), .B(n27132), .C(n25418), .D(n27133), .Y(n27131)
         );
  OAI22X1 U15935 ( .A(n25429), .B(n27134), .C(n25439), .D(n27135), .Y(n27130)
         );
  AOI22X1 U15936 ( .A(reg_file[2511]), .B(n25450), .C(reg_file[2383]), .D(
        n25461), .Y(n27128) );
  AOI22X1 U15937 ( .A(reg_file[2255]), .B(n25471), .C(reg_file[2127]), .D(
        n25482), .Y(n27127) );
  AOI21X1 U15938 ( .A(n27136), .B(n27137), .C(n25145), .Y(rd2data1040_78_) );
  NOR2X1 U15939 ( .A(n27138), .B(n27139), .Y(n27137) );
  NAND3X1 U15940 ( .A(n27140), .B(n27141), .C(n27142), .Y(n27139) );
  NOR2X1 U15941 ( .A(n27143), .B(n27144), .Y(n27142) );
  OAI22X1 U15942 ( .A(n25155), .B(n27145), .C(n25166), .D(n27146), .Y(n27144)
         );
  OAI22X1 U15943 ( .A(n25176), .B(n27147), .C(n25187), .D(n27148), .Y(n27143)
         );
  AOI22X1 U15944 ( .A(reg_file[1486]), .B(n25198), .C(reg_file[1358]), .D(
        n25208), .Y(n27141) );
  AOI22X1 U15945 ( .A(reg_file[1230]), .B(n25219), .C(reg_file[1102]), .D(
        n25229), .Y(n27140) );
  NAND3X1 U15946 ( .A(n27149), .B(n27150), .C(n27151), .Y(n27138) );
  NOR2X1 U15947 ( .A(n27152), .B(n27153), .Y(n27151) );
  OAI22X1 U15948 ( .A(n25239), .B(n27154), .C(n25250), .D(n27155), .Y(n27153)
         );
  OAI22X1 U15949 ( .A(n25260), .B(n27156), .C(n25271), .D(n27157), .Y(n27152)
         );
  AOI22X1 U15950 ( .A(reg_file[590]), .B(n25282), .C(reg_file[718]), .D(n25292), .Y(n27150) );
  AOI22X1 U15951 ( .A(reg_file[846]), .B(n25303), .C(reg_file[974]), .D(n25313), .Y(n27149) );
  NOR2X1 U15952 ( .A(n27158), .B(n27159), .Y(n27136) );
  NAND3X1 U15953 ( .A(n27160), .B(n27161), .C(n27162), .Y(n27159) );
  NOR2X1 U15954 ( .A(n27163), .B(n27164), .Y(n27162) );
  OAI22X1 U15955 ( .A(n25323), .B(n27165), .C(n25334), .D(n27166), .Y(n27164)
         );
  OAI22X1 U15956 ( .A(n25344), .B(n27167), .C(n25355), .D(n27168), .Y(n27163)
         );
  AOI22X1 U15957 ( .A(reg_file[3534]), .B(n25366), .C(reg_file[3406]), .D(
        n25376), .Y(n27161) );
  AOI22X1 U15958 ( .A(reg_file[3278]), .B(n25387), .C(reg_file[3150]), .D(
        n25397), .Y(n27160) );
  NAND3X1 U15959 ( .A(n27169), .B(n27170), .C(n27171), .Y(n27158) );
  NOR2X1 U15960 ( .A(n27172), .B(n27173), .Y(n27171) );
  OAI22X1 U15961 ( .A(n25407), .B(n27174), .C(n25418), .D(n27175), .Y(n27173)
         );
  OAI22X1 U15962 ( .A(n25428), .B(n27176), .C(n25439), .D(n27177), .Y(n27172)
         );
  AOI22X1 U15963 ( .A(reg_file[2510]), .B(n25450), .C(reg_file[2382]), .D(
        n25460), .Y(n27170) );
  AOI22X1 U15964 ( .A(reg_file[2254]), .B(n25471), .C(reg_file[2126]), .D(
        n25481), .Y(n27169) );
  AOI21X1 U15965 ( .A(n27178), .B(n27179), .C(n25145), .Y(rd2data1040_77_) );
  NOR2X1 U15966 ( .A(n27180), .B(n27181), .Y(n27179) );
  NAND3X1 U15967 ( .A(n27182), .B(n27183), .C(n27184), .Y(n27181) );
  NOR2X1 U15968 ( .A(n27185), .B(n27186), .Y(n27184) );
  OAI22X1 U15969 ( .A(n25155), .B(n27187), .C(n25166), .D(n27188), .Y(n27186)
         );
  OAI22X1 U15970 ( .A(n25176), .B(n27189), .C(n25187), .D(n27190), .Y(n27185)
         );
  AOI22X1 U15971 ( .A(reg_file[1485]), .B(n25198), .C(reg_file[1357]), .D(
        n25208), .Y(n27183) );
  AOI22X1 U15972 ( .A(reg_file[1229]), .B(n25219), .C(reg_file[1101]), .D(
        n25229), .Y(n27182) );
  NAND3X1 U15973 ( .A(n27191), .B(n27192), .C(n27193), .Y(n27180) );
  NOR2X1 U15974 ( .A(n27194), .B(n27195), .Y(n27193) );
  OAI22X1 U15975 ( .A(n25239), .B(n27196), .C(n25250), .D(n27197), .Y(n27195)
         );
  OAI22X1 U15976 ( .A(n25260), .B(n27198), .C(n25271), .D(n27199), .Y(n27194)
         );
  AOI22X1 U15977 ( .A(reg_file[589]), .B(n25282), .C(reg_file[717]), .D(n25292), .Y(n27192) );
  AOI22X1 U15978 ( .A(reg_file[845]), .B(n25303), .C(reg_file[973]), .D(n25313), .Y(n27191) );
  NOR2X1 U15979 ( .A(n27200), .B(n27201), .Y(n27178) );
  NAND3X1 U15980 ( .A(n27202), .B(n27203), .C(n27204), .Y(n27201) );
  NOR2X1 U15981 ( .A(n27205), .B(n27206), .Y(n27204) );
  OAI22X1 U15982 ( .A(n25323), .B(n27207), .C(n25334), .D(n27208), .Y(n27206)
         );
  OAI22X1 U15983 ( .A(n25344), .B(n27209), .C(n25355), .D(n27210), .Y(n27205)
         );
  AOI22X1 U15984 ( .A(reg_file[3533]), .B(n25366), .C(reg_file[3405]), .D(
        n25376), .Y(n27203) );
  AOI22X1 U15985 ( .A(reg_file[3277]), .B(n25387), .C(reg_file[3149]), .D(
        n25397), .Y(n27202) );
  NAND3X1 U15986 ( .A(n27211), .B(n27212), .C(n27213), .Y(n27200) );
  NOR2X1 U15987 ( .A(n27214), .B(n27215), .Y(n27213) );
  OAI22X1 U15988 ( .A(n25407), .B(n27216), .C(n25418), .D(n27217), .Y(n27215)
         );
  OAI22X1 U15989 ( .A(n25428), .B(n27218), .C(n25439), .D(n27219), .Y(n27214)
         );
  AOI22X1 U15990 ( .A(reg_file[2509]), .B(n25450), .C(reg_file[2381]), .D(
        n25460), .Y(n27212) );
  AOI22X1 U15991 ( .A(reg_file[2253]), .B(n25471), .C(reg_file[2125]), .D(
        n25481), .Y(n27211) );
  AOI21X1 U15992 ( .A(n27220), .B(n27221), .C(n25145), .Y(rd2data1040_76_) );
  NOR2X1 U15993 ( .A(n27222), .B(n27223), .Y(n27221) );
  NAND3X1 U15994 ( .A(n27224), .B(n27225), .C(n27226), .Y(n27223) );
  NOR2X1 U15995 ( .A(n27227), .B(n27228), .Y(n27226) );
  OAI22X1 U15996 ( .A(n25155), .B(n27229), .C(n25166), .D(n27230), .Y(n27228)
         );
  OAI22X1 U15997 ( .A(n25176), .B(n27231), .C(n25187), .D(n27232), .Y(n27227)
         );
  AOI22X1 U15998 ( .A(reg_file[1484]), .B(n25198), .C(reg_file[1356]), .D(
        n25208), .Y(n27225) );
  AOI22X1 U15999 ( .A(reg_file[1228]), .B(n25219), .C(reg_file[1100]), .D(
        n25229), .Y(n27224) );
  NAND3X1 U16000 ( .A(n27233), .B(n27234), .C(n27235), .Y(n27222) );
  NOR2X1 U16001 ( .A(n27236), .B(n27237), .Y(n27235) );
  OAI22X1 U16002 ( .A(n25239), .B(n27238), .C(n25250), .D(n27239), .Y(n27237)
         );
  OAI22X1 U16003 ( .A(n25260), .B(n27240), .C(n25271), .D(n27241), .Y(n27236)
         );
  AOI22X1 U16004 ( .A(reg_file[588]), .B(n25282), .C(reg_file[716]), .D(n25292), .Y(n27234) );
  AOI22X1 U16005 ( .A(reg_file[844]), .B(n25303), .C(reg_file[972]), .D(n25313), .Y(n27233) );
  NOR2X1 U16006 ( .A(n27242), .B(n27243), .Y(n27220) );
  NAND3X1 U16007 ( .A(n27244), .B(n27245), .C(n27246), .Y(n27243) );
  NOR2X1 U16008 ( .A(n27247), .B(n27248), .Y(n27246) );
  OAI22X1 U16009 ( .A(n25323), .B(n27249), .C(n25334), .D(n27250), .Y(n27248)
         );
  OAI22X1 U16010 ( .A(n25344), .B(n27251), .C(n25355), .D(n27252), .Y(n27247)
         );
  AOI22X1 U16011 ( .A(reg_file[3532]), .B(n25366), .C(reg_file[3404]), .D(
        n25376), .Y(n27245) );
  AOI22X1 U16012 ( .A(reg_file[3276]), .B(n25387), .C(reg_file[3148]), .D(
        n25397), .Y(n27244) );
  NAND3X1 U16013 ( .A(n27253), .B(n27254), .C(n27255), .Y(n27242) );
  NOR2X1 U16014 ( .A(n27256), .B(n27257), .Y(n27255) );
  OAI22X1 U16015 ( .A(n25407), .B(n27258), .C(n25418), .D(n27259), .Y(n27257)
         );
  OAI22X1 U16016 ( .A(n25428), .B(n27260), .C(n25439), .D(n27261), .Y(n27256)
         );
  AOI22X1 U16017 ( .A(reg_file[2508]), .B(n25450), .C(reg_file[2380]), .D(
        n25460), .Y(n27254) );
  AOI22X1 U16018 ( .A(reg_file[2252]), .B(n25471), .C(reg_file[2124]), .D(
        n25481), .Y(n27253) );
  AOI21X1 U16019 ( .A(n27262), .B(n27263), .C(n25145), .Y(rd2data1040_75_) );
  NOR2X1 U16020 ( .A(n27264), .B(n27265), .Y(n27263) );
  NAND3X1 U16021 ( .A(n27266), .B(n27267), .C(n27268), .Y(n27265) );
  NOR2X1 U16022 ( .A(n27269), .B(n27270), .Y(n27268) );
  OAI22X1 U16023 ( .A(n25155), .B(n27271), .C(n25166), .D(n27272), .Y(n27270)
         );
  OAI22X1 U16024 ( .A(n25176), .B(n27273), .C(n25187), .D(n27274), .Y(n27269)
         );
  AOI22X1 U16025 ( .A(reg_file[1483]), .B(n25198), .C(reg_file[1355]), .D(
        n25208), .Y(n27267) );
  AOI22X1 U16026 ( .A(reg_file[1227]), .B(n25219), .C(reg_file[1099]), .D(
        n25229), .Y(n27266) );
  NAND3X1 U16027 ( .A(n27275), .B(n27276), .C(n27277), .Y(n27264) );
  NOR2X1 U16028 ( .A(n27278), .B(n27279), .Y(n27277) );
  OAI22X1 U16029 ( .A(n25239), .B(n27280), .C(n25250), .D(n27281), .Y(n27279)
         );
  OAI22X1 U16030 ( .A(n25260), .B(n27282), .C(n25271), .D(n27283), .Y(n27278)
         );
  AOI22X1 U16031 ( .A(reg_file[587]), .B(n25282), .C(reg_file[715]), .D(n25292), .Y(n27276) );
  AOI22X1 U16032 ( .A(reg_file[843]), .B(n25303), .C(reg_file[971]), .D(n25313), .Y(n27275) );
  NOR2X1 U16033 ( .A(n27284), .B(n27285), .Y(n27262) );
  NAND3X1 U16034 ( .A(n27286), .B(n27287), .C(n27288), .Y(n27285) );
  NOR2X1 U16035 ( .A(n27289), .B(n27290), .Y(n27288) );
  OAI22X1 U16036 ( .A(n25323), .B(n27291), .C(n25334), .D(n27292), .Y(n27290)
         );
  OAI22X1 U16037 ( .A(n25344), .B(n27293), .C(n25355), .D(n27294), .Y(n27289)
         );
  AOI22X1 U16038 ( .A(reg_file[3531]), .B(n25366), .C(reg_file[3403]), .D(
        n25376), .Y(n27287) );
  AOI22X1 U16039 ( .A(reg_file[3275]), .B(n25387), .C(reg_file[3147]), .D(
        n25397), .Y(n27286) );
  NAND3X1 U16040 ( .A(n27295), .B(n27296), .C(n27297), .Y(n27284) );
  NOR2X1 U16041 ( .A(n27298), .B(n27299), .Y(n27297) );
  OAI22X1 U16042 ( .A(n25407), .B(n27300), .C(n25418), .D(n27301), .Y(n27299)
         );
  OAI22X1 U16043 ( .A(n25428), .B(n27302), .C(n25439), .D(n27303), .Y(n27298)
         );
  AOI22X1 U16044 ( .A(reg_file[2507]), .B(n25450), .C(reg_file[2379]), .D(
        n25460), .Y(n27296) );
  AOI22X1 U16045 ( .A(reg_file[2251]), .B(n25471), .C(reg_file[2123]), .D(
        n25481), .Y(n27295) );
  AOI21X1 U16046 ( .A(n27304), .B(n27305), .C(n25145), .Y(rd2data1040_74_) );
  NOR2X1 U16047 ( .A(n27306), .B(n27307), .Y(n27305) );
  NAND3X1 U16048 ( .A(n27308), .B(n27309), .C(n27310), .Y(n27307) );
  NOR2X1 U16049 ( .A(n27311), .B(n27312), .Y(n27310) );
  OAI22X1 U16050 ( .A(n25155), .B(n27313), .C(n25166), .D(n27314), .Y(n27312)
         );
  OAI22X1 U16051 ( .A(n25176), .B(n27315), .C(n25187), .D(n27316), .Y(n27311)
         );
  AOI22X1 U16052 ( .A(reg_file[1482]), .B(n25198), .C(reg_file[1354]), .D(
        n25208), .Y(n27309) );
  AOI22X1 U16053 ( .A(reg_file[1226]), .B(n25219), .C(reg_file[1098]), .D(
        n25229), .Y(n27308) );
  NAND3X1 U16054 ( .A(n27317), .B(n27318), .C(n27319), .Y(n27306) );
  NOR2X1 U16055 ( .A(n27320), .B(n27321), .Y(n27319) );
  OAI22X1 U16056 ( .A(n25239), .B(n27322), .C(n25250), .D(n27323), .Y(n27321)
         );
  OAI22X1 U16057 ( .A(n25260), .B(n27324), .C(n25271), .D(n27325), .Y(n27320)
         );
  AOI22X1 U16058 ( .A(reg_file[586]), .B(n25282), .C(reg_file[714]), .D(n25292), .Y(n27318) );
  AOI22X1 U16059 ( .A(reg_file[842]), .B(n25303), .C(reg_file[970]), .D(n25313), .Y(n27317) );
  NOR2X1 U16060 ( .A(n27326), .B(n27327), .Y(n27304) );
  NAND3X1 U16061 ( .A(n27328), .B(n27329), .C(n27330), .Y(n27327) );
  NOR2X1 U16062 ( .A(n27331), .B(n27332), .Y(n27330) );
  OAI22X1 U16063 ( .A(n25323), .B(n27333), .C(n25334), .D(n27334), .Y(n27332)
         );
  OAI22X1 U16064 ( .A(n25344), .B(n27335), .C(n25355), .D(n27336), .Y(n27331)
         );
  AOI22X1 U16065 ( .A(reg_file[3530]), .B(n25366), .C(reg_file[3402]), .D(
        n25376), .Y(n27329) );
  AOI22X1 U16066 ( .A(reg_file[3274]), .B(n25387), .C(reg_file[3146]), .D(
        n25397), .Y(n27328) );
  NAND3X1 U16067 ( .A(n27337), .B(n27338), .C(n27339), .Y(n27326) );
  NOR2X1 U16068 ( .A(n27340), .B(n27341), .Y(n27339) );
  OAI22X1 U16069 ( .A(n25407), .B(n27342), .C(n25418), .D(n27343), .Y(n27341)
         );
  OAI22X1 U16070 ( .A(n25428), .B(n27344), .C(n25439), .D(n27345), .Y(n27340)
         );
  AOI22X1 U16071 ( .A(reg_file[2506]), .B(n25450), .C(reg_file[2378]), .D(
        n25460), .Y(n27338) );
  AOI22X1 U16072 ( .A(reg_file[2250]), .B(n25471), .C(reg_file[2122]), .D(
        n25481), .Y(n27337) );
  AOI21X1 U16073 ( .A(n27346), .B(n27347), .C(n25145), .Y(rd2data1040_73_) );
  NOR2X1 U16074 ( .A(n27348), .B(n27349), .Y(n27347) );
  NAND3X1 U16075 ( .A(n27350), .B(n27351), .C(n27352), .Y(n27349) );
  NOR2X1 U16076 ( .A(n27353), .B(n27354), .Y(n27352) );
  OAI22X1 U16077 ( .A(n25155), .B(n27355), .C(n25166), .D(n27356), .Y(n27354)
         );
  OAI22X1 U16078 ( .A(n25176), .B(n27357), .C(n25187), .D(n27358), .Y(n27353)
         );
  AOI22X1 U16079 ( .A(reg_file[1481]), .B(n25198), .C(reg_file[1353]), .D(
        n25208), .Y(n27351) );
  AOI22X1 U16080 ( .A(reg_file[1225]), .B(n25219), .C(reg_file[1097]), .D(
        n25229), .Y(n27350) );
  NAND3X1 U16081 ( .A(n27359), .B(n27360), .C(n27361), .Y(n27348) );
  NOR2X1 U16082 ( .A(n27362), .B(n27363), .Y(n27361) );
  OAI22X1 U16083 ( .A(n25239), .B(n27364), .C(n25250), .D(n27365), .Y(n27363)
         );
  OAI22X1 U16084 ( .A(n25260), .B(n27366), .C(n25271), .D(n27367), .Y(n27362)
         );
  AOI22X1 U16085 ( .A(reg_file[585]), .B(n25282), .C(reg_file[713]), .D(n25292), .Y(n27360) );
  AOI22X1 U16086 ( .A(reg_file[841]), .B(n25303), .C(reg_file[969]), .D(n25313), .Y(n27359) );
  NOR2X1 U16087 ( .A(n27368), .B(n27369), .Y(n27346) );
  NAND3X1 U16088 ( .A(n27370), .B(n27371), .C(n27372), .Y(n27369) );
  NOR2X1 U16089 ( .A(n27373), .B(n27374), .Y(n27372) );
  OAI22X1 U16090 ( .A(n25323), .B(n27375), .C(n25334), .D(n27376), .Y(n27374)
         );
  OAI22X1 U16091 ( .A(n25344), .B(n27377), .C(n25355), .D(n27378), .Y(n27373)
         );
  AOI22X1 U16092 ( .A(reg_file[3529]), .B(n25366), .C(reg_file[3401]), .D(
        n25376), .Y(n27371) );
  AOI22X1 U16093 ( .A(reg_file[3273]), .B(n25387), .C(reg_file[3145]), .D(
        n25397), .Y(n27370) );
  NAND3X1 U16094 ( .A(n27379), .B(n27380), .C(n27381), .Y(n27368) );
  NOR2X1 U16095 ( .A(n27382), .B(n27383), .Y(n27381) );
  OAI22X1 U16096 ( .A(n25407), .B(n27384), .C(n25418), .D(n27385), .Y(n27383)
         );
  OAI22X1 U16097 ( .A(n25428), .B(n27386), .C(n25439), .D(n27387), .Y(n27382)
         );
  AOI22X1 U16098 ( .A(reg_file[2505]), .B(n25450), .C(reg_file[2377]), .D(
        n25460), .Y(n27380) );
  AOI22X1 U16099 ( .A(reg_file[2249]), .B(n25471), .C(reg_file[2121]), .D(
        n25481), .Y(n27379) );
  AOI21X1 U16100 ( .A(n27388), .B(n27389), .C(n25145), .Y(rd2data1040_72_) );
  NOR2X1 U16101 ( .A(n27390), .B(n27391), .Y(n27389) );
  NAND3X1 U16102 ( .A(n27392), .B(n27393), .C(n27394), .Y(n27391) );
  NOR2X1 U16103 ( .A(n27395), .B(n27396), .Y(n27394) );
  OAI22X1 U16104 ( .A(n25155), .B(n27397), .C(n25166), .D(n27398), .Y(n27396)
         );
  OAI22X1 U16105 ( .A(n25176), .B(n27399), .C(n25187), .D(n27400), .Y(n27395)
         );
  AOI22X1 U16106 ( .A(reg_file[1480]), .B(n25198), .C(reg_file[1352]), .D(
        n25208), .Y(n27393) );
  AOI22X1 U16107 ( .A(reg_file[1224]), .B(n25219), .C(reg_file[1096]), .D(
        n25229), .Y(n27392) );
  NAND3X1 U16108 ( .A(n27401), .B(n27402), .C(n27403), .Y(n27390) );
  NOR2X1 U16109 ( .A(n27404), .B(n27405), .Y(n27403) );
  OAI22X1 U16110 ( .A(n25239), .B(n27406), .C(n25250), .D(n27407), .Y(n27405)
         );
  OAI22X1 U16111 ( .A(n25260), .B(n27408), .C(n25271), .D(n27409), .Y(n27404)
         );
  AOI22X1 U16112 ( .A(reg_file[584]), .B(n25282), .C(reg_file[712]), .D(n25292), .Y(n27402) );
  AOI22X1 U16113 ( .A(reg_file[840]), .B(n25303), .C(reg_file[968]), .D(n25313), .Y(n27401) );
  NOR2X1 U16114 ( .A(n27410), .B(n27411), .Y(n27388) );
  NAND3X1 U16115 ( .A(n27412), .B(n27413), .C(n27414), .Y(n27411) );
  NOR2X1 U16116 ( .A(n27415), .B(n27416), .Y(n27414) );
  OAI22X1 U16117 ( .A(n25323), .B(n27417), .C(n25334), .D(n27418), .Y(n27416)
         );
  OAI22X1 U16118 ( .A(n25344), .B(n27419), .C(n25355), .D(n27420), .Y(n27415)
         );
  AOI22X1 U16119 ( .A(reg_file[3528]), .B(n25366), .C(reg_file[3400]), .D(
        n25376), .Y(n27413) );
  AOI22X1 U16120 ( .A(reg_file[3272]), .B(n25387), .C(reg_file[3144]), .D(
        n25397), .Y(n27412) );
  NAND3X1 U16121 ( .A(n27421), .B(n27422), .C(n27423), .Y(n27410) );
  NOR2X1 U16122 ( .A(n27424), .B(n27425), .Y(n27423) );
  OAI22X1 U16123 ( .A(n25407), .B(n27426), .C(n25418), .D(n27427), .Y(n27425)
         );
  OAI22X1 U16124 ( .A(n25428), .B(n27428), .C(n25439), .D(n27429), .Y(n27424)
         );
  AOI22X1 U16125 ( .A(reg_file[2504]), .B(n25450), .C(reg_file[2376]), .D(
        n25460), .Y(n27422) );
  AOI22X1 U16126 ( .A(reg_file[2248]), .B(n25471), .C(reg_file[2120]), .D(
        n25481), .Y(n27421) );
  AOI21X1 U16127 ( .A(n27430), .B(n27431), .C(n25145), .Y(rd2data1040_71_) );
  NOR2X1 U16128 ( .A(n27432), .B(n27433), .Y(n27431) );
  NAND3X1 U16129 ( .A(n27434), .B(n27435), .C(n27436), .Y(n27433) );
  NOR2X1 U16130 ( .A(n27437), .B(n27438), .Y(n27436) );
  OAI22X1 U16131 ( .A(n25155), .B(n27439), .C(n25166), .D(n27440), .Y(n27438)
         );
  OAI22X1 U16132 ( .A(n25176), .B(n27441), .C(n25187), .D(n27442), .Y(n27437)
         );
  AOI22X1 U16133 ( .A(reg_file[1479]), .B(n25198), .C(reg_file[1351]), .D(
        n25208), .Y(n27435) );
  AOI22X1 U16134 ( .A(reg_file[1223]), .B(n25219), .C(reg_file[1095]), .D(
        n25229), .Y(n27434) );
  NAND3X1 U16135 ( .A(n27443), .B(n27444), .C(n27445), .Y(n27432) );
  NOR2X1 U16136 ( .A(n27446), .B(n27447), .Y(n27445) );
  OAI22X1 U16137 ( .A(n25239), .B(n27448), .C(n25250), .D(n27449), .Y(n27447)
         );
  OAI22X1 U16138 ( .A(n25260), .B(n27450), .C(n25271), .D(n27451), .Y(n27446)
         );
  AOI22X1 U16139 ( .A(reg_file[583]), .B(n25282), .C(reg_file[711]), .D(n25292), .Y(n27444) );
  AOI22X1 U16140 ( .A(reg_file[839]), .B(n25303), .C(reg_file[967]), .D(n25313), .Y(n27443) );
  NOR2X1 U16141 ( .A(n27452), .B(n27453), .Y(n27430) );
  NAND3X1 U16142 ( .A(n27454), .B(n27455), .C(n27456), .Y(n27453) );
  NOR2X1 U16143 ( .A(n27457), .B(n27458), .Y(n27456) );
  OAI22X1 U16144 ( .A(n25323), .B(n27459), .C(n25334), .D(n27460), .Y(n27458)
         );
  OAI22X1 U16145 ( .A(n25344), .B(n27461), .C(n25355), .D(n27462), .Y(n27457)
         );
  AOI22X1 U16146 ( .A(reg_file[3527]), .B(n25366), .C(reg_file[3399]), .D(
        n25376), .Y(n27455) );
  AOI22X1 U16147 ( .A(reg_file[3271]), .B(n25387), .C(reg_file[3143]), .D(
        n25397), .Y(n27454) );
  NAND3X1 U16148 ( .A(n27463), .B(n27464), .C(n27465), .Y(n27452) );
  NOR2X1 U16149 ( .A(n27466), .B(n27467), .Y(n27465) );
  OAI22X1 U16150 ( .A(n25407), .B(n27468), .C(n25418), .D(n27469), .Y(n27467)
         );
  OAI22X1 U16151 ( .A(n25428), .B(n27470), .C(n25439), .D(n27471), .Y(n27466)
         );
  AOI22X1 U16152 ( .A(reg_file[2503]), .B(n25450), .C(reg_file[2375]), .D(
        n25460), .Y(n27464) );
  AOI22X1 U16153 ( .A(reg_file[2247]), .B(n25471), .C(reg_file[2119]), .D(
        n25481), .Y(n27463) );
  AOI21X1 U16154 ( .A(n27472), .B(n27473), .C(n25144), .Y(rd2data1040_70_) );
  NOR2X1 U16155 ( .A(n27474), .B(n27475), .Y(n27473) );
  NAND3X1 U16156 ( .A(n27476), .B(n27477), .C(n27478), .Y(n27475) );
  NOR2X1 U16157 ( .A(n27479), .B(n27480), .Y(n27478) );
  OAI22X1 U16158 ( .A(n25155), .B(n27481), .C(n25165), .D(n27482), .Y(n27480)
         );
  OAI22X1 U16159 ( .A(n25176), .B(n27483), .C(n25186), .D(n27484), .Y(n27479)
         );
  AOI22X1 U16160 ( .A(reg_file[1478]), .B(n25197), .C(reg_file[1350]), .D(
        n25208), .Y(n27477) );
  AOI22X1 U16161 ( .A(reg_file[1222]), .B(n25218), .C(reg_file[1094]), .D(
        n25229), .Y(n27476) );
  NAND3X1 U16162 ( .A(n27485), .B(n27486), .C(n27487), .Y(n27474) );
  NOR2X1 U16163 ( .A(n27488), .B(n27489), .Y(n27487) );
  OAI22X1 U16164 ( .A(n25239), .B(n27490), .C(n25249), .D(n27491), .Y(n27489)
         );
  OAI22X1 U16165 ( .A(n25260), .B(n27492), .C(n25270), .D(n27493), .Y(n27488)
         );
  AOI22X1 U16166 ( .A(reg_file[582]), .B(n25281), .C(reg_file[710]), .D(n25292), .Y(n27486) );
  AOI22X1 U16167 ( .A(reg_file[838]), .B(n25302), .C(reg_file[966]), .D(n25313), .Y(n27485) );
  NOR2X1 U16168 ( .A(n27494), .B(n27495), .Y(n27472) );
  NAND3X1 U16169 ( .A(n27496), .B(n27497), .C(n27498), .Y(n27495) );
  NOR2X1 U16170 ( .A(n27499), .B(n27500), .Y(n27498) );
  OAI22X1 U16171 ( .A(n25323), .B(n27501), .C(n25333), .D(n27502), .Y(n27500)
         );
  OAI22X1 U16172 ( .A(n25344), .B(n27503), .C(n25354), .D(n27504), .Y(n27499)
         );
  AOI22X1 U16173 ( .A(reg_file[3526]), .B(n25365), .C(reg_file[3398]), .D(
        n25376), .Y(n27497) );
  AOI22X1 U16174 ( .A(reg_file[3270]), .B(n25386), .C(reg_file[3142]), .D(
        n25397), .Y(n27496) );
  NAND3X1 U16175 ( .A(n27505), .B(n27506), .C(n27507), .Y(n27494) );
  NOR2X1 U16176 ( .A(n27508), .B(n27509), .Y(n27507) );
  OAI22X1 U16177 ( .A(n25407), .B(n27510), .C(n25417), .D(n27511), .Y(n27509)
         );
  OAI22X1 U16178 ( .A(n25428), .B(n27512), .C(n25438), .D(n27513), .Y(n27508)
         );
  AOI22X1 U16179 ( .A(reg_file[2502]), .B(n25449), .C(reg_file[2374]), .D(
        n25460), .Y(n27506) );
  AOI22X1 U16180 ( .A(reg_file[2246]), .B(n25470), .C(reg_file[2118]), .D(
        n25481), .Y(n27505) );
  AOI21X1 U16181 ( .A(n27514), .B(n27515), .C(n25144), .Y(rd2data1040_6_) );
  NOR2X1 U16182 ( .A(n27516), .B(n27517), .Y(n27515) );
  NAND3X1 U16183 ( .A(n27518), .B(n27519), .C(n27520), .Y(n27517) );
  NOR2X1 U16184 ( .A(n27521), .B(n27522), .Y(n27520) );
  OAI22X1 U16185 ( .A(n25155), .B(n27523), .C(n25165), .D(n27524), .Y(n27522)
         );
  OAI22X1 U16186 ( .A(n25176), .B(n27525), .C(n25186), .D(n27526), .Y(n27521)
         );
  AOI22X1 U16187 ( .A(reg_file[1414]), .B(n25197), .C(reg_file[1286]), .D(
        n25208), .Y(n27519) );
  AOI22X1 U16188 ( .A(reg_file[1158]), .B(n25218), .C(reg_file[1030]), .D(
        n25229), .Y(n27518) );
  NAND3X1 U16189 ( .A(n27527), .B(n27528), .C(n27529), .Y(n27516) );
  NOR2X1 U16190 ( .A(n27530), .B(n27531), .Y(n27529) );
  OAI22X1 U16191 ( .A(n25239), .B(n27532), .C(n25249), .D(n27533), .Y(n27531)
         );
  OAI22X1 U16192 ( .A(n25260), .B(n27534), .C(n25270), .D(n27535), .Y(n27530)
         );
  AOI22X1 U16193 ( .A(reg_file[518]), .B(n25281), .C(reg_file[646]), .D(n25292), .Y(n27528) );
  AOI22X1 U16194 ( .A(reg_file[774]), .B(n25302), .C(reg_file[902]), .D(n25313), .Y(n27527) );
  NOR2X1 U16195 ( .A(n27536), .B(n27537), .Y(n27514) );
  NAND3X1 U16196 ( .A(n27538), .B(n27539), .C(n27540), .Y(n27537) );
  NOR2X1 U16197 ( .A(n27541), .B(n27542), .Y(n27540) );
  OAI22X1 U16198 ( .A(n25323), .B(n27543), .C(n25333), .D(n27544), .Y(n27542)
         );
  OAI22X1 U16199 ( .A(n25344), .B(n27545), .C(n25354), .D(n27546), .Y(n27541)
         );
  AOI22X1 U16200 ( .A(reg_file[3462]), .B(n25365), .C(reg_file[3334]), .D(
        n25376), .Y(n27539) );
  AOI22X1 U16201 ( .A(reg_file[3206]), .B(n25386), .C(reg_file[3078]), .D(
        n25397), .Y(n27538) );
  NAND3X1 U16202 ( .A(n27547), .B(n27548), .C(n27549), .Y(n27536) );
  NOR2X1 U16203 ( .A(n27550), .B(n27551), .Y(n27549) );
  OAI22X1 U16204 ( .A(n25407), .B(n27552), .C(n25417), .D(n27553), .Y(n27551)
         );
  OAI22X1 U16205 ( .A(n25428), .B(n27554), .C(n25438), .D(n27555), .Y(n27550)
         );
  AOI22X1 U16206 ( .A(reg_file[2438]), .B(n25449), .C(reg_file[2310]), .D(
        n25460), .Y(n27548) );
  AOI22X1 U16207 ( .A(reg_file[2182]), .B(n25470), .C(reg_file[2054]), .D(
        n25481), .Y(n27547) );
  AOI21X1 U16208 ( .A(n27556), .B(n27557), .C(n25144), .Y(rd2data1040_69_) );
  NOR2X1 U16209 ( .A(n27558), .B(n27559), .Y(n27557) );
  NAND3X1 U16210 ( .A(n27560), .B(n27561), .C(n27562), .Y(n27559) );
  NOR2X1 U16211 ( .A(n27563), .B(n27564), .Y(n27562) );
  OAI22X1 U16212 ( .A(n25155), .B(n27565), .C(n25165), .D(n27566), .Y(n27564)
         );
  OAI22X1 U16213 ( .A(n25176), .B(n27567), .C(n25186), .D(n27568), .Y(n27563)
         );
  AOI22X1 U16214 ( .A(reg_file[1477]), .B(n25197), .C(reg_file[1349]), .D(
        n25208), .Y(n27561) );
  AOI22X1 U16215 ( .A(reg_file[1221]), .B(n25218), .C(reg_file[1093]), .D(
        n25229), .Y(n27560) );
  NAND3X1 U16216 ( .A(n27569), .B(n27570), .C(n27571), .Y(n27558) );
  NOR2X1 U16217 ( .A(n27572), .B(n27573), .Y(n27571) );
  OAI22X1 U16218 ( .A(n25239), .B(n27574), .C(n25249), .D(n27575), .Y(n27573)
         );
  OAI22X1 U16219 ( .A(n25260), .B(n27576), .C(n25270), .D(n27577), .Y(n27572)
         );
  AOI22X1 U16220 ( .A(reg_file[581]), .B(n25281), .C(reg_file[709]), .D(n25292), .Y(n27570) );
  AOI22X1 U16221 ( .A(reg_file[837]), .B(n25302), .C(reg_file[965]), .D(n25313), .Y(n27569) );
  NOR2X1 U16222 ( .A(n27578), .B(n27579), .Y(n27556) );
  NAND3X1 U16223 ( .A(n27580), .B(n27581), .C(n27582), .Y(n27579) );
  NOR2X1 U16224 ( .A(n27583), .B(n27584), .Y(n27582) );
  OAI22X1 U16225 ( .A(n25323), .B(n27585), .C(n25333), .D(n27586), .Y(n27584)
         );
  OAI22X1 U16226 ( .A(n25344), .B(n27587), .C(n25354), .D(n27588), .Y(n27583)
         );
  AOI22X1 U16227 ( .A(reg_file[3525]), .B(n25365), .C(reg_file[3397]), .D(
        n25376), .Y(n27581) );
  AOI22X1 U16228 ( .A(reg_file[3269]), .B(n25386), .C(reg_file[3141]), .D(
        n25397), .Y(n27580) );
  NAND3X1 U16229 ( .A(n27589), .B(n27590), .C(n27591), .Y(n27578) );
  NOR2X1 U16230 ( .A(n27592), .B(n27593), .Y(n27591) );
  OAI22X1 U16231 ( .A(n25407), .B(n27594), .C(n25417), .D(n27595), .Y(n27593)
         );
  OAI22X1 U16232 ( .A(n25428), .B(n27596), .C(n25438), .D(n27597), .Y(n27592)
         );
  AOI22X1 U16233 ( .A(reg_file[2501]), .B(n25449), .C(reg_file[2373]), .D(
        n25460), .Y(n27590) );
  AOI22X1 U16234 ( .A(reg_file[2245]), .B(n25470), .C(reg_file[2117]), .D(
        n25481), .Y(n27589) );
  AOI21X1 U16235 ( .A(n27598), .B(n27599), .C(n25144), .Y(rd2data1040_68_) );
  NOR2X1 U16236 ( .A(n27600), .B(n27601), .Y(n27599) );
  NAND3X1 U16237 ( .A(n27602), .B(n27603), .C(n27604), .Y(n27601) );
  NOR2X1 U16238 ( .A(n27605), .B(n27606), .Y(n27604) );
  OAI22X1 U16239 ( .A(n25155), .B(n27607), .C(n25165), .D(n27608), .Y(n27606)
         );
  OAI22X1 U16240 ( .A(n25176), .B(n27609), .C(n25186), .D(n27610), .Y(n27605)
         );
  AOI22X1 U16241 ( .A(reg_file[1476]), .B(n25197), .C(reg_file[1348]), .D(
        n25208), .Y(n27603) );
  AOI22X1 U16242 ( .A(reg_file[1220]), .B(n25218), .C(reg_file[1092]), .D(
        n25229), .Y(n27602) );
  NAND3X1 U16243 ( .A(n27611), .B(n27612), .C(n27613), .Y(n27600) );
  NOR2X1 U16244 ( .A(n27614), .B(n27615), .Y(n27613) );
  OAI22X1 U16245 ( .A(n25239), .B(n27616), .C(n25249), .D(n27617), .Y(n27615)
         );
  OAI22X1 U16246 ( .A(n25260), .B(n27618), .C(n25270), .D(n27619), .Y(n27614)
         );
  AOI22X1 U16247 ( .A(reg_file[580]), .B(n25281), .C(reg_file[708]), .D(n25292), .Y(n27612) );
  AOI22X1 U16248 ( .A(reg_file[836]), .B(n25302), .C(reg_file[964]), .D(n25313), .Y(n27611) );
  NOR2X1 U16249 ( .A(n27620), .B(n27621), .Y(n27598) );
  NAND3X1 U16250 ( .A(n27622), .B(n27623), .C(n27624), .Y(n27621) );
  NOR2X1 U16251 ( .A(n27625), .B(n27626), .Y(n27624) );
  OAI22X1 U16252 ( .A(n25323), .B(n27627), .C(n25333), .D(n27628), .Y(n27626)
         );
  OAI22X1 U16253 ( .A(n25344), .B(n27629), .C(n25354), .D(n27630), .Y(n27625)
         );
  AOI22X1 U16254 ( .A(reg_file[3524]), .B(n25365), .C(reg_file[3396]), .D(
        n25376), .Y(n27623) );
  AOI22X1 U16255 ( .A(reg_file[3268]), .B(n25386), .C(reg_file[3140]), .D(
        n25397), .Y(n27622) );
  NAND3X1 U16256 ( .A(n27631), .B(n27632), .C(n27633), .Y(n27620) );
  NOR2X1 U16257 ( .A(n27634), .B(n27635), .Y(n27633) );
  OAI22X1 U16258 ( .A(n25407), .B(n27636), .C(n25417), .D(n27637), .Y(n27635)
         );
  OAI22X1 U16259 ( .A(n25428), .B(n27638), .C(n25438), .D(n27639), .Y(n27634)
         );
  AOI22X1 U16260 ( .A(reg_file[2500]), .B(n25449), .C(reg_file[2372]), .D(
        n25460), .Y(n27632) );
  AOI22X1 U16261 ( .A(reg_file[2244]), .B(n25470), .C(reg_file[2116]), .D(
        n25481), .Y(n27631) );
  AOI21X1 U16262 ( .A(n27640), .B(n27641), .C(n25144), .Y(rd2data1040_67_) );
  NOR2X1 U16263 ( .A(n27642), .B(n27643), .Y(n27641) );
  NAND3X1 U16264 ( .A(n27644), .B(n27645), .C(n27646), .Y(n27643) );
  NOR2X1 U16265 ( .A(n27647), .B(n27648), .Y(n27646) );
  OAI22X1 U16266 ( .A(n25155), .B(n27649), .C(n25165), .D(n27650), .Y(n27648)
         );
  OAI22X1 U16267 ( .A(n25176), .B(n27651), .C(n25186), .D(n27652), .Y(n27647)
         );
  AOI22X1 U16268 ( .A(reg_file[1475]), .B(n25197), .C(reg_file[1347]), .D(
        n25208), .Y(n27645) );
  AOI22X1 U16269 ( .A(reg_file[1219]), .B(n25218), .C(reg_file[1091]), .D(
        n25229), .Y(n27644) );
  NAND3X1 U16270 ( .A(n27653), .B(n27654), .C(n27655), .Y(n27642) );
  NOR2X1 U16271 ( .A(n27656), .B(n27657), .Y(n27655) );
  OAI22X1 U16272 ( .A(n25239), .B(n27658), .C(n25249), .D(n27659), .Y(n27657)
         );
  OAI22X1 U16273 ( .A(n25260), .B(n27660), .C(n25270), .D(n27661), .Y(n27656)
         );
  AOI22X1 U16274 ( .A(reg_file[579]), .B(n25281), .C(reg_file[707]), .D(n25292), .Y(n27654) );
  AOI22X1 U16275 ( .A(reg_file[835]), .B(n25302), .C(reg_file[963]), .D(n25313), .Y(n27653) );
  NOR2X1 U16276 ( .A(n27662), .B(n27663), .Y(n27640) );
  NAND3X1 U16277 ( .A(n27664), .B(n27665), .C(n27666), .Y(n27663) );
  NOR2X1 U16278 ( .A(n27667), .B(n27668), .Y(n27666) );
  OAI22X1 U16279 ( .A(n25323), .B(n27669), .C(n25333), .D(n27670), .Y(n27668)
         );
  OAI22X1 U16280 ( .A(n25344), .B(n27671), .C(n25354), .D(n27672), .Y(n27667)
         );
  AOI22X1 U16281 ( .A(reg_file[3523]), .B(n25365), .C(reg_file[3395]), .D(
        n25376), .Y(n27665) );
  AOI22X1 U16282 ( .A(reg_file[3267]), .B(n25386), .C(reg_file[3139]), .D(
        n25397), .Y(n27664) );
  NAND3X1 U16283 ( .A(n27673), .B(n27674), .C(n27675), .Y(n27662) );
  NOR2X1 U16284 ( .A(n27676), .B(n27677), .Y(n27675) );
  OAI22X1 U16285 ( .A(n25407), .B(n27678), .C(n25417), .D(n27679), .Y(n27677)
         );
  OAI22X1 U16286 ( .A(n25428), .B(n27680), .C(n25438), .D(n27681), .Y(n27676)
         );
  AOI22X1 U16287 ( .A(reg_file[2499]), .B(n25449), .C(reg_file[2371]), .D(
        n25460), .Y(n27674) );
  AOI22X1 U16288 ( .A(reg_file[2243]), .B(n25470), .C(reg_file[2115]), .D(
        n25481), .Y(n27673) );
  AOI21X1 U16289 ( .A(n27682), .B(n27683), .C(n25144), .Y(rd2data1040_66_) );
  NOR2X1 U16290 ( .A(n27684), .B(n27685), .Y(n27683) );
  NAND3X1 U16291 ( .A(n27686), .B(n27687), .C(n27688), .Y(n27685) );
  NOR2X1 U16292 ( .A(n27689), .B(n27690), .Y(n27688) );
  OAI22X1 U16293 ( .A(n25154), .B(n27691), .C(n25165), .D(n27692), .Y(n27690)
         );
  OAI22X1 U16294 ( .A(n25175), .B(n27693), .C(n25186), .D(n27694), .Y(n27689)
         );
  AOI22X1 U16295 ( .A(reg_file[1474]), .B(n25197), .C(reg_file[1346]), .D(
        n25207), .Y(n27687) );
  AOI22X1 U16296 ( .A(reg_file[1218]), .B(n25218), .C(reg_file[1090]), .D(
        n25228), .Y(n27686) );
  NAND3X1 U16297 ( .A(n27695), .B(n27696), .C(n27697), .Y(n27684) );
  NOR2X1 U16298 ( .A(n27698), .B(n27699), .Y(n27697) );
  OAI22X1 U16299 ( .A(n25238), .B(n27700), .C(n25249), .D(n27701), .Y(n27699)
         );
  OAI22X1 U16300 ( .A(n25259), .B(n27702), .C(n25270), .D(n27703), .Y(n27698)
         );
  AOI22X1 U16301 ( .A(reg_file[578]), .B(n25281), .C(reg_file[706]), .D(n25291), .Y(n27696) );
  AOI22X1 U16302 ( .A(reg_file[834]), .B(n25302), .C(reg_file[962]), .D(n25312), .Y(n27695) );
  NOR2X1 U16303 ( .A(n27704), .B(n27705), .Y(n27682) );
  NAND3X1 U16304 ( .A(n27706), .B(n27707), .C(n27708), .Y(n27705) );
  NOR2X1 U16305 ( .A(n27709), .B(n27710), .Y(n27708) );
  OAI22X1 U16306 ( .A(n25322), .B(n27711), .C(n25333), .D(n27712), .Y(n27710)
         );
  OAI22X1 U16307 ( .A(n25343), .B(n27713), .C(n25354), .D(n27714), .Y(n27709)
         );
  AOI22X1 U16308 ( .A(reg_file[3522]), .B(n25365), .C(reg_file[3394]), .D(
        n25375), .Y(n27707) );
  AOI22X1 U16309 ( .A(reg_file[3266]), .B(n25386), .C(reg_file[3138]), .D(
        n25396), .Y(n27706) );
  NAND3X1 U16310 ( .A(n27715), .B(n27716), .C(n27717), .Y(n27704) );
  NOR2X1 U16311 ( .A(n27718), .B(n27719), .Y(n27717) );
  OAI22X1 U16312 ( .A(n25406), .B(n27720), .C(n25417), .D(n27721), .Y(n27719)
         );
  OAI22X1 U16313 ( .A(n25427), .B(n27722), .C(n25438), .D(n27723), .Y(n27718)
         );
  AOI22X1 U16314 ( .A(reg_file[2498]), .B(n25449), .C(reg_file[2370]), .D(
        n25459), .Y(n27716) );
  AOI22X1 U16315 ( .A(reg_file[2242]), .B(n25470), .C(reg_file[2114]), .D(
        n25480), .Y(n27715) );
  AOI21X1 U16316 ( .A(n27724), .B(n27725), .C(n25144), .Y(rd2data1040_65_) );
  NOR2X1 U16317 ( .A(n27726), .B(n27727), .Y(n27725) );
  NAND3X1 U16318 ( .A(n27728), .B(n27729), .C(n27730), .Y(n27727) );
  NOR2X1 U16319 ( .A(n27731), .B(n27732), .Y(n27730) );
  OAI22X1 U16320 ( .A(n25154), .B(n27733), .C(n25165), .D(n27734), .Y(n27732)
         );
  OAI22X1 U16321 ( .A(n25175), .B(n27735), .C(n25186), .D(n27736), .Y(n27731)
         );
  AOI22X1 U16322 ( .A(reg_file[1473]), .B(n25197), .C(reg_file[1345]), .D(
        n25207), .Y(n27729) );
  AOI22X1 U16323 ( .A(reg_file[1217]), .B(n25218), .C(reg_file[1089]), .D(
        n25228), .Y(n27728) );
  NAND3X1 U16324 ( .A(n27737), .B(n27738), .C(n27739), .Y(n27726) );
  NOR2X1 U16325 ( .A(n27740), .B(n27741), .Y(n27739) );
  OAI22X1 U16326 ( .A(n25238), .B(n27742), .C(n25249), .D(n27743), .Y(n27741)
         );
  OAI22X1 U16327 ( .A(n25259), .B(n27744), .C(n25270), .D(n27745), .Y(n27740)
         );
  AOI22X1 U16328 ( .A(reg_file[577]), .B(n25281), .C(reg_file[705]), .D(n25291), .Y(n27738) );
  AOI22X1 U16329 ( .A(reg_file[833]), .B(n25302), .C(reg_file[961]), .D(n25312), .Y(n27737) );
  NOR2X1 U16330 ( .A(n27746), .B(n27747), .Y(n27724) );
  NAND3X1 U16331 ( .A(n27748), .B(n27749), .C(n27750), .Y(n27747) );
  NOR2X1 U16332 ( .A(n27751), .B(n27752), .Y(n27750) );
  OAI22X1 U16333 ( .A(n25322), .B(n27753), .C(n25333), .D(n27754), .Y(n27752)
         );
  OAI22X1 U16334 ( .A(n25343), .B(n27755), .C(n25354), .D(n27756), .Y(n27751)
         );
  AOI22X1 U16335 ( .A(reg_file[3521]), .B(n25365), .C(reg_file[3393]), .D(
        n25375), .Y(n27749) );
  AOI22X1 U16336 ( .A(reg_file[3265]), .B(n25386), .C(reg_file[3137]), .D(
        n25396), .Y(n27748) );
  NAND3X1 U16337 ( .A(n27757), .B(n27758), .C(n27759), .Y(n27746) );
  NOR2X1 U16338 ( .A(n27760), .B(n27761), .Y(n27759) );
  OAI22X1 U16339 ( .A(n25406), .B(n27762), .C(n25417), .D(n27763), .Y(n27761)
         );
  OAI22X1 U16340 ( .A(n25427), .B(n27764), .C(n25438), .D(n27765), .Y(n27760)
         );
  AOI22X1 U16341 ( .A(reg_file[2497]), .B(n25449), .C(reg_file[2369]), .D(
        n25459), .Y(n27758) );
  AOI22X1 U16342 ( .A(reg_file[2241]), .B(n25470), .C(reg_file[2113]), .D(
        n25480), .Y(n27757) );
  AOI21X1 U16343 ( .A(n27766), .B(n27767), .C(n25144), .Y(rd2data1040_64_) );
  NOR2X1 U16344 ( .A(n27768), .B(n27769), .Y(n27767) );
  NAND3X1 U16345 ( .A(n27770), .B(n27771), .C(n27772), .Y(n27769) );
  NOR2X1 U16346 ( .A(n27773), .B(n27774), .Y(n27772) );
  OAI22X1 U16347 ( .A(n25154), .B(n27775), .C(n25165), .D(n27776), .Y(n27774)
         );
  OAI22X1 U16348 ( .A(n25175), .B(n27777), .C(n25186), .D(n27778), .Y(n27773)
         );
  AOI22X1 U16349 ( .A(reg_file[1472]), .B(n25197), .C(reg_file[1344]), .D(
        n25207), .Y(n27771) );
  AOI22X1 U16350 ( .A(reg_file[1216]), .B(n25218), .C(reg_file[1088]), .D(
        n25228), .Y(n27770) );
  NAND3X1 U16351 ( .A(n27779), .B(n27780), .C(n27781), .Y(n27768) );
  NOR2X1 U16352 ( .A(n27782), .B(n27783), .Y(n27781) );
  OAI22X1 U16353 ( .A(n25238), .B(n27784), .C(n25249), .D(n27785), .Y(n27783)
         );
  OAI22X1 U16354 ( .A(n25259), .B(n27786), .C(n25270), .D(n27787), .Y(n27782)
         );
  AOI22X1 U16355 ( .A(reg_file[576]), .B(n25281), .C(reg_file[704]), .D(n25291), .Y(n27780) );
  AOI22X1 U16356 ( .A(reg_file[832]), .B(n25302), .C(reg_file[960]), .D(n25312), .Y(n27779) );
  NOR2X1 U16357 ( .A(n27788), .B(n27789), .Y(n27766) );
  NAND3X1 U16358 ( .A(n27790), .B(n27791), .C(n27792), .Y(n27789) );
  NOR2X1 U16359 ( .A(n27793), .B(n27794), .Y(n27792) );
  OAI22X1 U16360 ( .A(n25322), .B(n27795), .C(n25333), .D(n27796), .Y(n27794)
         );
  OAI22X1 U16361 ( .A(n25343), .B(n27797), .C(n25354), .D(n27798), .Y(n27793)
         );
  AOI22X1 U16362 ( .A(reg_file[3520]), .B(n25365), .C(reg_file[3392]), .D(
        n25375), .Y(n27791) );
  AOI22X1 U16363 ( .A(reg_file[3264]), .B(n25386), .C(reg_file[3136]), .D(
        n25396), .Y(n27790) );
  NAND3X1 U16364 ( .A(n27799), .B(n27800), .C(n27801), .Y(n27788) );
  NOR2X1 U16365 ( .A(n27802), .B(n27803), .Y(n27801) );
  OAI22X1 U16366 ( .A(n25406), .B(n27804), .C(n25417), .D(n27805), .Y(n27803)
         );
  OAI22X1 U16367 ( .A(n25427), .B(n27806), .C(n25438), .D(n27807), .Y(n27802)
         );
  AOI22X1 U16368 ( .A(reg_file[2496]), .B(n25449), .C(reg_file[2368]), .D(
        n25459), .Y(n27800) );
  AOI22X1 U16369 ( .A(reg_file[2240]), .B(n25470), .C(reg_file[2112]), .D(
        n25480), .Y(n27799) );
  AOI21X1 U16370 ( .A(n27808), .B(n27809), .C(n25144), .Y(rd2data1040_63_) );
  NOR2X1 U16371 ( .A(n27810), .B(n27811), .Y(n27809) );
  NAND3X1 U16372 ( .A(n27812), .B(n27813), .C(n27814), .Y(n27811) );
  NOR2X1 U16373 ( .A(n27815), .B(n27816), .Y(n27814) );
  OAI22X1 U16374 ( .A(n25154), .B(n27817), .C(n25165), .D(n27818), .Y(n27816)
         );
  OAI22X1 U16375 ( .A(n25175), .B(n27819), .C(n25186), .D(n27820), .Y(n27815)
         );
  AOI22X1 U16376 ( .A(reg_file[1471]), .B(n25197), .C(reg_file[1343]), .D(
        n25207), .Y(n27813) );
  AOI22X1 U16377 ( .A(reg_file[1215]), .B(n25218), .C(reg_file[1087]), .D(
        n25228), .Y(n27812) );
  NAND3X1 U16378 ( .A(n27821), .B(n27822), .C(n27823), .Y(n27810) );
  NOR2X1 U16379 ( .A(n27824), .B(n27825), .Y(n27823) );
  OAI22X1 U16380 ( .A(n25238), .B(n27826), .C(n25249), .D(n27827), .Y(n27825)
         );
  OAI22X1 U16381 ( .A(n25259), .B(n27828), .C(n25270), .D(n27829), .Y(n27824)
         );
  AOI22X1 U16382 ( .A(reg_file[575]), .B(n25281), .C(reg_file[703]), .D(n25291), .Y(n27822) );
  AOI22X1 U16383 ( .A(reg_file[831]), .B(n25302), .C(reg_file[959]), .D(n25312), .Y(n27821) );
  NOR2X1 U16384 ( .A(n27830), .B(n27831), .Y(n27808) );
  NAND3X1 U16385 ( .A(n27832), .B(n27833), .C(n27834), .Y(n27831) );
  NOR2X1 U16386 ( .A(n27835), .B(n27836), .Y(n27834) );
  OAI22X1 U16387 ( .A(n25322), .B(n27837), .C(n25333), .D(n27838), .Y(n27836)
         );
  OAI22X1 U16388 ( .A(n25343), .B(n27839), .C(n25354), .D(n27840), .Y(n27835)
         );
  AOI22X1 U16389 ( .A(reg_file[3519]), .B(n25365), .C(reg_file[3391]), .D(
        n25375), .Y(n27833) );
  AOI22X1 U16390 ( .A(reg_file[3263]), .B(n25386), .C(reg_file[3135]), .D(
        n25396), .Y(n27832) );
  NAND3X1 U16391 ( .A(n27841), .B(n27842), .C(n27843), .Y(n27830) );
  NOR2X1 U16392 ( .A(n27844), .B(n27845), .Y(n27843) );
  OAI22X1 U16393 ( .A(n25406), .B(n27846), .C(n25417), .D(n27847), .Y(n27845)
         );
  OAI22X1 U16394 ( .A(n25427), .B(n27848), .C(n25438), .D(n27849), .Y(n27844)
         );
  AOI22X1 U16395 ( .A(reg_file[2495]), .B(n25449), .C(reg_file[2367]), .D(
        n25459), .Y(n27842) );
  AOI22X1 U16396 ( .A(reg_file[2239]), .B(n25470), .C(reg_file[2111]), .D(
        n25480), .Y(n27841) );
  AOI21X1 U16397 ( .A(n27850), .B(n27851), .C(n25144), .Y(rd2data1040_62_) );
  NOR2X1 U16398 ( .A(n27852), .B(n27853), .Y(n27851) );
  NAND3X1 U16399 ( .A(n27854), .B(n27855), .C(n27856), .Y(n27853) );
  NOR2X1 U16400 ( .A(n27857), .B(n27858), .Y(n27856) );
  OAI22X1 U16401 ( .A(n25154), .B(n27859), .C(n25165), .D(n27860), .Y(n27858)
         );
  OAI22X1 U16402 ( .A(n25175), .B(n27861), .C(n25186), .D(n27862), .Y(n27857)
         );
  AOI22X1 U16403 ( .A(reg_file[1470]), .B(n25197), .C(reg_file[1342]), .D(
        n25207), .Y(n27855) );
  AOI22X1 U16404 ( .A(reg_file[1214]), .B(n25218), .C(reg_file[1086]), .D(
        n25228), .Y(n27854) );
  NAND3X1 U16405 ( .A(n27863), .B(n27864), .C(n27865), .Y(n27852) );
  NOR2X1 U16406 ( .A(n27866), .B(n27867), .Y(n27865) );
  OAI22X1 U16407 ( .A(n25238), .B(n27868), .C(n25249), .D(n27869), .Y(n27867)
         );
  OAI22X1 U16408 ( .A(n25259), .B(n27870), .C(n25270), .D(n27871), .Y(n27866)
         );
  AOI22X1 U16409 ( .A(reg_file[574]), .B(n25281), .C(reg_file[702]), .D(n25291), .Y(n27864) );
  AOI22X1 U16410 ( .A(reg_file[830]), .B(n25302), .C(reg_file[958]), .D(n25312), .Y(n27863) );
  NOR2X1 U16411 ( .A(n27872), .B(n27873), .Y(n27850) );
  NAND3X1 U16412 ( .A(n27874), .B(n27875), .C(n27876), .Y(n27873) );
  NOR2X1 U16413 ( .A(n27877), .B(n27878), .Y(n27876) );
  OAI22X1 U16414 ( .A(n25322), .B(n27879), .C(n25333), .D(n27880), .Y(n27878)
         );
  OAI22X1 U16415 ( .A(n25343), .B(n27881), .C(n25354), .D(n27882), .Y(n27877)
         );
  AOI22X1 U16416 ( .A(reg_file[3518]), .B(n25365), .C(reg_file[3390]), .D(
        n25375), .Y(n27875) );
  AOI22X1 U16417 ( .A(reg_file[3262]), .B(n25386), .C(reg_file[3134]), .D(
        n25396), .Y(n27874) );
  NAND3X1 U16418 ( .A(n27883), .B(n27884), .C(n27885), .Y(n27872) );
  NOR2X1 U16419 ( .A(n27886), .B(n27887), .Y(n27885) );
  OAI22X1 U16420 ( .A(n25406), .B(n27888), .C(n25417), .D(n27889), .Y(n27887)
         );
  OAI22X1 U16421 ( .A(n25427), .B(n27890), .C(n25438), .D(n27891), .Y(n27886)
         );
  AOI22X1 U16422 ( .A(reg_file[2494]), .B(n25449), .C(reg_file[2366]), .D(
        n25459), .Y(n27884) );
  AOI22X1 U16423 ( .A(reg_file[2238]), .B(n25470), .C(reg_file[2110]), .D(
        n25480), .Y(n27883) );
  AOI21X1 U16424 ( .A(n27892), .B(n27893), .C(n25144), .Y(rd2data1040_61_) );
  NOR2X1 U16425 ( .A(n27894), .B(n27895), .Y(n27893) );
  NAND3X1 U16426 ( .A(n27896), .B(n27897), .C(n27898), .Y(n27895) );
  NOR2X1 U16427 ( .A(n27899), .B(n27900), .Y(n27898) );
  OAI22X1 U16428 ( .A(n25154), .B(n27901), .C(n25165), .D(n27902), .Y(n27900)
         );
  OAI22X1 U16429 ( .A(n25175), .B(n27903), .C(n25186), .D(n27904), .Y(n27899)
         );
  AOI22X1 U16430 ( .A(reg_file[1469]), .B(n25197), .C(reg_file[1341]), .D(
        n25207), .Y(n27897) );
  AOI22X1 U16431 ( .A(reg_file[1213]), .B(n25218), .C(reg_file[1085]), .D(
        n25228), .Y(n27896) );
  NAND3X1 U16432 ( .A(n27905), .B(n27906), .C(n27907), .Y(n27894) );
  NOR2X1 U16433 ( .A(n27908), .B(n27909), .Y(n27907) );
  OAI22X1 U16434 ( .A(n25238), .B(n27910), .C(n25249), .D(n27911), .Y(n27909)
         );
  OAI22X1 U16435 ( .A(n25259), .B(n27912), .C(n25270), .D(n27913), .Y(n27908)
         );
  AOI22X1 U16436 ( .A(reg_file[573]), .B(n25281), .C(reg_file[701]), .D(n25291), .Y(n27906) );
  AOI22X1 U16437 ( .A(reg_file[829]), .B(n25302), .C(reg_file[957]), .D(n25312), .Y(n27905) );
  NOR2X1 U16438 ( .A(n27914), .B(n27915), .Y(n27892) );
  NAND3X1 U16439 ( .A(n27916), .B(n27917), .C(n27918), .Y(n27915) );
  NOR2X1 U16440 ( .A(n27919), .B(n27920), .Y(n27918) );
  OAI22X1 U16441 ( .A(n25322), .B(n27921), .C(n25333), .D(n27922), .Y(n27920)
         );
  OAI22X1 U16442 ( .A(n25343), .B(n27923), .C(n25354), .D(n27924), .Y(n27919)
         );
  AOI22X1 U16443 ( .A(reg_file[3517]), .B(n25365), .C(reg_file[3389]), .D(
        n25375), .Y(n27917) );
  AOI22X1 U16444 ( .A(reg_file[3261]), .B(n25386), .C(reg_file[3133]), .D(
        n25396), .Y(n27916) );
  NAND3X1 U16445 ( .A(n27925), .B(n27926), .C(n27927), .Y(n27914) );
  NOR2X1 U16446 ( .A(n27928), .B(n27929), .Y(n27927) );
  OAI22X1 U16447 ( .A(n25406), .B(n27930), .C(n25417), .D(n27931), .Y(n27929)
         );
  OAI22X1 U16448 ( .A(n25427), .B(n27932), .C(n25438), .D(n27933), .Y(n27928)
         );
  AOI22X1 U16449 ( .A(reg_file[2493]), .B(n25449), .C(reg_file[2365]), .D(
        n25459), .Y(n27926) );
  AOI22X1 U16450 ( .A(reg_file[2237]), .B(n25470), .C(reg_file[2109]), .D(
        n25480), .Y(n27925) );
  AOI21X1 U16451 ( .A(n27934), .B(n27935), .C(n25144), .Y(rd2data1040_60_) );
  NOR2X1 U16452 ( .A(n27936), .B(n27937), .Y(n27935) );
  NAND3X1 U16453 ( .A(n27938), .B(n27939), .C(n27940), .Y(n27937) );
  NOR2X1 U16454 ( .A(n27941), .B(n27942), .Y(n27940) );
  OAI22X1 U16455 ( .A(n25154), .B(n27943), .C(n25165), .D(n27944), .Y(n27942)
         );
  OAI22X1 U16456 ( .A(n25175), .B(n27945), .C(n25186), .D(n27946), .Y(n27941)
         );
  AOI22X1 U16457 ( .A(reg_file[1468]), .B(n25197), .C(reg_file[1340]), .D(
        n25207), .Y(n27939) );
  AOI22X1 U16458 ( .A(reg_file[1212]), .B(n25218), .C(reg_file[1084]), .D(
        n25228), .Y(n27938) );
  NAND3X1 U16459 ( .A(n27947), .B(n27948), .C(n27949), .Y(n27936) );
  NOR2X1 U16460 ( .A(n27950), .B(n27951), .Y(n27949) );
  OAI22X1 U16461 ( .A(n25238), .B(n27952), .C(n25249), .D(n27953), .Y(n27951)
         );
  OAI22X1 U16462 ( .A(n25259), .B(n27954), .C(n25270), .D(n27955), .Y(n27950)
         );
  AOI22X1 U16463 ( .A(reg_file[572]), .B(n25281), .C(reg_file[700]), .D(n25291), .Y(n27948) );
  AOI22X1 U16464 ( .A(reg_file[828]), .B(n25302), .C(reg_file[956]), .D(n25312), .Y(n27947) );
  NOR2X1 U16465 ( .A(n27956), .B(n27957), .Y(n27934) );
  NAND3X1 U16466 ( .A(n27958), .B(n27959), .C(n27960), .Y(n27957) );
  NOR2X1 U16467 ( .A(n27961), .B(n27962), .Y(n27960) );
  OAI22X1 U16468 ( .A(n25322), .B(n27963), .C(n25333), .D(n27964), .Y(n27962)
         );
  OAI22X1 U16469 ( .A(n25343), .B(n27965), .C(n25354), .D(n27966), .Y(n27961)
         );
  AOI22X1 U16470 ( .A(reg_file[3516]), .B(n25365), .C(reg_file[3388]), .D(
        n25375), .Y(n27959) );
  AOI22X1 U16471 ( .A(reg_file[3260]), .B(n25386), .C(reg_file[3132]), .D(
        n25396), .Y(n27958) );
  NAND3X1 U16472 ( .A(n27967), .B(n27968), .C(n27969), .Y(n27956) );
  NOR2X1 U16473 ( .A(n27970), .B(n27971), .Y(n27969) );
  OAI22X1 U16474 ( .A(n25406), .B(n27972), .C(n25417), .D(n27973), .Y(n27971)
         );
  OAI22X1 U16475 ( .A(n25427), .B(n27974), .C(n25438), .D(n27975), .Y(n27970)
         );
  AOI22X1 U16476 ( .A(reg_file[2492]), .B(n25449), .C(reg_file[2364]), .D(
        n25459), .Y(n27968) );
  AOI22X1 U16477 ( .A(reg_file[2236]), .B(n25470), .C(reg_file[2108]), .D(
        n25480), .Y(n27967) );
  AOI21X1 U16478 ( .A(n27976), .B(n27977), .C(n25143), .Y(rd2data1040_5_) );
  NOR2X1 U16479 ( .A(n27978), .B(n27979), .Y(n27977) );
  NAND3X1 U16480 ( .A(n27980), .B(n27981), .C(n27982), .Y(n27979) );
  NOR2X1 U16481 ( .A(n27983), .B(n27984), .Y(n27982) );
  OAI22X1 U16482 ( .A(n25154), .B(n27985), .C(n25164), .D(n27986), .Y(n27984)
         );
  OAI22X1 U16483 ( .A(n25175), .B(n27987), .C(n25185), .D(n27988), .Y(n27983)
         );
  AOI22X1 U16484 ( .A(reg_file[1413]), .B(n25196), .C(reg_file[1285]), .D(
        n25207), .Y(n27981) );
  AOI22X1 U16485 ( .A(reg_file[1157]), .B(n25217), .C(reg_file[1029]), .D(
        n25228), .Y(n27980) );
  NAND3X1 U16486 ( .A(n27989), .B(n27990), .C(n27991), .Y(n27978) );
  NOR2X1 U16487 ( .A(n27992), .B(n27993), .Y(n27991) );
  OAI22X1 U16488 ( .A(n25238), .B(n27994), .C(n25248), .D(n27995), .Y(n27993)
         );
  OAI22X1 U16489 ( .A(n25259), .B(n27996), .C(n25269), .D(n27997), .Y(n27992)
         );
  AOI22X1 U16490 ( .A(reg_file[517]), .B(n25280), .C(reg_file[645]), .D(n25291), .Y(n27990) );
  AOI22X1 U16491 ( .A(reg_file[773]), .B(n25301), .C(reg_file[901]), .D(n25312), .Y(n27989) );
  NOR2X1 U16492 ( .A(n27998), .B(n27999), .Y(n27976) );
  NAND3X1 U16493 ( .A(n28000), .B(n28001), .C(n28002), .Y(n27999) );
  NOR2X1 U16494 ( .A(n28003), .B(n28004), .Y(n28002) );
  OAI22X1 U16495 ( .A(n25322), .B(n28005), .C(n25332), .D(n28006), .Y(n28004)
         );
  OAI22X1 U16496 ( .A(n25343), .B(n28007), .C(n25353), .D(n28008), .Y(n28003)
         );
  AOI22X1 U16497 ( .A(reg_file[3461]), .B(n25364), .C(reg_file[3333]), .D(
        n25375), .Y(n28001) );
  AOI22X1 U16498 ( .A(reg_file[3205]), .B(n25385), .C(reg_file[3077]), .D(
        n25396), .Y(n28000) );
  NAND3X1 U16499 ( .A(n28009), .B(n28010), .C(n28011), .Y(n27998) );
  NOR2X1 U16500 ( .A(n28012), .B(n28013), .Y(n28011) );
  OAI22X1 U16501 ( .A(n25406), .B(n28014), .C(n25416), .D(n28015), .Y(n28013)
         );
  OAI22X1 U16502 ( .A(n25427), .B(n28016), .C(n25437), .D(n28017), .Y(n28012)
         );
  AOI22X1 U16503 ( .A(reg_file[2437]), .B(n25448), .C(reg_file[2309]), .D(
        n25459), .Y(n28010) );
  AOI22X1 U16504 ( .A(reg_file[2181]), .B(n25469), .C(reg_file[2053]), .D(
        n25480), .Y(n28009) );
  AOI21X1 U16505 ( .A(n28018), .B(n28019), .C(n25143), .Y(rd2data1040_59_) );
  NOR2X1 U16506 ( .A(n28020), .B(n28021), .Y(n28019) );
  NAND3X1 U16507 ( .A(n28022), .B(n28023), .C(n28024), .Y(n28021) );
  NOR2X1 U16508 ( .A(n28025), .B(n28026), .Y(n28024) );
  OAI22X1 U16509 ( .A(n25154), .B(n28027), .C(n25164), .D(n28028), .Y(n28026)
         );
  OAI22X1 U16510 ( .A(n25175), .B(n28029), .C(n25185), .D(n28030), .Y(n28025)
         );
  AOI22X1 U16511 ( .A(reg_file[1467]), .B(n25196), .C(reg_file[1339]), .D(
        n25207), .Y(n28023) );
  AOI22X1 U16512 ( .A(reg_file[1211]), .B(n25217), .C(reg_file[1083]), .D(
        n25228), .Y(n28022) );
  NAND3X1 U16513 ( .A(n28031), .B(n28032), .C(n28033), .Y(n28020) );
  NOR2X1 U16514 ( .A(n28034), .B(n28035), .Y(n28033) );
  OAI22X1 U16515 ( .A(n25238), .B(n28036), .C(n25248), .D(n28037), .Y(n28035)
         );
  OAI22X1 U16516 ( .A(n25259), .B(n28038), .C(n25269), .D(n28039), .Y(n28034)
         );
  AOI22X1 U16517 ( .A(reg_file[571]), .B(n25280), .C(reg_file[699]), .D(n25291), .Y(n28032) );
  AOI22X1 U16518 ( .A(reg_file[827]), .B(n25301), .C(reg_file[955]), .D(n25312), .Y(n28031) );
  NOR2X1 U16519 ( .A(n28040), .B(n28041), .Y(n28018) );
  NAND3X1 U16520 ( .A(n28042), .B(n28043), .C(n28044), .Y(n28041) );
  NOR2X1 U16521 ( .A(n28045), .B(n28046), .Y(n28044) );
  OAI22X1 U16522 ( .A(n25322), .B(n28047), .C(n25332), .D(n28048), .Y(n28046)
         );
  OAI22X1 U16523 ( .A(n25343), .B(n28049), .C(n25353), .D(n28050), .Y(n28045)
         );
  AOI22X1 U16524 ( .A(reg_file[3515]), .B(n25364), .C(reg_file[3387]), .D(
        n25375), .Y(n28043) );
  AOI22X1 U16525 ( .A(reg_file[3259]), .B(n25385), .C(reg_file[3131]), .D(
        n25396), .Y(n28042) );
  NAND3X1 U16526 ( .A(n28051), .B(n28052), .C(n28053), .Y(n28040) );
  NOR2X1 U16527 ( .A(n28054), .B(n28055), .Y(n28053) );
  OAI22X1 U16528 ( .A(n25406), .B(n28056), .C(n25416), .D(n28057), .Y(n28055)
         );
  OAI22X1 U16529 ( .A(n25427), .B(n28058), .C(n25437), .D(n28059), .Y(n28054)
         );
  AOI22X1 U16530 ( .A(reg_file[2491]), .B(n25448), .C(reg_file[2363]), .D(
        n25459), .Y(n28052) );
  AOI22X1 U16531 ( .A(reg_file[2235]), .B(n25469), .C(reg_file[2107]), .D(
        n25480), .Y(n28051) );
  AOI21X1 U16532 ( .A(n28060), .B(n28061), .C(n25143), .Y(rd2data1040_58_) );
  NOR2X1 U16533 ( .A(n28062), .B(n28063), .Y(n28061) );
  NAND3X1 U16534 ( .A(n28064), .B(n28065), .C(n28066), .Y(n28063) );
  NOR2X1 U16535 ( .A(n28067), .B(n28068), .Y(n28066) );
  OAI22X1 U16536 ( .A(n25154), .B(n28069), .C(n25164), .D(n28070), .Y(n28068)
         );
  OAI22X1 U16537 ( .A(n25175), .B(n28071), .C(n25185), .D(n28072), .Y(n28067)
         );
  AOI22X1 U16538 ( .A(reg_file[1466]), .B(n25196), .C(reg_file[1338]), .D(
        n25207), .Y(n28065) );
  AOI22X1 U16539 ( .A(reg_file[1210]), .B(n25217), .C(reg_file[1082]), .D(
        n25228), .Y(n28064) );
  NAND3X1 U16540 ( .A(n28073), .B(n28074), .C(n28075), .Y(n28062) );
  NOR2X1 U16541 ( .A(n28076), .B(n28077), .Y(n28075) );
  OAI22X1 U16542 ( .A(n25238), .B(n28078), .C(n25248), .D(n28079), .Y(n28077)
         );
  OAI22X1 U16543 ( .A(n25259), .B(n28080), .C(n25269), .D(n28081), .Y(n28076)
         );
  AOI22X1 U16544 ( .A(reg_file[570]), .B(n25280), .C(reg_file[698]), .D(n25291), .Y(n28074) );
  AOI22X1 U16545 ( .A(reg_file[826]), .B(n25301), .C(reg_file[954]), .D(n25312), .Y(n28073) );
  NOR2X1 U16546 ( .A(n28082), .B(n28083), .Y(n28060) );
  NAND3X1 U16547 ( .A(n28084), .B(n28085), .C(n28086), .Y(n28083) );
  NOR2X1 U16548 ( .A(n28087), .B(n28088), .Y(n28086) );
  OAI22X1 U16549 ( .A(n25322), .B(n28089), .C(n25332), .D(n28090), .Y(n28088)
         );
  OAI22X1 U16550 ( .A(n25343), .B(n28091), .C(n25353), .D(n28092), .Y(n28087)
         );
  AOI22X1 U16551 ( .A(reg_file[3514]), .B(n25364), .C(reg_file[3386]), .D(
        n25375), .Y(n28085) );
  AOI22X1 U16552 ( .A(reg_file[3258]), .B(n25385), .C(reg_file[3130]), .D(
        n25396), .Y(n28084) );
  NAND3X1 U16553 ( .A(n28093), .B(n28094), .C(n28095), .Y(n28082) );
  NOR2X1 U16554 ( .A(n28096), .B(n28097), .Y(n28095) );
  OAI22X1 U16555 ( .A(n25406), .B(n28098), .C(n25416), .D(n28099), .Y(n28097)
         );
  OAI22X1 U16556 ( .A(n25427), .B(n28100), .C(n25437), .D(n28101), .Y(n28096)
         );
  AOI22X1 U16557 ( .A(reg_file[2490]), .B(n25448), .C(reg_file[2362]), .D(
        n25459), .Y(n28094) );
  AOI22X1 U16558 ( .A(reg_file[2234]), .B(n25469), .C(reg_file[2106]), .D(
        n25480), .Y(n28093) );
  AOI21X1 U16559 ( .A(n28102), .B(n28103), .C(n25143), .Y(rd2data1040_57_) );
  NOR2X1 U16560 ( .A(n28104), .B(n28105), .Y(n28103) );
  NAND3X1 U16561 ( .A(n28106), .B(n28107), .C(n28108), .Y(n28105) );
  NOR2X1 U16562 ( .A(n28109), .B(n28110), .Y(n28108) );
  OAI22X1 U16563 ( .A(n25154), .B(n28111), .C(n25164), .D(n28112), .Y(n28110)
         );
  OAI22X1 U16564 ( .A(n25175), .B(n28113), .C(n25185), .D(n28114), .Y(n28109)
         );
  AOI22X1 U16565 ( .A(reg_file[1465]), .B(n25196), .C(reg_file[1337]), .D(
        n25207), .Y(n28107) );
  AOI22X1 U16566 ( .A(reg_file[1209]), .B(n25217), .C(reg_file[1081]), .D(
        n25228), .Y(n28106) );
  NAND3X1 U16567 ( .A(n28115), .B(n28116), .C(n28117), .Y(n28104) );
  NOR2X1 U16568 ( .A(n28118), .B(n28119), .Y(n28117) );
  OAI22X1 U16569 ( .A(n25238), .B(n28120), .C(n25248), .D(n28121), .Y(n28119)
         );
  OAI22X1 U16570 ( .A(n25259), .B(n28122), .C(n25269), .D(n28123), .Y(n28118)
         );
  AOI22X1 U16571 ( .A(reg_file[569]), .B(n25280), .C(reg_file[697]), .D(n25291), .Y(n28116) );
  AOI22X1 U16572 ( .A(reg_file[825]), .B(n25301), .C(reg_file[953]), .D(n25312), .Y(n28115) );
  NOR2X1 U16573 ( .A(n28124), .B(n28125), .Y(n28102) );
  NAND3X1 U16574 ( .A(n28126), .B(n28127), .C(n28128), .Y(n28125) );
  NOR2X1 U16575 ( .A(n28129), .B(n28130), .Y(n28128) );
  OAI22X1 U16576 ( .A(n25322), .B(n28131), .C(n25332), .D(n28132), .Y(n28130)
         );
  OAI22X1 U16577 ( .A(n25343), .B(n28133), .C(n25353), .D(n28134), .Y(n28129)
         );
  AOI22X1 U16578 ( .A(reg_file[3513]), .B(n25364), .C(reg_file[3385]), .D(
        n25375), .Y(n28127) );
  AOI22X1 U16579 ( .A(reg_file[3257]), .B(n25385), .C(reg_file[3129]), .D(
        n25396), .Y(n28126) );
  NAND3X1 U16580 ( .A(n28135), .B(n28136), .C(n28137), .Y(n28124) );
  NOR2X1 U16581 ( .A(n28138), .B(n28139), .Y(n28137) );
  OAI22X1 U16582 ( .A(n25406), .B(n28140), .C(n25416), .D(n28141), .Y(n28139)
         );
  OAI22X1 U16583 ( .A(n25427), .B(n28142), .C(n25437), .D(n28143), .Y(n28138)
         );
  AOI22X1 U16584 ( .A(reg_file[2489]), .B(n25448), .C(reg_file[2361]), .D(
        n25459), .Y(n28136) );
  AOI22X1 U16585 ( .A(reg_file[2233]), .B(n25469), .C(reg_file[2105]), .D(
        n25480), .Y(n28135) );
  AOI21X1 U16586 ( .A(n28144), .B(n28145), .C(n25143), .Y(rd2data1040_56_) );
  NOR2X1 U16587 ( .A(n28146), .B(n28147), .Y(n28145) );
  NAND3X1 U16588 ( .A(n28148), .B(n28149), .C(n28150), .Y(n28147) );
  NOR2X1 U16589 ( .A(n28151), .B(n28152), .Y(n28150) );
  OAI22X1 U16590 ( .A(n25154), .B(n28153), .C(n25164), .D(n28154), .Y(n28152)
         );
  OAI22X1 U16591 ( .A(n25175), .B(n28155), .C(n25185), .D(n28156), .Y(n28151)
         );
  AOI22X1 U16592 ( .A(reg_file[1464]), .B(n25196), .C(reg_file[1336]), .D(
        n25207), .Y(n28149) );
  AOI22X1 U16593 ( .A(reg_file[1208]), .B(n25217), .C(reg_file[1080]), .D(
        n25228), .Y(n28148) );
  NAND3X1 U16594 ( .A(n28157), .B(n28158), .C(n28159), .Y(n28146) );
  NOR2X1 U16595 ( .A(n28160), .B(n28161), .Y(n28159) );
  OAI22X1 U16596 ( .A(n25238), .B(n28162), .C(n25248), .D(n28163), .Y(n28161)
         );
  OAI22X1 U16597 ( .A(n25259), .B(n28164), .C(n25269), .D(n28165), .Y(n28160)
         );
  AOI22X1 U16598 ( .A(reg_file[568]), .B(n25280), .C(reg_file[696]), .D(n25291), .Y(n28158) );
  AOI22X1 U16599 ( .A(reg_file[824]), .B(n25301), .C(reg_file[952]), .D(n25312), .Y(n28157) );
  NOR2X1 U16600 ( .A(n28166), .B(n28167), .Y(n28144) );
  NAND3X1 U16601 ( .A(n28168), .B(n28169), .C(n28170), .Y(n28167) );
  NOR2X1 U16602 ( .A(n28171), .B(n28172), .Y(n28170) );
  OAI22X1 U16603 ( .A(n25322), .B(n28173), .C(n25332), .D(n28174), .Y(n28172)
         );
  OAI22X1 U16604 ( .A(n25343), .B(n28175), .C(n25353), .D(n28176), .Y(n28171)
         );
  AOI22X1 U16605 ( .A(reg_file[3512]), .B(n25364), .C(reg_file[3384]), .D(
        n25375), .Y(n28169) );
  AOI22X1 U16606 ( .A(reg_file[3256]), .B(n25385), .C(reg_file[3128]), .D(
        n25396), .Y(n28168) );
  NAND3X1 U16607 ( .A(n28177), .B(n28178), .C(n28179), .Y(n28166) );
  NOR2X1 U16608 ( .A(n28180), .B(n28181), .Y(n28179) );
  OAI22X1 U16609 ( .A(n25406), .B(n28182), .C(n25416), .D(n28183), .Y(n28181)
         );
  OAI22X1 U16610 ( .A(n25427), .B(n28184), .C(n25437), .D(n28185), .Y(n28180)
         );
  AOI22X1 U16611 ( .A(reg_file[2488]), .B(n25448), .C(reg_file[2360]), .D(
        n25459), .Y(n28178) );
  AOI22X1 U16612 ( .A(reg_file[2232]), .B(n25469), .C(reg_file[2104]), .D(
        n25480), .Y(n28177) );
  AOI21X1 U16613 ( .A(n28186), .B(n28187), .C(n25143), .Y(rd2data1040_55_) );
  NOR2X1 U16614 ( .A(n28188), .B(n28189), .Y(n28187) );
  NAND3X1 U16615 ( .A(n28190), .B(n28191), .C(n28192), .Y(n28189) );
  NOR2X1 U16616 ( .A(n28193), .B(n28194), .Y(n28192) );
  OAI22X1 U16617 ( .A(n25154), .B(n28195), .C(n25164), .D(n28196), .Y(n28194)
         );
  OAI22X1 U16618 ( .A(n25175), .B(n28197), .C(n25185), .D(n28198), .Y(n28193)
         );
  AOI22X1 U16619 ( .A(reg_file[1463]), .B(n25196), .C(reg_file[1335]), .D(
        n25207), .Y(n28191) );
  AOI22X1 U16620 ( .A(reg_file[1207]), .B(n25217), .C(reg_file[1079]), .D(
        n25228), .Y(n28190) );
  NAND3X1 U16621 ( .A(n28199), .B(n28200), .C(n28201), .Y(n28188) );
  NOR2X1 U16622 ( .A(n28202), .B(n28203), .Y(n28201) );
  OAI22X1 U16623 ( .A(n25238), .B(n28204), .C(n25248), .D(n28205), .Y(n28203)
         );
  OAI22X1 U16624 ( .A(n25259), .B(n28206), .C(n25269), .D(n28207), .Y(n28202)
         );
  AOI22X1 U16625 ( .A(reg_file[567]), .B(n25280), .C(reg_file[695]), .D(n25291), .Y(n28200) );
  AOI22X1 U16626 ( .A(reg_file[823]), .B(n25301), .C(reg_file[951]), .D(n25312), .Y(n28199) );
  NOR2X1 U16627 ( .A(n28208), .B(n28209), .Y(n28186) );
  NAND3X1 U16628 ( .A(n28210), .B(n28211), .C(n28212), .Y(n28209) );
  NOR2X1 U16629 ( .A(n28213), .B(n28214), .Y(n28212) );
  OAI22X1 U16630 ( .A(n25322), .B(n28215), .C(n25332), .D(n28216), .Y(n28214)
         );
  OAI22X1 U16631 ( .A(n25343), .B(n28217), .C(n25353), .D(n28218), .Y(n28213)
         );
  AOI22X1 U16632 ( .A(reg_file[3511]), .B(n25364), .C(reg_file[3383]), .D(
        n25375), .Y(n28211) );
  AOI22X1 U16633 ( .A(reg_file[3255]), .B(n25385), .C(reg_file[3127]), .D(
        n25396), .Y(n28210) );
  NAND3X1 U16634 ( .A(n28219), .B(n28220), .C(n28221), .Y(n28208) );
  NOR2X1 U16635 ( .A(n28222), .B(n28223), .Y(n28221) );
  OAI22X1 U16636 ( .A(n25406), .B(n28224), .C(n25416), .D(n28225), .Y(n28223)
         );
  OAI22X1 U16637 ( .A(n25427), .B(n28226), .C(n25437), .D(n28227), .Y(n28222)
         );
  AOI22X1 U16638 ( .A(reg_file[2487]), .B(n25448), .C(reg_file[2359]), .D(
        n25459), .Y(n28220) );
  AOI22X1 U16639 ( .A(reg_file[2231]), .B(n25469), .C(reg_file[2103]), .D(
        n25480), .Y(n28219) );
  AOI21X1 U16640 ( .A(n28228), .B(n28229), .C(n25143), .Y(rd2data1040_54_) );
  NOR2X1 U16641 ( .A(n28230), .B(n28231), .Y(n28229) );
  NAND3X1 U16642 ( .A(n28232), .B(n28233), .C(n28234), .Y(n28231) );
  NOR2X1 U16643 ( .A(n28235), .B(n28236), .Y(n28234) );
  OAI22X1 U16644 ( .A(n25153), .B(n28237), .C(n25164), .D(n28238), .Y(n28236)
         );
  OAI22X1 U16645 ( .A(n25174), .B(n28239), .C(n25185), .D(n28240), .Y(n28235)
         );
  AOI22X1 U16646 ( .A(reg_file[1462]), .B(n25196), .C(reg_file[1334]), .D(
        n25206), .Y(n28233) );
  AOI22X1 U16647 ( .A(reg_file[1206]), .B(n25217), .C(reg_file[1078]), .D(
        n25227), .Y(n28232) );
  NAND3X1 U16648 ( .A(n28241), .B(n28242), .C(n28243), .Y(n28230) );
  NOR2X1 U16649 ( .A(n28244), .B(n28245), .Y(n28243) );
  OAI22X1 U16650 ( .A(n25237), .B(n28246), .C(n25248), .D(n28247), .Y(n28245)
         );
  OAI22X1 U16651 ( .A(n25258), .B(n28248), .C(n25269), .D(n28249), .Y(n28244)
         );
  AOI22X1 U16652 ( .A(reg_file[566]), .B(n25280), .C(reg_file[694]), .D(n25290), .Y(n28242) );
  AOI22X1 U16653 ( .A(reg_file[822]), .B(n25301), .C(reg_file[950]), .D(n25311), .Y(n28241) );
  NOR2X1 U16654 ( .A(n28250), .B(n28251), .Y(n28228) );
  NAND3X1 U16655 ( .A(n28252), .B(n28253), .C(n28254), .Y(n28251) );
  NOR2X1 U16656 ( .A(n28255), .B(n28256), .Y(n28254) );
  OAI22X1 U16657 ( .A(n25321), .B(n28257), .C(n25332), .D(n28258), .Y(n28256)
         );
  OAI22X1 U16658 ( .A(n25342), .B(n28259), .C(n25353), .D(n28260), .Y(n28255)
         );
  AOI22X1 U16659 ( .A(reg_file[3510]), .B(n25364), .C(reg_file[3382]), .D(
        n25374), .Y(n28253) );
  AOI22X1 U16660 ( .A(reg_file[3254]), .B(n25385), .C(reg_file[3126]), .D(
        n25395), .Y(n28252) );
  NAND3X1 U16661 ( .A(n28261), .B(n28262), .C(n28263), .Y(n28250) );
  NOR2X1 U16662 ( .A(n28264), .B(n28265), .Y(n28263) );
  OAI22X1 U16663 ( .A(n25405), .B(n28266), .C(n25416), .D(n28267), .Y(n28265)
         );
  OAI22X1 U16664 ( .A(n25426), .B(n28268), .C(n25437), .D(n28269), .Y(n28264)
         );
  AOI22X1 U16665 ( .A(reg_file[2486]), .B(n25448), .C(reg_file[2358]), .D(
        n25458), .Y(n28262) );
  AOI22X1 U16666 ( .A(reg_file[2230]), .B(n25469), .C(reg_file[2102]), .D(
        n25479), .Y(n28261) );
  AOI21X1 U16667 ( .A(n28270), .B(n28271), .C(n25143), .Y(rd2data1040_53_) );
  NOR2X1 U16668 ( .A(n28272), .B(n28273), .Y(n28271) );
  NAND3X1 U16669 ( .A(n28274), .B(n28275), .C(n28276), .Y(n28273) );
  NOR2X1 U16670 ( .A(n28277), .B(n28278), .Y(n28276) );
  OAI22X1 U16671 ( .A(n25153), .B(n28279), .C(n25164), .D(n28280), .Y(n28278)
         );
  OAI22X1 U16672 ( .A(n25174), .B(n28281), .C(n25185), .D(n28282), .Y(n28277)
         );
  AOI22X1 U16673 ( .A(reg_file[1461]), .B(n25196), .C(reg_file[1333]), .D(
        n25206), .Y(n28275) );
  AOI22X1 U16674 ( .A(reg_file[1205]), .B(n25217), .C(reg_file[1077]), .D(
        n25227), .Y(n28274) );
  NAND3X1 U16675 ( .A(n28283), .B(n28284), .C(n28285), .Y(n28272) );
  NOR2X1 U16676 ( .A(n28286), .B(n28287), .Y(n28285) );
  OAI22X1 U16677 ( .A(n25237), .B(n28288), .C(n25248), .D(n28289), .Y(n28287)
         );
  OAI22X1 U16678 ( .A(n25258), .B(n28290), .C(n25269), .D(n28291), .Y(n28286)
         );
  AOI22X1 U16679 ( .A(reg_file[565]), .B(n25280), .C(reg_file[693]), .D(n25290), .Y(n28284) );
  AOI22X1 U16680 ( .A(reg_file[821]), .B(n25301), .C(reg_file[949]), .D(n25311), .Y(n28283) );
  NOR2X1 U16681 ( .A(n28292), .B(n28293), .Y(n28270) );
  NAND3X1 U16682 ( .A(n28294), .B(n28295), .C(n28296), .Y(n28293) );
  NOR2X1 U16683 ( .A(n28297), .B(n28298), .Y(n28296) );
  OAI22X1 U16684 ( .A(n25321), .B(n28299), .C(n25332), .D(n28300), .Y(n28298)
         );
  OAI22X1 U16685 ( .A(n25342), .B(n28301), .C(n25353), .D(n28302), .Y(n28297)
         );
  AOI22X1 U16686 ( .A(reg_file[3509]), .B(n25364), .C(reg_file[3381]), .D(
        n25374), .Y(n28295) );
  AOI22X1 U16687 ( .A(reg_file[3253]), .B(n25385), .C(reg_file[3125]), .D(
        n25395), .Y(n28294) );
  NAND3X1 U16688 ( .A(n28303), .B(n28304), .C(n28305), .Y(n28292) );
  NOR2X1 U16689 ( .A(n28306), .B(n28307), .Y(n28305) );
  OAI22X1 U16690 ( .A(n25405), .B(n28308), .C(n25416), .D(n28309), .Y(n28307)
         );
  OAI22X1 U16691 ( .A(n25426), .B(n28310), .C(n25437), .D(n28311), .Y(n28306)
         );
  AOI22X1 U16692 ( .A(reg_file[2485]), .B(n25448), .C(reg_file[2357]), .D(
        n25458), .Y(n28304) );
  AOI22X1 U16693 ( .A(reg_file[2229]), .B(n25469), .C(reg_file[2101]), .D(
        n25479), .Y(n28303) );
  AOI21X1 U16694 ( .A(n28312), .B(n28313), .C(n25143), .Y(rd2data1040_52_) );
  NOR2X1 U16695 ( .A(n28314), .B(n28315), .Y(n28313) );
  NAND3X1 U16696 ( .A(n28316), .B(n28317), .C(n28318), .Y(n28315) );
  NOR2X1 U16697 ( .A(n28319), .B(n28320), .Y(n28318) );
  OAI22X1 U16698 ( .A(n25153), .B(n28321), .C(n25164), .D(n28322), .Y(n28320)
         );
  OAI22X1 U16699 ( .A(n25174), .B(n28323), .C(n25185), .D(n28324), .Y(n28319)
         );
  AOI22X1 U16700 ( .A(reg_file[1460]), .B(n25196), .C(reg_file[1332]), .D(
        n25206), .Y(n28317) );
  AOI22X1 U16701 ( .A(reg_file[1204]), .B(n25217), .C(reg_file[1076]), .D(
        n25227), .Y(n28316) );
  NAND3X1 U16702 ( .A(n28325), .B(n28326), .C(n28327), .Y(n28314) );
  NOR2X1 U16703 ( .A(n28328), .B(n28329), .Y(n28327) );
  OAI22X1 U16704 ( .A(n25237), .B(n28330), .C(n25248), .D(n28331), .Y(n28329)
         );
  OAI22X1 U16705 ( .A(n25258), .B(n28332), .C(n25269), .D(n28333), .Y(n28328)
         );
  AOI22X1 U16706 ( .A(reg_file[564]), .B(n25280), .C(reg_file[692]), .D(n25290), .Y(n28326) );
  AOI22X1 U16707 ( .A(reg_file[820]), .B(n25301), .C(reg_file[948]), .D(n25311), .Y(n28325) );
  NOR2X1 U16708 ( .A(n28334), .B(n28335), .Y(n28312) );
  NAND3X1 U16709 ( .A(n28336), .B(n28337), .C(n28338), .Y(n28335) );
  NOR2X1 U16710 ( .A(n28339), .B(n28340), .Y(n28338) );
  OAI22X1 U16711 ( .A(n25321), .B(n28341), .C(n25332), .D(n28342), .Y(n28340)
         );
  OAI22X1 U16712 ( .A(n25342), .B(n28343), .C(n25353), .D(n28344), .Y(n28339)
         );
  AOI22X1 U16713 ( .A(reg_file[3508]), .B(n25364), .C(reg_file[3380]), .D(
        n25374), .Y(n28337) );
  AOI22X1 U16714 ( .A(reg_file[3252]), .B(n25385), .C(reg_file[3124]), .D(
        n25395), .Y(n28336) );
  NAND3X1 U16715 ( .A(n28345), .B(n28346), .C(n28347), .Y(n28334) );
  NOR2X1 U16716 ( .A(n28348), .B(n28349), .Y(n28347) );
  OAI22X1 U16717 ( .A(n25405), .B(n28350), .C(n25416), .D(n28351), .Y(n28349)
         );
  OAI22X1 U16718 ( .A(n25426), .B(n28352), .C(n25437), .D(n28353), .Y(n28348)
         );
  AOI22X1 U16719 ( .A(reg_file[2484]), .B(n25448), .C(reg_file[2356]), .D(
        n25458), .Y(n28346) );
  AOI22X1 U16720 ( .A(reg_file[2228]), .B(n25469), .C(reg_file[2100]), .D(
        n25479), .Y(n28345) );
  AOI21X1 U16721 ( .A(n28354), .B(n28355), .C(n25143), .Y(rd2data1040_51_) );
  NOR2X1 U16722 ( .A(n28356), .B(n28357), .Y(n28355) );
  NAND3X1 U16723 ( .A(n28358), .B(n28359), .C(n28360), .Y(n28357) );
  NOR2X1 U16724 ( .A(n28361), .B(n28362), .Y(n28360) );
  OAI22X1 U16725 ( .A(n25153), .B(n28363), .C(n25164), .D(n28364), .Y(n28362)
         );
  OAI22X1 U16726 ( .A(n25174), .B(n28365), .C(n25185), .D(n28366), .Y(n28361)
         );
  AOI22X1 U16727 ( .A(reg_file[1459]), .B(n25196), .C(reg_file[1331]), .D(
        n25206), .Y(n28359) );
  AOI22X1 U16728 ( .A(reg_file[1203]), .B(n25217), .C(reg_file[1075]), .D(
        n25227), .Y(n28358) );
  NAND3X1 U16729 ( .A(n28367), .B(n28368), .C(n28369), .Y(n28356) );
  NOR2X1 U16730 ( .A(n28370), .B(n28371), .Y(n28369) );
  OAI22X1 U16731 ( .A(n25237), .B(n28372), .C(n25248), .D(n28373), .Y(n28371)
         );
  OAI22X1 U16732 ( .A(n25258), .B(n28374), .C(n25269), .D(n28375), .Y(n28370)
         );
  AOI22X1 U16733 ( .A(reg_file[563]), .B(n25280), .C(reg_file[691]), .D(n25290), .Y(n28368) );
  AOI22X1 U16734 ( .A(reg_file[819]), .B(n25301), .C(reg_file[947]), .D(n25311), .Y(n28367) );
  NOR2X1 U16735 ( .A(n28376), .B(n28377), .Y(n28354) );
  NAND3X1 U16736 ( .A(n28378), .B(n28379), .C(n28380), .Y(n28377) );
  NOR2X1 U16737 ( .A(n28381), .B(n28382), .Y(n28380) );
  OAI22X1 U16738 ( .A(n25321), .B(n28383), .C(n25332), .D(n28384), .Y(n28382)
         );
  OAI22X1 U16739 ( .A(n25342), .B(n28385), .C(n25353), .D(n28386), .Y(n28381)
         );
  AOI22X1 U16740 ( .A(reg_file[3507]), .B(n25364), .C(reg_file[3379]), .D(
        n25374), .Y(n28379) );
  AOI22X1 U16741 ( .A(reg_file[3251]), .B(n25385), .C(reg_file[3123]), .D(
        n25395), .Y(n28378) );
  NAND3X1 U16742 ( .A(n28387), .B(n28388), .C(n28389), .Y(n28376) );
  NOR2X1 U16743 ( .A(n28390), .B(n28391), .Y(n28389) );
  OAI22X1 U16744 ( .A(n25405), .B(n28392), .C(n25416), .D(n28393), .Y(n28391)
         );
  OAI22X1 U16745 ( .A(n25426), .B(n28394), .C(n25437), .D(n28395), .Y(n28390)
         );
  AOI22X1 U16746 ( .A(reg_file[2483]), .B(n25448), .C(reg_file[2355]), .D(
        n25458), .Y(n28388) );
  AOI22X1 U16747 ( .A(reg_file[2227]), .B(n25469), .C(reg_file[2099]), .D(
        n25479), .Y(n28387) );
  AOI21X1 U16748 ( .A(n28396), .B(n28397), .C(n25143), .Y(rd2data1040_50_) );
  NOR2X1 U16749 ( .A(n28398), .B(n28399), .Y(n28397) );
  NAND3X1 U16750 ( .A(n28400), .B(n28401), .C(n28402), .Y(n28399) );
  NOR2X1 U16751 ( .A(n28403), .B(n28404), .Y(n28402) );
  OAI22X1 U16752 ( .A(n25153), .B(n28405), .C(n25164), .D(n28406), .Y(n28404)
         );
  OAI22X1 U16753 ( .A(n25174), .B(n28407), .C(n25185), .D(n28408), .Y(n28403)
         );
  AOI22X1 U16754 ( .A(reg_file[1458]), .B(n25196), .C(reg_file[1330]), .D(
        n25206), .Y(n28401) );
  AOI22X1 U16755 ( .A(reg_file[1202]), .B(n25217), .C(reg_file[1074]), .D(
        n25227), .Y(n28400) );
  NAND3X1 U16756 ( .A(n28409), .B(n28410), .C(n28411), .Y(n28398) );
  NOR2X1 U16757 ( .A(n28412), .B(n28413), .Y(n28411) );
  OAI22X1 U16758 ( .A(n25237), .B(n28414), .C(n25248), .D(n28415), .Y(n28413)
         );
  OAI22X1 U16759 ( .A(n25258), .B(n28416), .C(n25269), .D(n28417), .Y(n28412)
         );
  AOI22X1 U16760 ( .A(reg_file[562]), .B(n25280), .C(reg_file[690]), .D(n25290), .Y(n28410) );
  AOI22X1 U16761 ( .A(reg_file[818]), .B(n25301), .C(reg_file[946]), .D(n25311), .Y(n28409) );
  NOR2X1 U16762 ( .A(n28418), .B(n28419), .Y(n28396) );
  NAND3X1 U16763 ( .A(n28420), .B(n28421), .C(n28422), .Y(n28419) );
  NOR2X1 U16764 ( .A(n28423), .B(n28424), .Y(n28422) );
  OAI22X1 U16765 ( .A(n25321), .B(n28425), .C(n25332), .D(n28426), .Y(n28424)
         );
  OAI22X1 U16766 ( .A(n25342), .B(n28427), .C(n25353), .D(n28428), .Y(n28423)
         );
  AOI22X1 U16767 ( .A(reg_file[3506]), .B(n25364), .C(reg_file[3378]), .D(
        n25374), .Y(n28421) );
  AOI22X1 U16768 ( .A(reg_file[3250]), .B(n25385), .C(reg_file[3122]), .D(
        n25395), .Y(n28420) );
  NAND3X1 U16769 ( .A(n28429), .B(n28430), .C(n28431), .Y(n28418) );
  NOR2X1 U16770 ( .A(n28432), .B(n28433), .Y(n28431) );
  OAI22X1 U16771 ( .A(n25405), .B(n28434), .C(n25416), .D(n28435), .Y(n28433)
         );
  OAI22X1 U16772 ( .A(n25426), .B(n28436), .C(n25437), .D(n28437), .Y(n28432)
         );
  AOI22X1 U16773 ( .A(reg_file[2482]), .B(n25448), .C(reg_file[2354]), .D(
        n25458), .Y(n28430) );
  AOI22X1 U16774 ( .A(reg_file[2226]), .B(n25469), .C(reg_file[2098]), .D(
        n25479), .Y(n28429) );
  AOI21X1 U16775 ( .A(n28438), .B(n28439), .C(n25143), .Y(rd2data1040_4_) );
  NOR2X1 U16776 ( .A(n28440), .B(n28441), .Y(n28439) );
  NAND3X1 U16777 ( .A(n28442), .B(n28443), .C(n28444), .Y(n28441) );
  NOR2X1 U16778 ( .A(n28445), .B(n28446), .Y(n28444) );
  OAI22X1 U16779 ( .A(n25153), .B(n28447), .C(n25164), .D(n28448), .Y(n28446)
         );
  OAI22X1 U16780 ( .A(n25174), .B(n28449), .C(n25185), .D(n28450), .Y(n28445)
         );
  AOI22X1 U16781 ( .A(reg_file[1412]), .B(n25196), .C(reg_file[1284]), .D(
        n25206), .Y(n28443) );
  AOI22X1 U16782 ( .A(reg_file[1156]), .B(n25217), .C(reg_file[1028]), .D(
        n25227), .Y(n28442) );
  NAND3X1 U16783 ( .A(n28451), .B(n28452), .C(n28453), .Y(n28440) );
  NOR2X1 U16784 ( .A(n28454), .B(n28455), .Y(n28453) );
  OAI22X1 U16785 ( .A(n25237), .B(n28456), .C(n25248), .D(n28457), .Y(n28455)
         );
  OAI22X1 U16786 ( .A(n25258), .B(n28458), .C(n25269), .D(n28459), .Y(n28454)
         );
  AOI22X1 U16787 ( .A(reg_file[516]), .B(n25280), .C(reg_file[644]), .D(n25290), .Y(n28452) );
  AOI22X1 U16788 ( .A(reg_file[772]), .B(n25301), .C(reg_file[900]), .D(n25311), .Y(n28451) );
  NOR2X1 U16789 ( .A(n28460), .B(n28461), .Y(n28438) );
  NAND3X1 U16790 ( .A(n28462), .B(n28463), .C(n28464), .Y(n28461) );
  NOR2X1 U16791 ( .A(n28465), .B(n28466), .Y(n28464) );
  OAI22X1 U16792 ( .A(n25321), .B(n28467), .C(n25332), .D(n28468), .Y(n28466)
         );
  OAI22X1 U16793 ( .A(n25342), .B(n28469), .C(n25353), .D(n28470), .Y(n28465)
         );
  AOI22X1 U16794 ( .A(reg_file[3460]), .B(n25364), .C(reg_file[3332]), .D(
        n25374), .Y(n28463) );
  AOI22X1 U16795 ( .A(reg_file[3204]), .B(n25385), .C(reg_file[3076]), .D(
        n25395), .Y(n28462) );
  NAND3X1 U16796 ( .A(n28471), .B(n28472), .C(n28473), .Y(n28460) );
  NOR2X1 U16797 ( .A(n28474), .B(n28475), .Y(n28473) );
  OAI22X1 U16798 ( .A(n25405), .B(n28476), .C(n25416), .D(n28477), .Y(n28475)
         );
  OAI22X1 U16799 ( .A(n25426), .B(n28478), .C(n25437), .D(n28479), .Y(n28474)
         );
  AOI22X1 U16800 ( .A(reg_file[2436]), .B(n25448), .C(reg_file[2308]), .D(
        n25458), .Y(n28472) );
  AOI22X1 U16801 ( .A(reg_file[2180]), .B(n25469), .C(reg_file[2052]), .D(
        n25479), .Y(n28471) );
  AOI21X1 U16802 ( .A(n28480), .B(n28481), .C(n25142), .Y(rd2data1040_49_) );
  NOR2X1 U16803 ( .A(n28482), .B(n28483), .Y(n28481) );
  NAND3X1 U16804 ( .A(n28484), .B(n28485), .C(n28486), .Y(n28483) );
  NOR2X1 U16805 ( .A(n28487), .B(n28488), .Y(n28486) );
  OAI22X1 U16806 ( .A(n25153), .B(n28489), .C(n25163), .D(n28490), .Y(n28488)
         );
  OAI22X1 U16807 ( .A(n25174), .B(n28491), .C(n25184), .D(n28492), .Y(n28487)
         );
  AOI22X1 U16808 ( .A(reg_file[1457]), .B(n25195), .C(reg_file[1329]), .D(
        n25206), .Y(n28485) );
  AOI22X1 U16809 ( .A(reg_file[1201]), .B(n25216), .C(reg_file[1073]), .D(
        n25227), .Y(n28484) );
  NAND3X1 U16810 ( .A(n28493), .B(n28494), .C(n28495), .Y(n28482) );
  NOR2X1 U16811 ( .A(n28496), .B(n28497), .Y(n28495) );
  OAI22X1 U16812 ( .A(n25237), .B(n28498), .C(n25247), .D(n28499), .Y(n28497)
         );
  OAI22X1 U16813 ( .A(n25258), .B(n28500), .C(n25268), .D(n28501), .Y(n28496)
         );
  AOI22X1 U16814 ( .A(reg_file[561]), .B(n25279), .C(reg_file[689]), .D(n25290), .Y(n28494) );
  AOI22X1 U16815 ( .A(reg_file[817]), .B(n25300), .C(reg_file[945]), .D(n25311), .Y(n28493) );
  NOR2X1 U16816 ( .A(n28502), .B(n28503), .Y(n28480) );
  NAND3X1 U16817 ( .A(n28504), .B(n28505), .C(n28506), .Y(n28503) );
  NOR2X1 U16818 ( .A(n28507), .B(n28508), .Y(n28506) );
  OAI22X1 U16819 ( .A(n25321), .B(n28509), .C(n25331), .D(n28510), .Y(n28508)
         );
  OAI22X1 U16820 ( .A(n25342), .B(n28511), .C(n25352), .D(n28512), .Y(n28507)
         );
  AOI22X1 U16821 ( .A(reg_file[3505]), .B(n25363), .C(reg_file[3377]), .D(
        n25374), .Y(n28505) );
  AOI22X1 U16822 ( .A(reg_file[3249]), .B(n25384), .C(reg_file[3121]), .D(
        n25395), .Y(n28504) );
  NAND3X1 U16823 ( .A(n28513), .B(n28514), .C(n28515), .Y(n28502) );
  NOR2X1 U16824 ( .A(n28516), .B(n28517), .Y(n28515) );
  OAI22X1 U16825 ( .A(n25405), .B(n28518), .C(n25415), .D(n28519), .Y(n28517)
         );
  OAI22X1 U16826 ( .A(n25426), .B(n28520), .C(n25436), .D(n28521), .Y(n28516)
         );
  AOI22X1 U16827 ( .A(reg_file[2481]), .B(n25447), .C(reg_file[2353]), .D(
        n25458), .Y(n28514) );
  AOI22X1 U16828 ( .A(reg_file[2225]), .B(n25468), .C(reg_file[2097]), .D(
        n25479), .Y(n28513) );
  AOI21X1 U16829 ( .A(n28522), .B(n28523), .C(n25142), .Y(rd2data1040_48_) );
  NOR2X1 U16830 ( .A(n28524), .B(n28525), .Y(n28523) );
  NAND3X1 U16831 ( .A(n28526), .B(n28527), .C(n28528), .Y(n28525) );
  NOR2X1 U16832 ( .A(n28529), .B(n28530), .Y(n28528) );
  OAI22X1 U16833 ( .A(n25153), .B(n28531), .C(n25163), .D(n28532), .Y(n28530)
         );
  OAI22X1 U16834 ( .A(n25174), .B(n28533), .C(n25184), .D(n28534), .Y(n28529)
         );
  AOI22X1 U16835 ( .A(reg_file[1456]), .B(n25195), .C(reg_file[1328]), .D(
        n25206), .Y(n28527) );
  AOI22X1 U16836 ( .A(reg_file[1200]), .B(n25216), .C(reg_file[1072]), .D(
        n25227), .Y(n28526) );
  NAND3X1 U16837 ( .A(n28535), .B(n28536), .C(n28537), .Y(n28524) );
  NOR2X1 U16838 ( .A(n28538), .B(n28539), .Y(n28537) );
  OAI22X1 U16839 ( .A(n25237), .B(n28540), .C(n25247), .D(n28541), .Y(n28539)
         );
  OAI22X1 U16840 ( .A(n25258), .B(n28542), .C(n25268), .D(n28543), .Y(n28538)
         );
  AOI22X1 U16841 ( .A(reg_file[560]), .B(n25279), .C(reg_file[688]), .D(n25290), .Y(n28536) );
  AOI22X1 U16842 ( .A(reg_file[816]), .B(n25300), .C(reg_file[944]), .D(n25311), .Y(n28535) );
  NOR2X1 U16843 ( .A(n28544), .B(n28545), .Y(n28522) );
  NAND3X1 U16844 ( .A(n28546), .B(n28547), .C(n28548), .Y(n28545) );
  NOR2X1 U16845 ( .A(n28549), .B(n28550), .Y(n28548) );
  OAI22X1 U16846 ( .A(n25321), .B(n28551), .C(n25331), .D(n28552), .Y(n28550)
         );
  OAI22X1 U16847 ( .A(n25342), .B(n28553), .C(n25352), .D(n28554), .Y(n28549)
         );
  AOI22X1 U16848 ( .A(reg_file[3504]), .B(n25363), .C(reg_file[3376]), .D(
        n25374), .Y(n28547) );
  AOI22X1 U16849 ( .A(reg_file[3248]), .B(n25384), .C(reg_file[3120]), .D(
        n25395), .Y(n28546) );
  NAND3X1 U16850 ( .A(n28555), .B(n28556), .C(n28557), .Y(n28544) );
  NOR2X1 U16851 ( .A(n28558), .B(n28559), .Y(n28557) );
  OAI22X1 U16852 ( .A(n25405), .B(n28560), .C(n25415), .D(n28561), .Y(n28559)
         );
  OAI22X1 U16853 ( .A(n25426), .B(n28562), .C(n25436), .D(n28563), .Y(n28558)
         );
  AOI22X1 U16854 ( .A(reg_file[2480]), .B(n25447), .C(reg_file[2352]), .D(
        n25458), .Y(n28556) );
  AOI22X1 U16855 ( .A(reg_file[2224]), .B(n25468), .C(reg_file[2096]), .D(
        n25479), .Y(n28555) );
  AOI21X1 U16856 ( .A(n28564), .B(n28565), .C(n25142), .Y(rd2data1040_47_) );
  NOR2X1 U16857 ( .A(n28566), .B(n28567), .Y(n28565) );
  NAND3X1 U16858 ( .A(n28568), .B(n28569), .C(n28570), .Y(n28567) );
  NOR2X1 U16859 ( .A(n28571), .B(n28572), .Y(n28570) );
  OAI22X1 U16860 ( .A(n25153), .B(n28573), .C(n25163), .D(n28574), .Y(n28572)
         );
  OAI22X1 U16861 ( .A(n25174), .B(n28575), .C(n25184), .D(n28576), .Y(n28571)
         );
  AOI22X1 U16862 ( .A(reg_file[1455]), .B(n25195), .C(reg_file[1327]), .D(
        n25206), .Y(n28569) );
  AOI22X1 U16863 ( .A(reg_file[1199]), .B(n25216), .C(reg_file[1071]), .D(
        n25227), .Y(n28568) );
  NAND3X1 U16864 ( .A(n28577), .B(n28578), .C(n28579), .Y(n28566) );
  NOR2X1 U16865 ( .A(n28580), .B(n28581), .Y(n28579) );
  OAI22X1 U16866 ( .A(n25237), .B(n28582), .C(n25247), .D(n28583), .Y(n28581)
         );
  OAI22X1 U16867 ( .A(n25258), .B(n28584), .C(n25268), .D(n28585), .Y(n28580)
         );
  AOI22X1 U16868 ( .A(reg_file[559]), .B(n25279), .C(reg_file[687]), .D(n25290), .Y(n28578) );
  AOI22X1 U16869 ( .A(reg_file[815]), .B(n25300), .C(reg_file[943]), .D(n25311), .Y(n28577) );
  NOR2X1 U16870 ( .A(n28586), .B(n28587), .Y(n28564) );
  NAND3X1 U16871 ( .A(n28588), .B(n28589), .C(n28590), .Y(n28587) );
  NOR2X1 U16872 ( .A(n28591), .B(n28592), .Y(n28590) );
  OAI22X1 U16873 ( .A(n25321), .B(n28593), .C(n25331), .D(n28594), .Y(n28592)
         );
  OAI22X1 U16874 ( .A(n25342), .B(n28595), .C(n25352), .D(n28596), .Y(n28591)
         );
  AOI22X1 U16875 ( .A(reg_file[3503]), .B(n25363), .C(reg_file[3375]), .D(
        n25374), .Y(n28589) );
  AOI22X1 U16876 ( .A(reg_file[3247]), .B(n25384), .C(reg_file[3119]), .D(
        n25395), .Y(n28588) );
  NAND3X1 U16877 ( .A(n28597), .B(n28598), .C(n28599), .Y(n28586) );
  NOR2X1 U16878 ( .A(n28600), .B(n28601), .Y(n28599) );
  OAI22X1 U16879 ( .A(n25405), .B(n28602), .C(n25415), .D(n28603), .Y(n28601)
         );
  OAI22X1 U16880 ( .A(n25426), .B(n28604), .C(n25436), .D(n28605), .Y(n28600)
         );
  AOI22X1 U16881 ( .A(reg_file[2479]), .B(n25447), .C(reg_file[2351]), .D(
        n25458), .Y(n28598) );
  AOI22X1 U16882 ( .A(reg_file[2223]), .B(n25468), .C(reg_file[2095]), .D(
        n25479), .Y(n28597) );
  AOI21X1 U16883 ( .A(n28606), .B(n28607), .C(n25142), .Y(rd2data1040_46_) );
  NOR2X1 U16884 ( .A(n28608), .B(n28609), .Y(n28607) );
  NAND3X1 U16885 ( .A(n28610), .B(n28611), .C(n28612), .Y(n28609) );
  NOR2X1 U16886 ( .A(n28613), .B(n28614), .Y(n28612) );
  OAI22X1 U16887 ( .A(n25153), .B(n28615), .C(n25163), .D(n28616), .Y(n28614)
         );
  OAI22X1 U16888 ( .A(n25174), .B(n28617), .C(n25184), .D(n28618), .Y(n28613)
         );
  AOI22X1 U16889 ( .A(reg_file[1454]), .B(n25195), .C(reg_file[1326]), .D(
        n25206), .Y(n28611) );
  AOI22X1 U16890 ( .A(reg_file[1198]), .B(n25216), .C(reg_file[1070]), .D(
        n25227), .Y(n28610) );
  NAND3X1 U16891 ( .A(n28619), .B(n28620), .C(n28621), .Y(n28608) );
  NOR2X1 U16892 ( .A(n28622), .B(n28623), .Y(n28621) );
  OAI22X1 U16893 ( .A(n25237), .B(n28624), .C(n25247), .D(n28625), .Y(n28623)
         );
  OAI22X1 U16894 ( .A(n25258), .B(n28626), .C(n25268), .D(n28627), .Y(n28622)
         );
  AOI22X1 U16895 ( .A(reg_file[558]), .B(n25279), .C(reg_file[686]), .D(n25290), .Y(n28620) );
  AOI22X1 U16896 ( .A(reg_file[814]), .B(n25300), .C(reg_file[942]), .D(n25311), .Y(n28619) );
  NOR2X1 U16897 ( .A(n28628), .B(n28629), .Y(n28606) );
  NAND3X1 U16898 ( .A(n28630), .B(n28631), .C(n28632), .Y(n28629) );
  NOR2X1 U16899 ( .A(n28633), .B(n28634), .Y(n28632) );
  OAI22X1 U16900 ( .A(n25321), .B(n28635), .C(n25331), .D(n28636), .Y(n28634)
         );
  OAI22X1 U16901 ( .A(n25342), .B(n28637), .C(n25352), .D(n28638), .Y(n28633)
         );
  AOI22X1 U16902 ( .A(reg_file[3502]), .B(n25363), .C(reg_file[3374]), .D(
        n25374), .Y(n28631) );
  AOI22X1 U16903 ( .A(reg_file[3246]), .B(n25384), .C(reg_file[3118]), .D(
        n25395), .Y(n28630) );
  NAND3X1 U16904 ( .A(n28639), .B(n28640), .C(n28641), .Y(n28628) );
  NOR2X1 U16905 ( .A(n28642), .B(n28643), .Y(n28641) );
  OAI22X1 U16906 ( .A(n25405), .B(n28644), .C(n25415), .D(n28645), .Y(n28643)
         );
  OAI22X1 U16907 ( .A(n25426), .B(n28646), .C(n25436), .D(n28647), .Y(n28642)
         );
  AOI22X1 U16908 ( .A(reg_file[2478]), .B(n25447), .C(reg_file[2350]), .D(
        n25458), .Y(n28640) );
  AOI22X1 U16909 ( .A(reg_file[2222]), .B(n25468), .C(reg_file[2094]), .D(
        n25479), .Y(n28639) );
  AOI21X1 U16910 ( .A(n28648), .B(n28649), .C(n25142), .Y(rd2data1040_45_) );
  NOR2X1 U16911 ( .A(n28650), .B(n28651), .Y(n28649) );
  NAND3X1 U16912 ( .A(n28652), .B(n28653), .C(n28654), .Y(n28651) );
  NOR2X1 U16913 ( .A(n28655), .B(n28656), .Y(n28654) );
  OAI22X1 U16914 ( .A(n25153), .B(n28657), .C(n25163), .D(n28658), .Y(n28656)
         );
  OAI22X1 U16915 ( .A(n25174), .B(n28659), .C(n25184), .D(n28660), .Y(n28655)
         );
  AOI22X1 U16916 ( .A(reg_file[1453]), .B(n25195), .C(reg_file[1325]), .D(
        n25206), .Y(n28653) );
  AOI22X1 U16917 ( .A(reg_file[1197]), .B(n25216), .C(reg_file[1069]), .D(
        n25227), .Y(n28652) );
  NAND3X1 U16918 ( .A(n28661), .B(n28662), .C(n28663), .Y(n28650) );
  NOR2X1 U16919 ( .A(n28664), .B(n28665), .Y(n28663) );
  OAI22X1 U16920 ( .A(n25237), .B(n28666), .C(n25247), .D(n28667), .Y(n28665)
         );
  OAI22X1 U16921 ( .A(n25258), .B(n28668), .C(n25268), .D(n28669), .Y(n28664)
         );
  AOI22X1 U16922 ( .A(reg_file[557]), .B(n25279), .C(reg_file[685]), .D(n25290), .Y(n28662) );
  AOI22X1 U16923 ( .A(reg_file[813]), .B(n25300), .C(reg_file[941]), .D(n25311), .Y(n28661) );
  NOR2X1 U16924 ( .A(n28670), .B(n28671), .Y(n28648) );
  NAND3X1 U16925 ( .A(n28672), .B(n28673), .C(n28674), .Y(n28671) );
  NOR2X1 U16926 ( .A(n28675), .B(n28676), .Y(n28674) );
  OAI22X1 U16927 ( .A(n25321), .B(n28677), .C(n25331), .D(n28678), .Y(n28676)
         );
  OAI22X1 U16928 ( .A(n25342), .B(n28679), .C(n25352), .D(n28680), .Y(n28675)
         );
  AOI22X1 U16929 ( .A(reg_file[3501]), .B(n25363), .C(reg_file[3373]), .D(
        n25374), .Y(n28673) );
  AOI22X1 U16930 ( .A(reg_file[3245]), .B(n25384), .C(reg_file[3117]), .D(
        n25395), .Y(n28672) );
  NAND3X1 U16931 ( .A(n28681), .B(n28682), .C(n28683), .Y(n28670) );
  NOR2X1 U16932 ( .A(n28684), .B(n28685), .Y(n28683) );
  OAI22X1 U16933 ( .A(n25405), .B(n28686), .C(n25415), .D(n28687), .Y(n28685)
         );
  OAI22X1 U16934 ( .A(n25426), .B(n28688), .C(n25436), .D(n28689), .Y(n28684)
         );
  AOI22X1 U16935 ( .A(reg_file[2477]), .B(n25447), .C(reg_file[2349]), .D(
        n25458), .Y(n28682) );
  AOI22X1 U16936 ( .A(reg_file[2221]), .B(n25468), .C(reg_file[2093]), .D(
        n25479), .Y(n28681) );
  AOI21X1 U16937 ( .A(n28690), .B(n28691), .C(n25142), .Y(rd2data1040_44_) );
  NOR2X1 U16938 ( .A(n28692), .B(n28693), .Y(n28691) );
  NAND3X1 U16939 ( .A(n28694), .B(n28695), .C(n28696), .Y(n28693) );
  NOR2X1 U16940 ( .A(n28697), .B(n28698), .Y(n28696) );
  OAI22X1 U16941 ( .A(n25153), .B(n28699), .C(n25163), .D(n28700), .Y(n28698)
         );
  OAI22X1 U16942 ( .A(n25174), .B(n28701), .C(n25184), .D(n28702), .Y(n28697)
         );
  AOI22X1 U16943 ( .A(reg_file[1452]), .B(n25195), .C(reg_file[1324]), .D(
        n25206), .Y(n28695) );
  AOI22X1 U16944 ( .A(reg_file[1196]), .B(n25216), .C(reg_file[1068]), .D(
        n25227), .Y(n28694) );
  NAND3X1 U16945 ( .A(n28703), .B(n28704), .C(n28705), .Y(n28692) );
  NOR2X1 U16946 ( .A(n28706), .B(n28707), .Y(n28705) );
  OAI22X1 U16947 ( .A(n25237), .B(n28708), .C(n25247), .D(n28709), .Y(n28707)
         );
  OAI22X1 U16948 ( .A(n25258), .B(n28710), .C(n25268), .D(n28711), .Y(n28706)
         );
  AOI22X1 U16949 ( .A(reg_file[556]), .B(n25279), .C(reg_file[684]), .D(n25290), .Y(n28704) );
  AOI22X1 U16950 ( .A(reg_file[812]), .B(n25300), .C(reg_file[940]), .D(n25311), .Y(n28703) );
  NOR2X1 U16951 ( .A(n28712), .B(n28713), .Y(n28690) );
  NAND3X1 U16952 ( .A(n28714), .B(n28715), .C(n28716), .Y(n28713) );
  NOR2X1 U16953 ( .A(n28717), .B(n28718), .Y(n28716) );
  OAI22X1 U16954 ( .A(n25321), .B(n28719), .C(n25331), .D(n28720), .Y(n28718)
         );
  OAI22X1 U16955 ( .A(n25342), .B(n28721), .C(n25352), .D(n28722), .Y(n28717)
         );
  AOI22X1 U16956 ( .A(reg_file[3500]), .B(n25363), .C(reg_file[3372]), .D(
        n25374), .Y(n28715) );
  AOI22X1 U16957 ( .A(reg_file[3244]), .B(n25384), .C(reg_file[3116]), .D(
        n25395), .Y(n28714) );
  NAND3X1 U16958 ( .A(n28723), .B(n28724), .C(n28725), .Y(n28712) );
  NOR2X1 U16959 ( .A(n28726), .B(n28727), .Y(n28725) );
  OAI22X1 U16960 ( .A(n25405), .B(n28728), .C(n25415), .D(n28729), .Y(n28727)
         );
  OAI22X1 U16961 ( .A(n25426), .B(n28730), .C(n25436), .D(n28731), .Y(n28726)
         );
  AOI22X1 U16962 ( .A(reg_file[2476]), .B(n25447), .C(reg_file[2348]), .D(
        n25458), .Y(n28724) );
  AOI22X1 U16963 ( .A(reg_file[2220]), .B(n25468), .C(reg_file[2092]), .D(
        n25479), .Y(n28723) );
  AOI21X1 U16964 ( .A(n28732), .B(n28733), .C(n25142), .Y(rd2data1040_43_) );
  NOR2X1 U16965 ( .A(n28734), .B(n28735), .Y(n28733) );
  NAND3X1 U16966 ( .A(n28736), .B(n28737), .C(n28738), .Y(n28735) );
  NOR2X1 U16967 ( .A(n28739), .B(n28740), .Y(n28738) );
  OAI22X1 U16968 ( .A(n25153), .B(n28741), .C(n25163), .D(n28742), .Y(n28740)
         );
  OAI22X1 U16969 ( .A(n25174), .B(n28743), .C(n25184), .D(n28744), .Y(n28739)
         );
  AOI22X1 U16970 ( .A(reg_file[1451]), .B(n25195), .C(reg_file[1323]), .D(
        n25206), .Y(n28737) );
  AOI22X1 U16971 ( .A(reg_file[1195]), .B(n25216), .C(reg_file[1067]), .D(
        n25227), .Y(n28736) );
  NAND3X1 U16972 ( .A(n28745), .B(n28746), .C(n28747), .Y(n28734) );
  NOR2X1 U16973 ( .A(n28748), .B(n28749), .Y(n28747) );
  OAI22X1 U16974 ( .A(n25237), .B(n28750), .C(n25247), .D(n28751), .Y(n28749)
         );
  OAI22X1 U16975 ( .A(n25258), .B(n28752), .C(n25268), .D(n28753), .Y(n28748)
         );
  AOI22X1 U16976 ( .A(reg_file[555]), .B(n25279), .C(reg_file[683]), .D(n25290), .Y(n28746) );
  AOI22X1 U16977 ( .A(reg_file[811]), .B(n25300), .C(reg_file[939]), .D(n25311), .Y(n28745) );
  NOR2X1 U16978 ( .A(n28754), .B(n28755), .Y(n28732) );
  NAND3X1 U16979 ( .A(n28756), .B(n28757), .C(n28758), .Y(n28755) );
  NOR2X1 U16980 ( .A(n28759), .B(n28760), .Y(n28758) );
  OAI22X1 U16981 ( .A(n25321), .B(n28761), .C(n25331), .D(n28762), .Y(n28760)
         );
  OAI22X1 U16982 ( .A(n25342), .B(n28763), .C(n25352), .D(n28764), .Y(n28759)
         );
  AOI22X1 U16983 ( .A(reg_file[3499]), .B(n25363), .C(reg_file[3371]), .D(
        n25374), .Y(n28757) );
  AOI22X1 U16984 ( .A(reg_file[3243]), .B(n25384), .C(reg_file[3115]), .D(
        n25395), .Y(n28756) );
  NAND3X1 U16985 ( .A(n28765), .B(n28766), .C(n28767), .Y(n28754) );
  NOR2X1 U16986 ( .A(n28768), .B(n28769), .Y(n28767) );
  OAI22X1 U16987 ( .A(n25405), .B(n28770), .C(n25415), .D(n28771), .Y(n28769)
         );
  OAI22X1 U16988 ( .A(n25426), .B(n28772), .C(n25436), .D(n28773), .Y(n28768)
         );
  AOI22X1 U16989 ( .A(reg_file[2475]), .B(n25447), .C(reg_file[2347]), .D(
        n25458), .Y(n28766) );
  AOI22X1 U16990 ( .A(reg_file[2219]), .B(n25468), .C(reg_file[2091]), .D(
        n25479), .Y(n28765) );
  AOI21X1 U16991 ( .A(n28774), .B(n28775), .C(n25142), .Y(rd2data1040_42_) );
  NOR2X1 U16992 ( .A(n28776), .B(n28777), .Y(n28775) );
  NAND3X1 U16993 ( .A(n28778), .B(n28779), .C(n28780), .Y(n28777) );
  NOR2X1 U16994 ( .A(n28781), .B(n28782), .Y(n28780) );
  OAI22X1 U16995 ( .A(n25152), .B(n28783), .C(n25163), .D(n28784), .Y(n28782)
         );
  OAI22X1 U16996 ( .A(n25173), .B(n28785), .C(n25184), .D(n28786), .Y(n28781)
         );
  AOI22X1 U16997 ( .A(reg_file[1450]), .B(n25195), .C(reg_file[1322]), .D(
        n25205), .Y(n28779) );
  AOI22X1 U16998 ( .A(reg_file[1194]), .B(n25216), .C(reg_file[1066]), .D(
        n25226), .Y(n28778) );
  NAND3X1 U16999 ( .A(n28787), .B(n28788), .C(n28789), .Y(n28776) );
  NOR2X1 U17000 ( .A(n28790), .B(n28791), .Y(n28789) );
  OAI22X1 U17001 ( .A(n25236), .B(n28792), .C(n25247), .D(n28793), .Y(n28791)
         );
  OAI22X1 U17002 ( .A(n25257), .B(n28794), .C(n25268), .D(n28795), .Y(n28790)
         );
  AOI22X1 U17003 ( .A(reg_file[554]), .B(n25279), .C(reg_file[682]), .D(n25289), .Y(n28788) );
  AOI22X1 U17004 ( .A(reg_file[810]), .B(n25300), .C(reg_file[938]), .D(n25310), .Y(n28787) );
  NOR2X1 U17005 ( .A(n28796), .B(n28797), .Y(n28774) );
  NAND3X1 U17006 ( .A(n28798), .B(n28799), .C(n28800), .Y(n28797) );
  NOR2X1 U17007 ( .A(n28801), .B(n28802), .Y(n28800) );
  OAI22X1 U17008 ( .A(n25320), .B(n28803), .C(n25331), .D(n28804), .Y(n28802)
         );
  OAI22X1 U17009 ( .A(n25341), .B(n28805), .C(n25352), .D(n28806), .Y(n28801)
         );
  AOI22X1 U17010 ( .A(reg_file[3498]), .B(n25363), .C(reg_file[3370]), .D(
        n25373), .Y(n28799) );
  AOI22X1 U17011 ( .A(reg_file[3242]), .B(n25384), .C(reg_file[3114]), .D(
        n25394), .Y(n28798) );
  NAND3X1 U17012 ( .A(n28807), .B(n28808), .C(n28809), .Y(n28796) );
  NOR2X1 U17013 ( .A(n28810), .B(n28811), .Y(n28809) );
  OAI22X1 U17014 ( .A(n25404), .B(n28812), .C(n25415), .D(n28813), .Y(n28811)
         );
  OAI22X1 U17015 ( .A(n25425), .B(n28814), .C(n25436), .D(n28815), .Y(n28810)
         );
  AOI22X1 U17016 ( .A(reg_file[2474]), .B(n25447), .C(reg_file[2346]), .D(
        n25457), .Y(n28808) );
  AOI22X1 U17017 ( .A(reg_file[2218]), .B(n25468), .C(reg_file[2090]), .D(
        n25478), .Y(n28807) );
  AOI21X1 U17018 ( .A(n28816), .B(n28817), .C(n25142), .Y(rd2data1040_41_) );
  NOR2X1 U17019 ( .A(n28818), .B(n28819), .Y(n28817) );
  NAND3X1 U17020 ( .A(n28820), .B(n28821), .C(n28822), .Y(n28819) );
  NOR2X1 U17021 ( .A(n28823), .B(n28824), .Y(n28822) );
  OAI22X1 U17022 ( .A(n25152), .B(n28825), .C(n25163), .D(n28826), .Y(n28824)
         );
  OAI22X1 U17023 ( .A(n25173), .B(n28827), .C(n25184), .D(n28828), .Y(n28823)
         );
  AOI22X1 U17024 ( .A(reg_file[1449]), .B(n25195), .C(reg_file[1321]), .D(
        n25205), .Y(n28821) );
  AOI22X1 U17025 ( .A(reg_file[1193]), .B(n25216), .C(reg_file[1065]), .D(
        n25226), .Y(n28820) );
  NAND3X1 U17026 ( .A(n28829), .B(n28830), .C(n28831), .Y(n28818) );
  NOR2X1 U17027 ( .A(n28832), .B(n28833), .Y(n28831) );
  OAI22X1 U17028 ( .A(n25236), .B(n28834), .C(n25247), .D(n28835), .Y(n28833)
         );
  OAI22X1 U17029 ( .A(n25257), .B(n28836), .C(n25268), .D(n28837), .Y(n28832)
         );
  AOI22X1 U17030 ( .A(reg_file[553]), .B(n25279), .C(reg_file[681]), .D(n25289), .Y(n28830) );
  AOI22X1 U17031 ( .A(reg_file[809]), .B(n25300), .C(reg_file[937]), .D(n25310), .Y(n28829) );
  NOR2X1 U17032 ( .A(n28838), .B(n28839), .Y(n28816) );
  NAND3X1 U17033 ( .A(n28840), .B(n28841), .C(n28842), .Y(n28839) );
  NOR2X1 U17034 ( .A(n28843), .B(n28844), .Y(n28842) );
  OAI22X1 U17035 ( .A(n25320), .B(n28845), .C(n25331), .D(n28846), .Y(n28844)
         );
  OAI22X1 U17036 ( .A(n25341), .B(n28847), .C(n25352), .D(n28848), .Y(n28843)
         );
  AOI22X1 U17037 ( .A(reg_file[3497]), .B(n25363), .C(reg_file[3369]), .D(
        n25373), .Y(n28841) );
  AOI22X1 U17038 ( .A(reg_file[3241]), .B(n25384), .C(reg_file[3113]), .D(
        n25394), .Y(n28840) );
  NAND3X1 U17039 ( .A(n28849), .B(n28850), .C(n28851), .Y(n28838) );
  NOR2X1 U17040 ( .A(n28852), .B(n28853), .Y(n28851) );
  OAI22X1 U17041 ( .A(n25404), .B(n28854), .C(n25415), .D(n28855), .Y(n28853)
         );
  OAI22X1 U17042 ( .A(n25425), .B(n28856), .C(n25436), .D(n28857), .Y(n28852)
         );
  AOI22X1 U17043 ( .A(reg_file[2473]), .B(n25447), .C(reg_file[2345]), .D(
        n25457), .Y(n28850) );
  AOI22X1 U17044 ( .A(reg_file[2217]), .B(n25468), .C(reg_file[2089]), .D(
        n25478), .Y(n28849) );
  AOI21X1 U17045 ( .A(n28858), .B(n28859), .C(n25142), .Y(rd2data1040_40_) );
  NOR2X1 U17046 ( .A(n28860), .B(n28861), .Y(n28859) );
  NAND3X1 U17047 ( .A(n28862), .B(n28863), .C(n28864), .Y(n28861) );
  NOR2X1 U17048 ( .A(n28865), .B(n28866), .Y(n28864) );
  OAI22X1 U17049 ( .A(n25152), .B(n28867), .C(n25163), .D(n28868), .Y(n28866)
         );
  OAI22X1 U17050 ( .A(n25173), .B(n28869), .C(n25184), .D(n28870), .Y(n28865)
         );
  AOI22X1 U17051 ( .A(reg_file[1448]), .B(n25195), .C(reg_file[1320]), .D(
        n25205), .Y(n28863) );
  AOI22X1 U17052 ( .A(reg_file[1192]), .B(n25216), .C(reg_file[1064]), .D(
        n25226), .Y(n28862) );
  NAND3X1 U17053 ( .A(n28871), .B(n28872), .C(n28873), .Y(n28860) );
  NOR2X1 U17054 ( .A(n28874), .B(n28875), .Y(n28873) );
  OAI22X1 U17055 ( .A(n25236), .B(n28876), .C(n25247), .D(n28877), .Y(n28875)
         );
  OAI22X1 U17056 ( .A(n25257), .B(n28878), .C(n25268), .D(n28879), .Y(n28874)
         );
  AOI22X1 U17057 ( .A(reg_file[552]), .B(n25279), .C(reg_file[680]), .D(n25289), .Y(n28872) );
  AOI22X1 U17058 ( .A(reg_file[808]), .B(n25300), .C(reg_file[936]), .D(n25310), .Y(n28871) );
  NOR2X1 U17059 ( .A(n28880), .B(n28881), .Y(n28858) );
  NAND3X1 U17060 ( .A(n28882), .B(n28883), .C(n28884), .Y(n28881) );
  NOR2X1 U17061 ( .A(n28885), .B(n28886), .Y(n28884) );
  OAI22X1 U17062 ( .A(n25320), .B(n28887), .C(n25331), .D(n28888), .Y(n28886)
         );
  OAI22X1 U17063 ( .A(n25341), .B(n28889), .C(n25352), .D(n28890), .Y(n28885)
         );
  AOI22X1 U17064 ( .A(reg_file[3496]), .B(n25363), .C(reg_file[3368]), .D(
        n25373), .Y(n28883) );
  AOI22X1 U17065 ( .A(reg_file[3240]), .B(n25384), .C(reg_file[3112]), .D(
        n25394), .Y(n28882) );
  NAND3X1 U17066 ( .A(n28891), .B(n28892), .C(n28893), .Y(n28880) );
  NOR2X1 U17067 ( .A(n28894), .B(n28895), .Y(n28893) );
  OAI22X1 U17068 ( .A(n25404), .B(n28896), .C(n25415), .D(n28897), .Y(n28895)
         );
  OAI22X1 U17069 ( .A(n25425), .B(n28898), .C(n25436), .D(n28899), .Y(n28894)
         );
  AOI22X1 U17070 ( .A(reg_file[2472]), .B(n25447), .C(reg_file[2344]), .D(
        n25457), .Y(n28892) );
  AOI22X1 U17071 ( .A(reg_file[2216]), .B(n25468), .C(reg_file[2088]), .D(
        n25478), .Y(n28891) );
  AOI21X1 U17072 ( .A(n28900), .B(n28901), .C(n25142), .Y(rd2data1040_3_) );
  NOR2X1 U17073 ( .A(n28902), .B(n28903), .Y(n28901) );
  NAND3X1 U17074 ( .A(n28904), .B(n28905), .C(n28906), .Y(n28903) );
  NOR2X1 U17075 ( .A(n28907), .B(n28908), .Y(n28906) );
  OAI22X1 U17076 ( .A(n25152), .B(n28909), .C(n25163), .D(n28910), .Y(n28908)
         );
  OAI22X1 U17077 ( .A(n25173), .B(n28911), .C(n25184), .D(n28912), .Y(n28907)
         );
  AOI22X1 U17078 ( .A(reg_file[1411]), .B(n25195), .C(reg_file[1283]), .D(
        n25205), .Y(n28905) );
  AOI22X1 U17079 ( .A(reg_file[1155]), .B(n25216), .C(reg_file[1027]), .D(
        n25226), .Y(n28904) );
  NAND3X1 U17080 ( .A(n28913), .B(n28914), .C(n28915), .Y(n28902) );
  NOR2X1 U17081 ( .A(n28916), .B(n28917), .Y(n28915) );
  OAI22X1 U17082 ( .A(n25236), .B(n28918), .C(n25247), .D(n28919), .Y(n28917)
         );
  OAI22X1 U17083 ( .A(n25257), .B(n28920), .C(n25268), .D(n28921), .Y(n28916)
         );
  AOI22X1 U17084 ( .A(reg_file[515]), .B(n25279), .C(reg_file[643]), .D(n25289), .Y(n28914) );
  AOI22X1 U17085 ( .A(reg_file[771]), .B(n25300), .C(reg_file[899]), .D(n25310), .Y(n28913) );
  NOR2X1 U17086 ( .A(n28922), .B(n28923), .Y(n28900) );
  NAND3X1 U17087 ( .A(n28924), .B(n28925), .C(n28926), .Y(n28923) );
  NOR2X1 U17088 ( .A(n28927), .B(n28928), .Y(n28926) );
  OAI22X1 U17089 ( .A(n25320), .B(n28929), .C(n25331), .D(n28930), .Y(n28928)
         );
  OAI22X1 U17090 ( .A(n25341), .B(n28931), .C(n25352), .D(n28932), .Y(n28927)
         );
  AOI22X1 U17091 ( .A(reg_file[3459]), .B(n25363), .C(reg_file[3331]), .D(
        n25373), .Y(n28925) );
  AOI22X1 U17092 ( .A(reg_file[3203]), .B(n25384), .C(reg_file[3075]), .D(
        n25394), .Y(n28924) );
  NAND3X1 U17093 ( .A(n28933), .B(n28934), .C(n28935), .Y(n28922) );
  NOR2X1 U17094 ( .A(n28936), .B(n28937), .Y(n28935) );
  OAI22X1 U17095 ( .A(n25404), .B(n28938), .C(n25415), .D(n28939), .Y(n28937)
         );
  OAI22X1 U17096 ( .A(n25425), .B(n28940), .C(n25436), .D(n28941), .Y(n28936)
         );
  AOI22X1 U17097 ( .A(reg_file[2435]), .B(n25447), .C(reg_file[2307]), .D(
        n25457), .Y(n28934) );
  AOI22X1 U17098 ( .A(reg_file[2179]), .B(n25468), .C(reg_file[2051]), .D(
        n25478), .Y(n28933) );
  AOI21X1 U17099 ( .A(n28942), .B(n28943), .C(n25142), .Y(rd2data1040_39_) );
  NOR2X1 U17100 ( .A(n28944), .B(n28945), .Y(n28943) );
  NAND3X1 U17101 ( .A(n28946), .B(n28947), .C(n28948), .Y(n28945) );
  NOR2X1 U17102 ( .A(n28949), .B(n28950), .Y(n28948) );
  OAI22X1 U17103 ( .A(n25152), .B(n28951), .C(n25163), .D(n28952), .Y(n28950)
         );
  OAI22X1 U17104 ( .A(n25173), .B(n28953), .C(n25184), .D(n28954), .Y(n28949)
         );
  AOI22X1 U17105 ( .A(reg_file[1447]), .B(n25195), .C(reg_file[1319]), .D(
        n25205), .Y(n28947) );
  AOI22X1 U17106 ( .A(reg_file[1191]), .B(n25216), .C(reg_file[1063]), .D(
        n25226), .Y(n28946) );
  NAND3X1 U17107 ( .A(n28955), .B(n28956), .C(n28957), .Y(n28944) );
  NOR2X1 U17108 ( .A(n28958), .B(n28959), .Y(n28957) );
  OAI22X1 U17109 ( .A(n25236), .B(n28960), .C(n25247), .D(n28961), .Y(n28959)
         );
  OAI22X1 U17110 ( .A(n25257), .B(n28962), .C(n25268), .D(n28963), .Y(n28958)
         );
  AOI22X1 U17111 ( .A(reg_file[551]), .B(n25279), .C(reg_file[679]), .D(n25289), .Y(n28956) );
  AOI22X1 U17112 ( .A(reg_file[807]), .B(n25300), .C(reg_file[935]), .D(n25310), .Y(n28955) );
  NOR2X1 U17113 ( .A(n28964), .B(n28965), .Y(n28942) );
  NAND3X1 U17114 ( .A(n28966), .B(n28967), .C(n28968), .Y(n28965) );
  NOR2X1 U17115 ( .A(n28969), .B(n28970), .Y(n28968) );
  OAI22X1 U17116 ( .A(n25320), .B(n28971), .C(n25331), .D(n28972), .Y(n28970)
         );
  OAI22X1 U17117 ( .A(n25341), .B(n28973), .C(n25352), .D(n28974), .Y(n28969)
         );
  AOI22X1 U17118 ( .A(reg_file[3495]), .B(n25363), .C(reg_file[3367]), .D(
        n25373), .Y(n28967) );
  AOI22X1 U17119 ( .A(reg_file[3239]), .B(n25384), .C(reg_file[3111]), .D(
        n25394), .Y(n28966) );
  NAND3X1 U17120 ( .A(n28975), .B(n28976), .C(n28977), .Y(n28964) );
  NOR2X1 U17121 ( .A(n28978), .B(n28979), .Y(n28977) );
  OAI22X1 U17122 ( .A(n25404), .B(n28980), .C(n25415), .D(n28981), .Y(n28979)
         );
  OAI22X1 U17123 ( .A(n25425), .B(n28982), .C(n25436), .D(n28983), .Y(n28978)
         );
  AOI22X1 U17124 ( .A(reg_file[2471]), .B(n25447), .C(reg_file[2343]), .D(
        n25457), .Y(n28976) );
  AOI22X1 U17125 ( .A(reg_file[2215]), .B(n25468), .C(reg_file[2087]), .D(
        n25478), .Y(n28975) );
  AOI21X1 U17126 ( .A(n28984), .B(n28985), .C(n25141), .Y(rd2data1040_38_) );
  NOR2X1 U17127 ( .A(n28986), .B(n28987), .Y(n28985) );
  NAND3X1 U17128 ( .A(n28988), .B(n28989), .C(n28990), .Y(n28987) );
  NOR2X1 U17129 ( .A(n28991), .B(n28992), .Y(n28990) );
  OAI22X1 U17130 ( .A(n25152), .B(n28993), .C(n25162), .D(n28994), .Y(n28992)
         );
  OAI22X1 U17131 ( .A(n25173), .B(n28995), .C(n25183), .D(n28996), .Y(n28991)
         );
  AOI22X1 U17132 ( .A(reg_file[1446]), .B(n25194), .C(reg_file[1318]), .D(
        n25205), .Y(n28989) );
  AOI22X1 U17133 ( .A(reg_file[1190]), .B(n25215), .C(reg_file[1062]), .D(
        n25226), .Y(n28988) );
  NAND3X1 U17134 ( .A(n28997), .B(n28998), .C(n28999), .Y(n28986) );
  NOR2X1 U17135 ( .A(n29000), .B(n29001), .Y(n28999) );
  OAI22X1 U17136 ( .A(n25236), .B(n29002), .C(n25246), .D(n29003), .Y(n29001)
         );
  OAI22X1 U17137 ( .A(n25257), .B(n29004), .C(n25267), .D(n29005), .Y(n29000)
         );
  AOI22X1 U17138 ( .A(reg_file[550]), .B(n25278), .C(reg_file[678]), .D(n25289), .Y(n28998) );
  AOI22X1 U17139 ( .A(reg_file[806]), .B(n25299), .C(reg_file[934]), .D(n25310), .Y(n28997) );
  NOR2X1 U17140 ( .A(n29006), .B(n29007), .Y(n28984) );
  NAND3X1 U17141 ( .A(n29008), .B(n29009), .C(n29010), .Y(n29007) );
  NOR2X1 U17142 ( .A(n29011), .B(n29012), .Y(n29010) );
  OAI22X1 U17143 ( .A(n25320), .B(n29013), .C(n25330), .D(n29014), .Y(n29012)
         );
  OAI22X1 U17144 ( .A(n25341), .B(n29015), .C(n25351), .D(n29016), .Y(n29011)
         );
  AOI22X1 U17145 ( .A(reg_file[3494]), .B(n25362), .C(reg_file[3366]), .D(
        n25373), .Y(n29009) );
  AOI22X1 U17146 ( .A(reg_file[3238]), .B(n25383), .C(reg_file[3110]), .D(
        n25394), .Y(n29008) );
  NAND3X1 U17147 ( .A(n29017), .B(n29018), .C(n29019), .Y(n29006) );
  NOR2X1 U17148 ( .A(n29020), .B(n29021), .Y(n29019) );
  OAI22X1 U17149 ( .A(n25404), .B(n29022), .C(n25414), .D(n29023), .Y(n29021)
         );
  OAI22X1 U17150 ( .A(n25425), .B(n29024), .C(n25435), .D(n29025), .Y(n29020)
         );
  AOI22X1 U17151 ( .A(reg_file[2470]), .B(n25446), .C(reg_file[2342]), .D(
        n25457), .Y(n29018) );
  AOI22X1 U17152 ( .A(reg_file[2214]), .B(n25467), .C(reg_file[2086]), .D(
        n25478), .Y(n29017) );
  AOI21X1 U17153 ( .A(n29026), .B(n29027), .C(n25141), .Y(rd2data1040_37_) );
  NOR2X1 U17154 ( .A(n29028), .B(n29029), .Y(n29027) );
  NAND3X1 U17155 ( .A(n29030), .B(n29031), .C(n29032), .Y(n29029) );
  NOR2X1 U17156 ( .A(n29033), .B(n29034), .Y(n29032) );
  OAI22X1 U17157 ( .A(n25152), .B(n29035), .C(n25162), .D(n29036), .Y(n29034)
         );
  OAI22X1 U17158 ( .A(n25173), .B(n29037), .C(n25183), .D(n29038), .Y(n29033)
         );
  AOI22X1 U17159 ( .A(reg_file[1445]), .B(n25194), .C(reg_file[1317]), .D(
        n25205), .Y(n29031) );
  AOI22X1 U17160 ( .A(reg_file[1189]), .B(n25215), .C(reg_file[1061]), .D(
        n25226), .Y(n29030) );
  NAND3X1 U17161 ( .A(n29039), .B(n29040), .C(n29041), .Y(n29028) );
  NOR2X1 U17162 ( .A(n29042), .B(n29043), .Y(n29041) );
  OAI22X1 U17163 ( .A(n25236), .B(n29044), .C(n25246), .D(n29045), .Y(n29043)
         );
  OAI22X1 U17164 ( .A(n25257), .B(n29046), .C(n25267), .D(n29047), .Y(n29042)
         );
  AOI22X1 U17165 ( .A(reg_file[549]), .B(n25278), .C(reg_file[677]), .D(n25289), .Y(n29040) );
  AOI22X1 U17166 ( .A(reg_file[805]), .B(n25299), .C(reg_file[933]), .D(n25310), .Y(n29039) );
  NOR2X1 U17167 ( .A(n29048), .B(n29049), .Y(n29026) );
  NAND3X1 U17168 ( .A(n29050), .B(n29051), .C(n29052), .Y(n29049) );
  NOR2X1 U17169 ( .A(n29053), .B(n29054), .Y(n29052) );
  OAI22X1 U17170 ( .A(n25320), .B(n29055), .C(n25330), .D(n29056), .Y(n29054)
         );
  OAI22X1 U17171 ( .A(n25341), .B(n29057), .C(n25351), .D(n29058), .Y(n29053)
         );
  AOI22X1 U17172 ( .A(reg_file[3493]), .B(n25362), .C(reg_file[3365]), .D(
        n25373), .Y(n29051) );
  AOI22X1 U17173 ( .A(reg_file[3237]), .B(n25383), .C(reg_file[3109]), .D(
        n25394), .Y(n29050) );
  NAND3X1 U17174 ( .A(n29059), .B(n29060), .C(n29061), .Y(n29048) );
  NOR2X1 U17175 ( .A(n29062), .B(n29063), .Y(n29061) );
  OAI22X1 U17176 ( .A(n25404), .B(n29064), .C(n25414), .D(n29065), .Y(n29063)
         );
  OAI22X1 U17177 ( .A(n25425), .B(n29066), .C(n25435), .D(n29067), .Y(n29062)
         );
  AOI22X1 U17178 ( .A(reg_file[2469]), .B(n25446), .C(reg_file[2341]), .D(
        n25457), .Y(n29060) );
  AOI22X1 U17179 ( .A(reg_file[2213]), .B(n25467), .C(reg_file[2085]), .D(
        n25478), .Y(n29059) );
  AOI21X1 U17180 ( .A(n29068), .B(n29069), .C(n25141), .Y(rd2data1040_36_) );
  NOR2X1 U17181 ( .A(n29070), .B(n29071), .Y(n29069) );
  NAND3X1 U17182 ( .A(n29072), .B(n29073), .C(n29074), .Y(n29071) );
  NOR2X1 U17183 ( .A(n29075), .B(n29076), .Y(n29074) );
  OAI22X1 U17184 ( .A(n25152), .B(n29077), .C(n25162), .D(n29078), .Y(n29076)
         );
  OAI22X1 U17185 ( .A(n25173), .B(n29079), .C(n25183), .D(n29080), .Y(n29075)
         );
  AOI22X1 U17186 ( .A(reg_file[1444]), .B(n25194), .C(reg_file[1316]), .D(
        n25205), .Y(n29073) );
  AOI22X1 U17187 ( .A(reg_file[1188]), .B(n25215), .C(reg_file[1060]), .D(
        n25226), .Y(n29072) );
  NAND3X1 U17188 ( .A(n29081), .B(n29082), .C(n29083), .Y(n29070) );
  NOR2X1 U17189 ( .A(n29084), .B(n29085), .Y(n29083) );
  OAI22X1 U17190 ( .A(n25236), .B(n29086), .C(n25246), .D(n29087), .Y(n29085)
         );
  OAI22X1 U17191 ( .A(n25257), .B(n29088), .C(n25267), .D(n29089), .Y(n29084)
         );
  AOI22X1 U17192 ( .A(reg_file[548]), .B(n25278), .C(reg_file[676]), .D(n25289), .Y(n29082) );
  AOI22X1 U17193 ( .A(reg_file[804]), .B(n25299), .C(reg_file[932]), .D(n25310), .Y(n29081) );
  NOR2X1 U17194 ( .A(n29090), .B(n29091), .Y(n29068) );
  NAND3X1 U17195 ( .A(n29092), .B(n29093), .C(n29094), .Y(n29091) );
  NOR2X1 U17196 ( .A(n29095), .B(n29096), .Y(n29094) );
  OAI22X1 U17197 ( .A(n25320), .B(n29097), .C(n25330), .D(n29098), .Y(n29096)
         );
  OAI22X1 U17198 ( .A(n25341), .B(n29099), .C(n25351), .D(n29100), .Y(n29095)
         );
  AOI22X1 U17199 ( .A(reg_file[3492]), .B(n25362), .C(reg_file[3364]), .D(
        n25373), .Y(n29093) );
  AOI22X1 U17200 ( .A(reg_file[3236]), .B(n25383), .C(reg_file[3108]), .D(
        n25394), .Y(n29092) );
  NAND3X1 U17201 ( .A(n29101), .B(n29102), .C(n29103), .Y(n29090) );
  NOR2X1 U17202 ( .A(n29104), .B(n29105), .Y(n29103) );
  OAI22X1 U17203 ( .A(n25404), .B(n29106), .C(n25414), .D(n29107), .Y(n29105)
         );
  OAI22X1 U17204 ( .A(n25425), .B(n29108), .C(n25435), .D(n29109), .Y(n29104)
         );
  AOI22X1 U17205 ( .A(reg_file[2468]), .B(n25446), .C(reg_file[2340]), .D(
        n25457), .Y(n29102) );
  AOI22X1 U17206 ( .A(reg_file[2212]), .B(n25467), .C(reg_file[2084]), .D(
        n25478), .Y(n29101) );
  AOI21X1 U17207 ( .A(n29110), .B(n29111), .C(n25141), .Y(rd2data1040_35_) );
  NOR2X1 U17208 ( .A(n29112), .B(n29113), .Y(n29111) );
  NAND3X1 U17209 ( .A(n29114), .B(n29115), .C(n29116), .Y(n29113) );
  NOR2X1 U17210 ( .A(n29117), .B(n29118), .Y(n29116) );
  OAI22X1 U17211 ( .A(n25152), .B(n29119), .C(n25162), .D(n29120), .Y(n29118)
         );
  OAI22X1 U17212 ( .A(n25173), .B(n29121), .C(n25183), .D(n29122), .Y(n29117)
         );
  AOI22X1 U17213 ( .A(reg_file[1443]), .B(n25194), .C(reg_file[1315]), .D(
        n25205), .Y(n29115) );
  AOI22X1 U17214 ( .A(reg_file[1187]), .B(n25215), .C(reg_file[1059]), .D(
        n25226), .Y(n29114) );
  NAND3X1 U17215 ( .A(n29123), .B(n29124), .C(n29125), .Y(n29112) );
  NOR2X1 U17216 ( .A(n29126), .B(n29127), .Y(n29125) );
  OAI22X1 U17217 ( .A(n25236), .B(n29128), .C(n25246), .D(n29129), .Y(n29127)
         );
  OAI22X1 U17218 ( .A(n25257), .B(n29130), .C(n25267), .D(n29131), .Y(n29126)
         );
  AOI22X1 U17219 ( .A(reg_file[547]), .B(n25278), .C(reg_file[675]), .D(n25289), .Y(n29124) );
  AOI22X1 U17220 ( .A(reg_file[803]), .B(n25299), .C(reg_file[931]), .D(n25310), .Y(n29123) );
  NOR2X1 U17221 ( .A(n29132), .B(n29133), .Y(n29110) );
  NAND3X1 U17222 ( .A(n29134), .B(n29135), .C(n29136), .Y(n29133) );
  NOR2X1 U17223 ( .A(n29137), .B(n29138), .Y(n29136) );
  OAI22X1 U17224 ( .A(n25320), .B(n29139), .C(n25330), .D(n29140), .Y(n29138)
         );
  OAI22X1 U17225 ( .A(n25341), .B(n29141), .C(n25351), .D(n29142), .Y(n29137)
         );
  AOI22X1 U17226 ( .A(reg_file[3491]), .B(n25362), .C(reg_file[3363]), .D(
        n25373), .Y(n29135) );
  AOI22X1 U17227 ( .A(reg_file[3235]), .B(n25383), .C(reg_file[3107]), .D(
        n25394), .Y(n29134) );
  NAND3X1 U17228 ( .A(n29143), .B(n29144), .C(n29145), .Y(n29132) );
  NOR2X1 U17229 ( .A(n29146), .B(n29147), .Y(n29145) );
  OAI22X1 U17230 ( .A(n25404), .B(n29148), .C(n25414), .D(n29149), .Y(n29147)
         );
  OAI22X1 U17231 ( .A(n25425), .B(n29150), .C(n25435), .D(n29151), .Y(n29146)
         );
  AOI22X1 U17232 ( .A(reg_file[2467]), .B(n25446), .C(reg_file[2339]), .D(
        n25457), .Y(n29144) );
  AOI22X1 U17233 ( .A(reg_file[2211]), .B(n25467), .C(reg_file[2083]), .D(
        n25478), .Y(n29143) );
  AOI21X1 U17234 ( .A(n29152), .B(n29153), .C(n25141), .Y(rd2data1040_34_) );
  NOR2X1 U17235 ( .A(n29154), .B(n29155), .Y(n29153) );
  NAND3X1 U17236 ( .A(n29156), .B(n29157), .C(n29158), .Y(n29155) );
  NOR2X1 U17237 ( .A(n29159), .B(n29160), .Y(n29158) );
  OAI22X1 U17238 ( .A(n25152), .B(n29161), .C(n25162), .D(n29162), .Y(n29160)
         );
  OAI22X1 U17239 ( .A(n25173), .B(n29163), .C(n25183), .D(n29164), .Y(n29159)
         );
  AOI22X1 U17240 ( .A(reg_file[1442]), .B(n25194), .C(reg_file[1314]), .D(
        n25205), .Y(n29157) );
  AOI22X1 U17241 ( .A(reg_file[1186]), .B(n25215), .C(reg_file[1058]), .D(
        n25226), .Y(n29156) );
  NAND3X1 U17242 ( .A(n29165), .B(n29166), .C(n29167), .Y(n29154) );
  NOR2X1 U17243 ( .A(n29168), .B(n29169), .Y(n29167) );
  OAI22X1 U17244 ( .A(n25236), .B(n29170), .C(n25246), .D(n29171), .Y(n29169)
         );
  OAI22X1 U17245 ( .A(n25257), .B(n29172), .C(n25267), .D(n29173), .Y(n29168)
         );
  AOI22X1 U17246 ( .A(reg_file[546]), .B(n25278), .C(reg_file[674]), .D(n25289), .Y(n29166) );
  AOI22X1 U17247 ( .A(reg_file[802]), .B(n25299), .C(reg_file[930]), .D(n25310), .Y(n29165) );
  NOR2X1 U17248 ( .A(n29174), .B(n29175), .Y(n29152) );
  NAND3X1 U17249 ( .A(n29176), .B(n29177), .C(n29178), .Y(n29175) );
  NOR2X1 U17250 ( .A(n29179), .B(n29180), .Y(n29178) );
  OAI22X1 U17251 ( .A(n25320), .B(n29181), .C(n25330), .D(n29182), .Y(n29180)
         );
  OAI22X1 U17252 ( .A(n25341), .B(n29183), .C(n25351), .D(n29184), .Y(n29179)
         );
  AOI22X1 U17253 ( .A(reg_file[3490]), .B(n25362), .C(reg_file[3362]), .D(
        n25373), .Y(n29177) );
  AOI22X1 U17254 ( .A(reg_file[3234]), .B(n25383), .C(reg_file[3106]), .D(
        n25394), .Y(n29176) );
  NAND3X1 U17255 ( .A(n29185), .B(n29186), .C(n29187), .Y(n29174) );
  NOR2X1 U17256 ( .A(n29188), .B(n29189), .Y(n29187) );
  OAI22X1 U17257 ( .A(n25404), .B(n29190), .C(n25414), .D(n29191), .Y(n29189)
         );
  OAI22X1 U17258 ( .A(n25425), .B(n29192), .C(n25435), .D(n29193), .Y(n29188)
         );
  AOI22X1 U17259 ( .A(reg_file[2466]), .B(n25446), .C(reg_file[2338]), .D(
        n25457), .Y(n29186) );
  AOI22X1 U17260 ( .A(reg_file[2210]), .B(n25467), .C(reg_file[2082]), .D(
        n25478), .Y(n29185) );
  AOI21X1 U17261 ( .A(n29194), .B(n29195), .C(n25141), .Y(rd2data1040_33_) );
  NOR2X1 U17262 ( .A(n29196), .B(n29197), .Y(n29195) );
  NAND3X1 U17263 ( .A(n29198), .B(n29199), .C(n29200), .Y(n29197) );
  NOR2X1 U17264 ( .A(n29201), .B(n29202), .Y(n29200) );
  OAI22X1 U17265 ( .A(n25152), .B(n29203), .C(n25162), .D(n29204), .Y(n29202)
         );
  OAI22X1 U17266 ( .A(n25173), .B(n29205), .C(n25183), .D(n29206), .Y(n29201)
         );
  AOI22X1 U17267 ( .A(reg_file[1441]), .B(n25194), .C(reg_file[1313]), .D(
        n25205), .Y(n29199) );
  AOI22X1 U17268 ( .A(reg_file[1185]), .B(n25215), .C(reg_file[1057]), .D(
        n25226), .Y(n29198) );
  NAND3X1 U17269 ( .A(n29207), .B(n29208), .C(n29209), .Y(n29196) );
  NOR2X1 U17270 ( .A(n29210), .B(n29211), .Y(n29209) );
  OAI22X1 U17271 ( .A(n25236), .B(n29212), .C(n25246), .D(n29213), .Y(n29211)
         );
  OAI22X1 U17272 ( .A(n25257), .B(n29214), .C(n25267), .D(n29215), .Y(n29210)
         );
  AOI22X1 U17273 ( .A(reg_file[545]), .B(n25278), .C(reg_file[673]), .D(n25289), .Y(n29208) );
  AOI22X1 U17274 ( .A(reg_file[801]), .B(n25299), .C(reg_file[929]), .D(n25310), .Y(n29207) );
  NOR2X1 U17275 ( .A(n29216), .B(n29217), .Y(n29194) );
  NAND3X1 U17276 ( .A(n29218), .B(n29219), .C(n29220), .Y(n29217) );
  NOR2X1 U17277 ( .A(n29221), .B(n29222), .Y(n29220) );
  OAI22X1 U17278 ( .A(n25320), .B(n29223), .C(n25330), .D(n29224), .Y(n29222)
         );
  OAI22X1 U17279 ( .A(n25341), .B(n29225), .C(n25351), .D(n29226), .Y(n29221)
         );
  AOI22X1 U17280 ( .A(reg_file[3489]), .B(n25362), .C(reg_file[3361]), .D(
        n25373), .Y(n29219) );
  AOI22X1 U17281 ( .A(reg_file[3233]), .B(n25383), .C(reg_file[3105]), .D(
        n25394), .Y(n29218) );
  NAND3X1 U17282 ( .A(n29227), .B(n29228), .C(n29229), .Y(n29216) );
  NOR2X1 U17283 ( .A(n29230), .B(n29231), .Y(n29229) );
  OAI22X1 U17284 ( .A(n25404), .B(n29232), .C(n25414), .D(n29233), .Y(n29231)
         );
  OAI22X1 U17285 ( .A(n25425), .B(n29234), .C(n25435), .D(n29235), .Y(n29230)
         );
  AOI22X1 U17286 ( .A(reg_file[2465]), .B(n25446), .C(reg_file[2337]), .D(
        n25457), .Y(n29228) );
  AOI22X1 U17287 ( .A(reg_file[2209]), .B(n25467), .C(reg_file[2081]), .D(
        n25478), .Y(n29227) );
  AOI21X1 U17288 ( .A(n29236), .B(n29237), .C(n25141), .Y(rd2data1040_32_) );
  NOR2X1 U17289 ( .A(n29238), .B(n29239), .Y(n29237) );
  NAND3X1 U17290 ( .A(n29240), .B(n29241), .C(n29242), .Y(n29239) );
  NOR2X1 U17291 ( .A(n29243), .B(n29244), .Y(n29242) );
  OAI22X1 U17292 ( .A(n25152), .B(n29245), .C(n25162), .D(n29246), .Y(n29244)
         );
  OAI22X1 U17293 ( .A(n25173), .B(n29247), .C(n25183), .D(n29248), .Y(n29243)
         );
  AOI22X1 U17294 ( .A(reg_file[1440]), .B(n25194), .C(reg_file[1312]), .D(
        n25205), .Y(n29241) );
  AOI22X1 U17295 ( .A(reg_file[1184]), .B(n25215), .C(reg_file[1056]), .D(
        n25226), .Y(n29240) );
  NAND3X1 U17296 ( .A(n29249), .B(n29250), .C(n29251), .Y(n29238) );
  NOR2X1 U17297 ( .A(n29252), .B(n29253), .Y(n29251) );
  OAI22X1 U17298 ( .A(n25236), .B(n29254), .C(n25246), .D(n29255), .Y(n29253)
         );
  OAI22X1 U17299 ( .A(n25257), .B(n29256), .C(n25267), .D(n29257), .Y(n29252)
         );
  AOI22X1 U17300 ( .A(reg_file[544]), .B(n25278), .C(reg_file[672]), .D(n25289), .Y(n29250) );
  AOI22X1 U17301 ( .A(reg_file[800]), .B(n25299), .C(reg_file[928]), .D(n25310), .Y(n29249) );
  NOR2X1 U17302 ( .A(n29258), .B(n29259), .Y(n29236) );
  NAND3X1 U17303 ( .A(n29260), .B(n29261), .C(n29262), .Y(n29259) );
  NOR2X1 U17304 ( .A(n29263), .B(n29264), .Y(n29262) );
  OAI22X1 U17305 ( .A(n25320), .B(n29265), .C(n25330), .D(n29266), .Y(n29264)
         );
  OAI22X1 U17306 ( .A(n25341), .B(n29267), .C(n25351), .D(n29268), .Y(n29263)
         );
  AOI22X1 U17307 ( .A(reg_file[3488]), .B(n25362), .C(reg_file[3360]), .D(
        n25373), .Y(n29261) );
  AOI22X1 U17308 ( .A(reg_file[3232]), .B(n25383), .C(reg_file[3104]), .D(
        n25394), .Y(n29260) );
  NAND3X1 U17309 ( .A(n29269), .B(n29270), .C(n29271), .Y(n29258) );
  NOR2X1 U17310 ( .A(n29272), .B(n29273), .Y(n29271) );
  OAI22X1 U17311 ( .A(n25404), .B(n29274), .C(n25414), .D(n29275), .Y(n29273)
         );
  OAI22X1 U17312 ( .A(n25425), .B(n29276), .C(n25435), .D(n29277), .Y(n29272)
         );
  AOI22X1 U17313 ( .A(reg_file[2464]), .B(n25446), .C(reg_file[2336]), .D(
        n25457), .Y(n29270) );
  AOI22X1 U17314 ( .A(reg_file[2208]), .B(n25467), .C(reg_file[2080]), .D(
        n25478), .Y(n29269) );
  AOI21X1 U17315 ( .A(n29278), .B(n29279), .C(n25141), .Y(rd2data1040_31_) );
  NOR2X1 U17316 ( .A(n29280), .B(n29281), .Y(n29279) );
  NAND3X1 U17317 ( .A(n29282), .B(n29283), .C(n29284), .Y(n29281) );
  NOR2X1 U17318 ( .A(n29285), .B(n29286), .Y(n29284) );
  OAI22X1 U17319 ( .A(n25152), .B(n29287), .C(n25162), .D(n29288), .Y(n29286)
         );
  OAI22X1 U17320 ( .A(n25173), .B(n29289), .C(n25183), .D(n29290), .Y(n29285)
         );
  AOI22X1 U17321 ( .A(reg_file[1439]), .B(n25194), .C(reg_file[1311]), .D(
        n25205), .Y(n29283) );
  AOI22X1 U17322 ( .A(reg_file[1183]), .B(n25215), .C(reg_file[1055]), .D(
        n25226), .Y(n29282) );
  NAND3X1 U17323 ( .A(n29291), .B(n29292), .C(n29293), .Y(n29280) );
  NOR2X1 U17324 ( .A(n29294), .B(n29295), .Y(n29293) );
  OAI22X1 U17325 ( .A(n25236), .B(n29296), .C(n25246), .D(n29297), .Y(n29295)
         );
  OAI22X1 U17326 ( .A(n25257), .B(n29298), .C(n25267), .D(n29299), .Y(n29294)
         );
  AOI22X1 U17327 ( .A(reg_file[543]), .B(n25278), .C(reg_file[671]), .D(n25289), .Y(n29292) );
  AOI22X1 U17328 ( .A(reg_file[799]), .B(n25299), .C(reg_file[927]), .D(n25310), .Y(n29291) );
  NOR2X1 U17329 ( .A(n29300), .B(n29301), .Y(n29278) );
  NAND3X1 U17330 ( .A(n29302), .B(n29303), .C(n29304), .Y(n29301) );
  NOR2X1 U17331 ( .A(n29305), .B(n29306), .Y(n29304) );
  OAI22X1 U17332 ( .A(n25320), .B(n29307), .C(n25330), .D(n29308), .Y(n29306)
         );
  OAI22X1 U17333 ( .A(n25341), .B(n29309), .C(n25351), .D(n29310), .Y(n29305)
         );
  AOI22X1 U17334 ( .A(reg_file[3487]), .B(n25362), .C(reg_file[3359]), .D(
        n25373), .Y(n29303) );
  AOI22X1 U17335 ( .A(reg_file[3231]), .B(n25383), .C(reg_file[3103]), .D(
        n25394), .Y(n29302) );
  NAND3X1 U17336 ( .A(n29311), .B(n29312), .C(n29313), .Y(n29300) );
  NOR2X1 U17337 ( .A(n29314), .B(n29315), .Y(n29313) );
  OAI22X1 U17338 ( .A(n25404), .B(n29316), .C(n25414), .D(n29317), .Y(n29315)
         );
  OAI22X1 U17339 ( .A(n25425), .B(n29318), .C(n25435), .D(n29319), .Y(n29314)
         );
  AOI22X1 U17340 ( .A(reg_file[2463]), .B(n25446), .C(reg_file[2335]), .D(
        n25457), .Y(n29312) );
  AOI22X1 U17341 ( .A(reg_file[2207]), .B(n25467), .C(reg_file[2079]), .D(
        n25478), .Y(n29311) );
  AOI21X1 U17342 ( .A(n29320), .B(n29321), .C(n25141), .Y(rd2data1040_30_) );
  NOR2X1 U17343 ( .A(n29322), .B(n29323), .Y(n29321) );
  NAND3X1 U17344 ( .A(n29324), .B(n29325), .C(n29326), .Y(n29323) );
  NOR2X1 U17345 ( .A(n29327), .B(n29328), .Y(n29326) );
  OAI22X1 U17346 ( .A(n25151), .B(n29329), .C(n25162), .D(n29330), .Y(n29328)
         );
  OAI22X1 U17347 ( .A(n25172), .B(n29331), .C(n25183), .D(n29332), .Y(n29327)
         );
  AOI22X1 U17348 ( .A(reg_file[1438]), .B(n25194), .C(reg_file[1310]), .D(
        n25204), .Y(n29325) );
  AOI22X1 U17349 ( .A(reg_file[1182]), .B(n25215), .C(reg_file[1054]), .D(
        n25225), .Y(n29324) );
  NAND3X1 U17350 ( .A(n29333), .B(n29334), .C(n29335), .Y(n29322) );
  NOR2X1 U17351 ( .A(n29336), .B(n29337), .Y(n29335) );
  OAI22X1 U17352 ( .A(n25235), .B(n29338), .C(n25246), .D(n29339), .Y(n29337)
         );
  OAI22X1 U17353 ( .A(n25256), .B(n29340), .C(n25267), .D(n29341), .Y(n29336)
         );
  AOI22X1 U17354 ( .A(reg_file[542]), .B(n25278), .C(reg_file[670]), .D(n25288), .Y(n29334) );
  AOI22X1 U17355 ( .A(reg_file[798]), .B(n25299), .C(reg_file[926]), .D(n25309), .Y(n29333) );
  NOR2X1 U17356 ( .A(n29342), .B(n29343), .Y(n29320) );
  NAND3X1 U17357 ( .A(n29344), .B(n29345), .C(n29346), .Y(n29343) );
  NOR2X1 U17358 ( .A(n29347), .B(n29348), .Y(n29346) );
  OAI22X1 U17359 ( .A(n25319), .B(n29349), .C(n25330), .D(n29350), .Y(n29348)
         );
  OAI22X1 U17360 ( .A(n25340), .B(n29351), .C(n25351), .D(n29352), .Y(n29347)
         );
  AOI22X1 U17361 ( .A(reg_file[3486]), .B(n25362), .C(reg_file[3358]), .D(
        n25372), .Y(n29345) );
  AOI22X1 U17362 ( .A(reg_file[3230]), .B(n25383), .C(reg_file[3102]), .D(
        n25393), .Y(n29344) );
  NAND3X1 U17363 ( .A(n29353), .B(n29354), .C(n29355), .Y(n29342) );
  NOR2X1 U17364 ( .A(n29356), .B(n29357), .Y(n29355) );
  OAI22X1 U17365 ( .A(n25403), .B(n29358), .C(n25414), .D(n29359), .Y(n29357)
         );
  OAI22X1 U17366 ( .A(n25424), .B(n29360), .C(n25435), .D(n29361), .Y(n29356)
         );
  AOI22X1 U17367 ( .A(reg_file[2462]), .B(n25446), .C(reg_file[2334]), .D(
        n25456), .Y(n29354) );
  AOI22X1 U17368 ( .A(reg_file[2206]), .B(n25467), .C(reg_file[2078]), .D(
        n25477), .Y(n29353) );
  AOI21X1 U17369 ( .A(n29362), .B(n29363), .C(n25141), .Y(rd2data1040_2_) );
  NOR2X1 U17370 ( .A(n29364), .B(n29365), .Y(n29363) );
  NAND3X1 U17371 ( .A(n29366), .B(n29367), .C(n29368), .Y(n29365) );
  NOR2X1 U17372 ( .A(n29369), .B(n29370), .Y(n29368) );
  OAI22X1 U17373 ( .A(n25151), .B(n29371), .C(n25162), .D(n29372), .Y(n29370)
         );
  OAI22X1 U17374 ( .A(n25172), .B(n29373), .C(n25183), .D(n29374), .Y(n29369)
         );
  AOI22X1 U17375 ( .A(reg_file[1410]), .B(n25194), .C(reg_file[1282]), .D(
        n25204), .Y(n29367) );
  AOI22X1 U17376 ( .A(reg_file[1154]), .B(n25215), .C(reg_file[1026]), .D(
        n25225), .Y(n29366) );
  NAND3X1 U17377 ( .A(n29375), .B(n29376), .C(n29377), .Y(n29364) );
  NOR2X1 U17378 ( .A(n29378), .B(n29379), .Y(n29377) );
  OAI22X1 U17379 ( .A(n25235), .B(n29380), .C(n25246), .D(n29381), .Y(n29379)
         );
  OAI22X1 U17380 ( .A(n25256), .B(n29382), .C(n25267), .D(n29383), .Y(n29378)
         );
  AOI22X1 U17381 ( .A(reg_file[514]), .B(n25278), .C(reg_file[642]), .D(n25288), .Y(n29376) );
  AOI22X1 U17382 ( .A(reg_file[770]), .B(n25299), .C(reg_file[898]), .D(n25309), .Y(n29375) );
  NOR2X1 U17383 ( .A(n29384), .B(n29385), .Y(n29362) );
  NAND3X1 U17384 ( .A(n29386), .B(n29387), .C(n29388), .Y(n29385) );
  NOR2X1 U17385 ( .A(n29389), .B(n29390), .Y(n29388) );
  OAI22X1 U17386 ( .A(n25319), .B(n29391), .C(n25330), .D(n29392), .Y(n29390)
         );
  OAI22X1 U17387 ( .A(n25340), .B(n29393), .C(n25351), .D(n29394), .Y(n29389)
         );
  AOI22X1 U17388 ( .A(reg_file[3458]), .B(n25362), .C(reg_file[3330]), .D(
        n25372), .Y(n29387) );
  AOI22X1 U17389 ( .A(reg_file[3202]), .B(n25383), .C(reg_file[3074]), .D(
        n25393), .Y(n29386) );
  NAND3X1 U17390 ( .A(n29395), .B(n29396), .C(n29397), .Y(n29384) );
  NOR2X1 U17391 ( .A(n29398), .B(n29399), .Y(n29397) );
  OAI22X1 U17392 ( .A(n25403), .B(n29400), .C(n25414), .D(n29401), .Y(n29399)
         );
  OAI22X1 U17393 ( .A(n25424), .B(n29402), .C(n25435), .D(n29403), .Y(n29398)
         );
  AOI22X1 U17394 ( .A(reg_file[2434]), .B(n25446), .C(reg_file[2306]), .D(
        n25456), .Y(n29396) );
  AOI22X1 U17395 ( .A(reg_file[2178]), .B(n25467), .C(reg_file[2050]), .D(
        n25477), .Y(n29395) );
  AOI21X1 U17396 ( .A(n29404), .B(n29405), .C(n25141), .Y(rd2data1040_29_) );
  NOR2X1 U17397 ( .A(n29406), .B(n29407), .Y(n29405) );
  NAND3X1 U17398 ( .A(n29408), .B(n29409), .C(n29410), .Y(n29407) );
  NOR2X1 U17399 ( .A(n29411), .B(n29412), .Y(n29410) );
  OAI22X1 U17400 ( .A(n25151), .B(n29413), .C(n25162), .D(n29414), .Y(n29412)
         );
  OAI22X1 U17401 ( .A(n25172), .B(n29415), .C(n25183), .D(n29416), .Y(n29411)
         );
  AOI22X1 U17402 ( .A(reg_file[1437]), .B(n25194), .C(reg_file[1309]), .D(
        n25204), .Y(n29409) );
  AOI22X1 U17403 ( .A(reg_file[1181]), .B(n25215), .C(reg_file[1053]), .D(
        n25225), .Y(n29408) );
  NAND3X1 U17404 ( .A(n29417), .B(n29418), .C(n29419), .Y(n29406) );
  NOR2X1 U17405 ( .A(n29420), .B(n29421), .Y(n29419) );
  OAI22X1 U17406 ( .A(n25235), .B(n29422), .C(n25246), .D(n29423), .Y(n29421)
         );
  OAI22X1 U17407 ( .A(n25256), .B(n29424), .C(n25267), .D(n29425), .Y(n29420)
         );
  AOI22X1 U17408 ( .A(reg_file[541]), .B(n25278), .C(reg_file[669]), .D(n25288), .Y(n29418) );
  AOI22X1 U17409 ( .A(reg_file[797]), .B(n25299), .C(reg_file[925]), .D(n25309), .Y(n29417) );
  NOR2X1 U17410 ( .A(n29426), .B(n29427), .Y(n29404) );
  NAND3X1 U17411 ( .A(n29428), .B(n29429), .C(n29430), .Y(n29427) );
  NOR2X1 U17412 ( .A(n29431), .B(n29432), .Y(n29430) );
  OAI22X1 U17413 ( .A(n25319), .B(n29433), .C(n25330), .D(n29434), .Y(n29432)
         );
  OAI22X1 U17414 ( .A(n25340), .B(n29435), .C(n25351), .D(n29436), .Y(n29431)
         );
  AOI22X1 U17415 ( .A(reg_file[3485]), .B(n25362), .C(reg_file[3357]), .D(
        n25372), .Y(n29429) );
  AOI22X1 U17416 ( .A(reg_file[3229]), .B(n25383), .C(reg_file[3101]), .D(
        n25393), .Y(n29428) );
  NAND3X1 U17417 ( .A(n29437), .B(n29438), .C(n29439), .Y(n29426) );
  NOR2X1 U17418 ( .A(n29440), .B(n29441), .Y(n29439) );
  OAI22X1 U17419 ( .A(n25403), .B(n29442), .C(n25414), .D(n29443), .Y(n29441)
         );
  OAI22X1 U17420 ( .A(n25424), .B(n29444), .C(n25435), .D(n29445), .Y(n29440)
         );
  AOI22X1 U17421 ( .A(reg_file[2461]), .B(n25446), .C(reg_file[2333]), .D(
        n25456), .Y(n29438) );
  AOI22X1 U17422 ( .A(reg_file[2205]), .B(n25467), .C(reg_file[2077]), .D(
        n25477), .Y(n29437) );
  AOI21X1 U17423 ( .A(n29446), .B(n29447), .C(n25141), .Y(rd2data1040_28_) );
  NOR2X1 U17424 ( .A(n29448), .B(n29449), .Y(n29447) );
  NAND3X1 U17425 ( .A(n29450), .B(n29451), .C(n29452), .Y(n29449) );
  NOR2X1 U17426 ( .A(n29453), .B(n29454), .Y(n29452) );
  OAI22X1 U17427 ( .A(n25151), .B(n29455), .C(n25162), .D(n29456), .Y(n29454)
         );
  OAI22X1 U17428 ( .A(n25172), .B(n29457), .C(n25183), .D(n29458), .Y(n29453)
         );
  AOI22X1 U17429 ( .A(reg_file[1436]), .B(n25194), .C(reg_file[1308]), .D(
        n25204), .Y(n29451) );
  AOI22X1 U17430 ( .A(reg_file[1180]), .B(n25215), .C(reg_file[1052]), .D(
        n25225), .Y(n29450) );
  NAND3X1 U17431 ( .A(n29459), .B(n29460), .C(n29461), .Y(n29448) );
  NOR2X1 U17432 ( .A(n29462), .B(n29463), .Y(n29461) );
  OAI22X1 U17433 ( .A(n25235), .B(n29464), .C(n25246), .D(n29465), .Y(n29463)
         );
  OAI22X1 U17434 ( .A(n25256), .B(n29466), .C(n25267), .D(n29467), .Y(n29462)
         );
  AOI22X1 U17435 ( .A(reg_file[540]), .B(n25278), .C(reg_file[668]), .D(n25288), .Y(n29460) );
  AOI22X1 U17436 ( .A(reg_file[796]), .B(n25299), .C(reg_file[924]), .D(n25309), .Y(n29459) );
  NOR2X1 U17437 ( .A(n29468), .B(n29469), .Y(n29446) );
  NAND3X1 U17438 ( .A(n29470), .B(n29471), .C(n29472), .Y(n29469) );
  NOR2X1 U17439 ( .A(n29473), .B(n29474), .Y(n29472) );
  OAI22X1 U17440 ( .A(n25319), .B(n29475), .C(n25330), .D(n29476), .Y(n29474)
         );
  OAI22X1 U17441 ( .A(n25340), .B(n29477), .C(n25351), .D(n29478), .Y(n29473)
         );
  AOI22X1 U17442 ( .A(reg_file[3484]), .B(n25362), .C(reg_file[3356]), .D(
        n25372), .Y(n29471) );
  AOI22X1 U17443 ( .A(reg_file[3228]), .B(n25383), .C(reg_file[3100]), .D(
        n25393), .Y(n29470) );
  NAND3X1 U17444 ( .A(n29479), .B(n29480), .C(n29481), .Y(n29468) );
  NOR2X1 U17445 ( .A(n29482), .B(n29483), .Y(n29481) );
  OAI22X1 U17446 ( .A(n25403), .B(n29484), .C(n25414), .D(n29485), .Y(n29483)
         );
  OAI22X1 U17447 ( .A(n25424), .B(n29486), .C(n25435), .D(n29487), .Y(n29482)
         );
  AOI22X1 U17448 ( .A(reg_file[2460]), .B(n25446), .C(reg_file[2332]), .D(
        n25456), .Y(n29480) );
  AOI22X1 U17449 ( .A(reg_file[2204]), .B(n25467), .C(reg_file[2076]), .D(
        n25477), .Y(n29479) );
  AOI21X1 U17450 ( .A(n29488), .B(n29489), .C(n25140), .Y(rd2data1040_27_) );
  NOR2X1 U17451 ( .A(n29490), .B(n29491), .Y(n29489) );
  NAND3X1 U17452 ( .A(n29492), .B(n29493), .C(n29494), .Y(n29491) );
  NOR2X1 U17453 ( .A(n29495), .B(n29496), .Y(n29494) );
  OAI22X1 U17454 ( .A(n25151), .B(n29497), .C(n25161), .D(n29498), .Y(n29496)
         );
  OAI22X1 U17455 ( .A(n25172), .B(n29499), .C(n25182), .D(n29500), .Y(n29495)
         );
  AOI22X1 U17456 ( .A(reg_file[1435]), .B(n25193), .C(reg_file[1307]), .D(
        n25204), .Y(n29493) );
  AOI22X1 U17457 ( .A(reg_file[1179]), .B(n25214), .C(reg_file[1051]), .D(
        n25225), .Y(n29492) );
  NAND3X1 U17458 ( .A(n29501), .B(n29502), .C(n29503), .Y(n29490) );
  NOR2X1 U17459 ( .A(n29504), .B(n29505), .Y(n29503) );
  OAI22X1 U17460 ( .A(n25235), .B(n29506), .C(n25245), .D(n29507), .Y(n29505)
         );
  OAI22X1 U17461 ( .A(n25256), .B(n29508), .C(n25266), .D(n29509), .Y(n29504)
         );
  AOI22X1 U17462 ( .A(reg_file[539]), .B(n25277), .C(reg_file[667]), .D(n25288), .Y(n29502) );
  AOI22X1 U17463 ( .A(reg_file[795]), .B(n25298), .C(reg_file[923]), .D(n25309), .Y(n29501) );
  NOR2X1 U17464 ( .A(n29510), .B(n29511), .Y(n29488) );
  NAND3X1 U17465 ( .A(n29512), .B(n29513), .C(n29514), .Y(n29511) );
  NOR2X1 U17466 ( .A(n29515), .B(n29516), .Y(n29514) );
  OAI22X1 U17467 ( .A(n25319), .B(n29517), .C(n25329), .D(n29518), .Y(n29516)
         );
  OAI22X1 U17468 ( .A(n25340), .B(n29519), .C(n25350), .D(n29520), .Y(n29515)
         );
  AOI22X1 U17469 ( .A(reg_file[3483]), .B(n25361), .C(reg_file[3355]), .D(
        n25372), .Y(n29513) );
  AOI22X1 U17470 ( .A(reg_file[3227]), .B(n25382), .C(reg_file[3099]), .D(
        n25393), .Y(n29512) );
  NAND3X1 U17471 ( .A(n29521), .B(n29522), .C(n29523), .Y(n29510) );
  NOR2X1 U17472 ( .A(n29524), .B(n29525), .Y(n29523) );
  OAI22X1 U17473 ( .A(n25403), .B(n29526), .C(n25413), .D(n29527), .Y(n29525)
         );
  OAI22X1 U17474 ( .A(n25424), .B(n29528), .C(n25434), .D(n29529), .Y(n29524)
         );
  AOI22X1 U17475 ( .A(reg_file[2459]), .B(n25445), .C(reg_file[2331]), .D(
        n25456), .Y(n29522) );
  AOI22X1 U17476 ( .A(reg_file[2203]), .B(n25466), .C(reg_file[2075]), .D(
        n25477), .Y(n29521) );
  AOI21X1 U17477 ( .A(n29530), .B(n29531), .C(n25140), .Y(rd2data1040_26_) );
  NOR2X1 U17478 ( .A(n29532), .B(n29533), .Y(n29531) );
  NAND3X1 U17479 ( .A(n29534), .B(n29535), .C(n29536), .Y(n29533) );
  NOR2X1 U17480 ( .A(n29537), .B(n29538), .Y(n29536) );
  OAI22X1 U17481 ( .A(n25151), .B(n29539), .C(n25161), .D(n29540), .Y(n29538)
         );
  OAI22X1 U17482 ( .A(n25172), .B(n29541), .C(n25182), .D(n29542), .Y(n29537)
         );
  AOI22X1 U17483 ( .A(reg_file[1434]), .B(n25193), .C(reg_file[1306]), .D(
        n25204), .Y(n29535) );
  AOI22X1 U17484 ( .A(reg_file[1178]), .B(n25214), .C(reg_file[1050]), .D(
        n25225), .Y(n29534) );
  NAND3X1 U17485 ( .A(n29543), .B(n29544), .C(n29545), .Y(n29532) );
  NOR2X1 U17486 ( .A(n29546), .B(n29547), .Y(n29545) );
  OAI22X1 U17487 ( .A(n25235), .B(n29548), .C(n25245), .D(n29549), .Y(n29547)
         );
  OAI22X1 U17488 ( .A(n25256), .B(n29550), .C(n25266), .D(n29551), .Y(n29546)
         );
  AOI22X1 U17489 ( .A(reg_file[538]), .B(n25277), .C(reg_file[666]), .D(n25288), .Y(n29544) );
  AOI22X1 U17490 ( .A(reg_file[794]), .B(n25298), .C(reg_file[922]), .D(n25309), .Y(n29543) );
  NOR2X1 U17491 ( .A(n29552), .B(n29553), .Y(n29530) );
  NAND3X1 U17492 ( .A(n29554), .B(n29555), .C(n29556), .Y(n29553) );
  NOR2X1 U17493 ( .A(n29557), .B(n29558), .Y(n29556) );
  OAI22X1 U17494 ( .A(n25319), .B(n29559), .C(n25329), .D(n29560), .Y(n29558)
         );
  OAI22X1 U17495 ( .A(n25340), .B(n29561), .C(n25350), .D(n29562), .Y(n29557)
         );
  AOI22X1 U17496 ( .A(reg_file[3482]), .B(n25361), .C(reg_file[3354]), .D(
        n25372), .Y(n29555) );
  AOI22X1 U17497 ( .A(reg_file[3226]), .B(n25382), .C(reg_file[3098]), .D(
        n25393), .Y(n29554) );
  NAND3X1 U17498 ( .A(n29563), .B(n29564), .C(n29565), .Y(n29552) );
  NOR2X1 U17499 ( .A(n29566), .B(n29567), .Y(n29565) );
  OAI22X1 U17500 ( .A(n25403), .B(n29568), .C(n25413), .D(n29569), .Y(n29567)
         );
  OAI22X1 U17501 ( .A(n25424), .B(n29570), .C(n25434), .D(n29571), .Y(n29566)
         );
  AOI22X1 U17502 ( .A(reg_file[2458]), .B(n25445), .C(reg_file[2330]), .D(
        n25456), .Y(n29564) );
  AOI22X1 U17503 ( .A(reg_file[2202]), .B(n25466), .C(reg_file[2074]), .D(
        n25477), .Y(n29563) );
  AOI21X1 U17504 ( .A(n29572), .B(n29573), .C(n25140), .Y(rd2data1040_25_) );
  NOR2X1 U17505 ( .A(n29574), .B(n29575), .Y(n29573) );
  NAND3X1 U17506 ( .A(n29576), .B(n29577), .C(n29578), .Y(n29575) );
  NOR2X1 U17507 ( .A(n29579), .B(n29580), .Y(n29578) );
  OAI22X1 U17508 ( .A(n25151), .B(n29581), .C(n25161), .D(n29582), .Y(n29580)
         );
  OAI22X1 U17509 ( .A(n25172), .B(n29583), .C(n25182), .D(n29584), .Y(n29579)
         );
  AOI22X1 U17510 ( .A(reg_file[1433]), .B(n25193), .C(reg_file[1305]), .D(
        n25204), .Y(n29577) );
  AOI22X1 U17511 ( .A(reg_file[1177]), .B(n25214), .C(reg_file[1049]), .D(
        n25225), .Y(n29576) );
  NAND3X1 U17512 ( .A(n29585), .B(n29586), .C(n29587), .Y(n29574) );
  NOR2X1 U17513 ( .A(n29588), .B(n29589), .Y(n29587) );
  OAI22X1 U17514 ( .A(n25235), .B(n29590), .C(n25245), .D(n29591), .Y(n29589)
         );
  OAI22X1 U17515 ( .A(n25256), .B(n29592), .C(n25266), .D(n29593), .Y(n29588)
         );
  AOI22X1 U17516 ( .A(reg_file[537]), .B(n25277), .C(reg_file[665]), .D(n25288), .Y(n29586) );
  AOI22X1 U17517 ( .A(reg_file[793]), .B(n25298), .C(reg_file[921]), .D(n25309), .Y(n29585) );
  NOR2X1 U17518 ( .A(n29594), .B(n29595), .Y(n29572) );
  NAND3X1 U17519 ( .A(n29596), .B(n29597), .C(n29598), .Y(n29595) );
  NOR2X1 U17520 ( .A(n29599), .B(n29600), .Y(n29598) );
  OAI22X1 U17521 ( .A(n25319), .B(n29601), .C(n25329), .D(n29602), .Y(n29600)
         );
  OAI22X1 U17522 ( .A(n25340), .B(n29603), .C(n25350), .D(n29604), .Y(n29599)
         );
  AOI22X1 U17523 ( .A(reg_file[3481]), .B(n25361), .C(reg_file[3353]), .D(
        n25372), .Y(n29597) );
  AOI22X1 U17524 ( .A(reg_file[3225]), .B(n25382), .C(reg_file[3097]), .D(
        n25393), .Y(n29596) );
  NAND3X1 U17525 ( .A(n29605), .B(n29606), .C(n29607), .Y(n29594) );
  NOR2X1 U17526 ( .A(n29608), .B(n29609), .Y(n29607) );
  OAI22X1 U17527 ( .A(n25403), .B(n29610), .C(n25413), .D(n29611), .Y(n29609)
         );
  OAI22X1 U17528 ( .A(n25424), .B(n29612), .C(n25434), .D(n29613), .Y(n29608)
         );
  AOI22X1 U17529 ( .A(reg_file[2457]), .B(n25445), .C(reg_file[2329]), .D(
        n25456), .Y(n29606) );
  AOI22X1 U17530 ( .A(reg_file[2201]), .B(n25466), .C(reg_file[2073]), .D(
        n25477), .Y(n29605) );
  AOI21X1 U17531 ( .A(n29614), .B(n29615), .C(n25140), .Y(rd2data1040_24_) );
  NOR2X1 U17532 ( .A(n29616), .B(n29617), .Y(n29615) );
  NAND3X1 U17533 ( .A(n29618), .B(n29619), .C(n29620), .Y(n29617) );
  NOR2X1 U17534 ( .A(n29621), .B(n29622), .Y(n29620) );
  OAI22X1 U17535 ( .A(n25151), .B(n29623), .C(n25161), .D(n29624), .Y(n29622)
         );
  OAI22X1 U17536 ( .A(n25172), .B(n29625), .C(n25182), .D(n29626), .Y(n29621)
         );
  AOI22X1 U17537 ( .A(reg_file[1432]), .B(n25193), .C(reg_file[1304]), .D(
        n25204), .Y(n29619) );
  AOI22X1 U17538 ( .A(reg_file[1176]), .B(n25214), .C(reg_file[1048]), .D(
        n25225), .Y(n29618) );
  NAND3X1 U17539 ( .A(n29627), .B(n29628), .C(n29629), .Y(n29616) );
  NOR2X1 U17540 ( .A(n29630), .B(n29631), .Y(n29629) );
  OAI22X1 U17541 ( .A(n25235), .B(n29632), .C(n25245), .D(n29633), .Y(n29631)
         );
  OAI22X1 U17542 ( .A(n25256), .B(n29634), .C(n25266), .D(n29635), .Y(n29630)
         );
  AOI22X1 U17543 ( .A(reg_file[536]), .B(n25277), .C(reg_file[664]), .D(n25288), .Y(n29628) );
  AOI22X1 U17544 ( .A(reg_file[792]), .B(n25298), .C(reg_file[920]), .D(n25309), .Y(n29627) );
  NOR2X1 U17545 ( .A(n29636), .B(n29637), .Y(n29614) );
  NAND3X1 U17546 ( .A(n29638), .B(n29639), .C(n29640), .Y(n29637) );
  NOR2X1 U17547 ( .A(n29641), .B(n29642), .Y(n29640) );
  OAI22X1 U17548 ( .A(n25319), .B(n29643), .C(n25329), .D(n29644), .Y(n29642)
         );
  OAI22X1 U17549 ( .A(n25340), .B(n29645), .C(n25350), .D(n29646), .Y(n29641)
         );
  AOI22X1 U17550 ( .A(reg_file[3480]), .B(n25361), .C(reg_file[3352]), .D(
        n25372), .Y(n29639) );
  AOI22X1 U17551 ( .A(reg_file[3224]), .B(n25382), .C(reg_file[3096]), .D(
        n25393), .Y(n29638) );
  NAND3X1 U17552 ( .A(n29647), .B(n29648), .C(n29649), .Y(n29636) );
  NOR2X1 U17553 ( .A(n29650), .B(n29651), .Y(n29649) );
  OAI22X1 U17554 ( .A(n25403), .B(n29652), .C(n25413), .D(n29653), .Y(n29651)
         );
  OAI22X1 U17555 ( .A(n25424), .B(n29654), .C(n25434), .D(n29655), .Y(n29650)
         );
  AOI22X1 U17556 ( .A(reg_file[2456]), .B(n25445), .C(reg_file[2328]), .D(
        n25456), .Y(n29648) );
  AOI22X1 U17557 ( .A(reg_file[2200]), .B(n25466), .C(reg_file[2072]), .D(
        n25477), .Y(n29647) );
  AOI21X1 U17558 ( .A(n29656), .B(n29657), .C(n25140), .Y(rd2data1040_23_) );
  NOR2X1 U17559 ( .A(n29658), .B(n29659), .Y(n29657) );
  NAND3X1 U17560 ( .A(n29660), .B(n29661), .C(n29662), .Y(n29659) );
  NOR2X1 U17561 ( .A(n29663), .B(n29664), .Y(n29662) );
  OAI22X1 U17562 ( .A(n25151), .B(n29665), .C(n25161), .D(n29666), .Y(n29664)
         );
  OAI22X1 U17563 ( .A(n25172), .B(n29667), .C(n25182), .D(n29668), .Y(n29663)
         );
  AOI22X1 U17564 ( .A(reg_file[1431]), .B(n25193), .C(reg_file[1303]), .D(
        n25204), .Y(n29661) );
  AOI22X1 U17565 ( .A(reg_file[1175]), .B(n25214), .C(reg_file[1047]), .D(
        n25225), .Y(n29660) );
  NAND3X1 U17566 ( .A(n29669), .B(n29670), .C(n29671), .Y(n29658) );
  NOR2X1 U17567 ( .A(n29672), .B(n29673), .Y(n29671) );
  OAI22X1 U17568 ( .A(n25235), .B(n29674), .C(n25245), .D(n29675), .Y(n29673)
         );
  OAI22X1 U17569 ( .A(n25256), .B(n29676), .C(n25266), .D(n29677), .Y(n29672)
         );
  AOI22X1 U17570 ( .A(reg_file[535]), .B(n25277), .C(reg_file[663]), .D(n25288), .Y(n29670) );
  AOI22X1 U17571 ( .A(reg_file[791]), .B(n25298), .C(reg_file[919]), .D(n25309), .Y(n29669) );
  NOR2X1 U17572 ( .A(n29678), .B(n29679), .Y(n29656) );
  NAND3X1 U17573 ( .A(n29680), .B(n29681), .C(n29682), .Y(n29679) );
  NOR2X1 U17574 ( .A(n29683), .B(n29684), .Y(n29682) );
  OAI22X1 U17575 ( .A(n25319), .B(n29685), .C(n25329), .D(n29686), .Y(n29684)
         );
  OAI22X1 U17576 ( .A(n25340), .B(n29687), .C(n25350), .D(n29688), .Y(n29683)
         );
  AOI22X1 U17577 ( .A(reg_file[3479]), .B(n25361), .C(reg_file[3351]), .D(
        n25372), .Y(n29681) );
  AOI22X1 U17578 ( .A(reg_file[3223]), .B(n25382), .C(reg_file[3095]), .D(
        n25393), .Y(n29680) );
  NAND3X1 U17579 ( .A(n29689), .B(n29690), .C(n29691), .Y(n29678) );
  NOR2X1 U17580 ( .A(n29692), .B(n29693), .Y(n29691) );
  OAI22X1 U17581 ( .A(n25403), .B(n29694), .C(n25413), .D(n29695), .Y(n29693)
         );
  OAI22X1 U17582 ( .A(n25424), .B(n29696), .C(n25434), .D(n29697), .Y(n29692)
         );
  AOI22X1 U17583 ( .A(reg_file[2455]), .B(n25445), .C(reg_file[2327]), .D(
        n25456), .Y(n29690) );
  AOI22X1 U17584 ( .A(reg_file[2199]), .B(n25466), .C(reg_file[2071]), .D(
        n25477), .Y(n29689) );
  AOI21X1 U17585 ( .A(n29698), .B(n29699), .C(n25140), .Y(rd2data1040_22_) );
  NOR2X1 U17586 ( .A(n29700), .B(n29701), .Y(n29699) );
  NAND3X1 U17587 ( .A(n29702), .B(n29703), .C(n29704), .Y(n29701) );
  NOR2X1 U17588 ( .A(n29705), .B(n29706), .Y(n29704) );
  OAI22X1 U17589 ( .A(n25151), .B(n29707), .C(n25161), .D(n29708), .Y(n29706)
         );
  OAI22X1 U17590 ( .A(n25172), .B(n29709), .C(n25182), .D(n29710), .Y(n29705)
         );
  AOI22X1 U17591 ( .A(reg_file[1430]), .B(n25193), .C(reg_file[1302]), .D(
        n25204), .Y(n29703) );
  AOI22X1 U17592 ( .A(reg_file[1174]), .B(n25214), .C(reg_file[1046]), .D(
        n25225), .Y(n29702) );
  NAND3X1 U17593 ( .A(n29711), .B(n29712), .C(n29713), .Y(n29700) );
  NOR2X1 U17594 ( .A(n29714), .B(n29715), .Y(n29713) );
  OAI22X1 U17595 ( .A(n25235), .B(n29716), .C(n25245), .D(n29717), .Y(n29715)
         );
  OAI22X1 U17596 ( .A(n25256), .B(n29718), .C(n25266), .D(n29719), .Y(n29714)
         );
  AOI22X1 U17597 ( .A(reg_file[534]), .B(n25277), .C(reg_file[662]), .D(n25288), .Y(n29712) );
  AOI22X1 U17598 ( .A(reg_file[790]), .B(n25298), .C(reg_file[918]), .D(n25309), .Y(n29711) );
  NOR2X1 U17599 ( .A(n29720), .B(n29721), .Y(n29698) );
  NAND3X1 U17600 ( .A(n29722), .B(n29723), .C(n29724), .Y(n29721) );
  NOR2X1 U17601 ( .A(n29725), .B(n29726), .Y(n29724) );
  OAI22X1 U17602 ( .A(n25319), .B(n29727), .C(n25329), .D(n29728), .Y(n29726)
         );
  OAI22X1 U17603 ( .A(n25340), .B(n29729), .C(n25350), .D(n29730), .Y(n29725)
         );
  AOI22X1 U17604 ( .A(reg_file[3478]), .B(n25361), .C(reg_file[3350]), .D(
        n25372), .Y(n29723) );
  AOI22X1 U17605 ( .A(reg_file[3222]), .B(n25382), .C(reg_file[3094]), .D(
        n25393), .Y(n29722) );
  NAND3X1 U17606 ( .A(n29731), .B(n29732), .C(n29733), .Y(n29720) );
  NOR2X1 U17607 ( .A(n29734), .B(n29735), .Y(n29733) );
  OAI22X1 U17608 ( .A(n25403), .B(n29736), .C(n25413), .D(n29737), .Y(n29735)
         );
  OAI22X1 U17609 ( .A(n25424), .B(n29738), .C(n25434), .D(n29739), .Y(n29734)
         );
  AOI22X1 U17610 ( .A(reg_file[2454]), .B(n25445), .C(reg_file[2326]), .D(
        n25456), .Y(n29732) );
  AOI22X1 U17611 ( .A(reg_file[2198]), .B(n25466), .C(reg_file[2070]), .D(
        n25477), .Y(n29731) );
  AOI21X1 U17612 ( .A(n29740), .B(n29741), .C(n25140), .Y(rd2data1040_21_) );
  NOR2X1 U17613 ( .A(n29742), .B(n29743), .Y(n29741) );
  NAND3X1 U17614 ( .A(n29744), .B(n29745), .C(n29746), .Y(n29743) );
  NOR2X1 U17615 ( .A(n29747), .B(n29748), .Y(n29746) );
  OAI22X1 U17616 ( .A(n25151), .B(n29749), .C(n25161), .D(n29750), .Y(n29748)
         );
  OAI22X1 U17617 ( .A(n25172), .B(n29751), .C(n25182), .D(n29752), .Y(n29747)
         );
  AOI22X1 U17618 ( .A(reg_file[1429]), .B(n25193), .C(reg_file[1301]), .D(
        n25204), .Y(n29745) );
  AOI22X1 U17619 ( .A(reg_file[1173]), .B(n25214), .C(reg_file[1045]), .D(
        n25225), .Y(n29744) );
  NAND3X1 U17620 ( .A(n29753), .B(n29754), .C(n29755), .Y(n29742) );
  NOR2X1 U17621 ( .A(n29756), .B(n29757), .Y(n29755) );
  OAI22X1 U17622 ( .A(n25235), .B(n29758), .C(n25245), .D(n29759), .Y(n29757)
         );
  OAI22X1 U17623 ( .A(n25256), .B(n29760), .C(n25266), .D(n29761), .Y(n29756)
         );
  AOI22X1 U17624 ( .A(reg_file[533]), .B(n25277), .C(reg_file[661]), .D(n25288), .Y(n29754) );
  AOI22X1 U17625 ( .A(reg_file[789]), .B(n25298), .C(reg_file[917]), .D(n25309), .Y(n29753) );
  NOR2X1 U17626 ( .A(n29762), .B(n29763), .Y(n29740) );
  NAND3X1 U17627 ( .A(n29764), .B(n29765), .C(n29766), .Y(n29763) );
  NOR2X1 U17628 ( .A(n29767), .B(n29768), .Y(n29766) );
  OAI22X1 U17629 ( .A(n25319), .B(n29769), .C(n25329), .D(n29770), .Y(n29768)
         );
  OAI22X1 U17630 ( .A(n25340), .B(n29771), .C(n25350), .D(n29772), .Y(n29767)
         );
  AOI22X1 U17631 ( .A(reg_file[3477]), .B(n25361), .C(reg_file[3349]), .D(
        n25372), .Y(n29765) );
  AOI22X1 U17632 ( .A(reg_file[3221]), .B(n25382), .C(reg_file[3093]), .D(
        n25393), .Y(n29764) );
  NAND3X1 U17633 ( .A(n29773), .B(n29774), .C(n29775), .Y(n29762) );
  NOR2X1 U17634 ( .A(n29776), .B(n29777), .Y(n29775) );
  OAI22X1 U17635 ( .A(n25403), .B(n29778), .C(n25413), .D(n29779), .Y(n29777)
         );
  OAI22X1 U17636 ( .A(n25424), .B(n29780), .C(n25434), .D(n29781), .Y(n29776)
         );
  AOI22X1 U17637 ( .A(reg_file[2453]), .B(n25445), .C(reg_file[2325]), .D(
        n25456), .Y(n29774) );
  AOI22X1 U17638 ( .A(reg_file[2197]), .B(n25466), .C(reg_file[2069]), .D(
        n25477), .Y(n29773) );
  AOI21X1 U17639 ( .A(n29782), .B(n29783), .C(n25140), .Y(rd2data1040_20_) );
  NOR2X1 U17640 ( .A(n29784), .B(n29785), .Y(n29783) );
  NAND3X1 U17641 ( .A(n29786), .B(n29787), .C(n29788), .Y(n29785) );
  NOR2X1 U17642 ( .A(n29789), .B(n29790), .Y(n29788) );
  OAI22X1 U17643 ( .A(n25151), .B(n29791), .C(n25161), .D(n29792), .Y(n29790)
         );
  OAI22X1 U17644 ( .A(n25172), .B(n29793), .C(n25182), .D(n29794), .Y(n29789)
         );
  AOI22X1 U17645 ( .A(reg_file[1428]), .B(n25193), .C(reg_file[1300]), .D(
        n25204), .Y(n29787) );
  AOI22X1 U17646 ( .A(reg_file[1172]), .B(n25214), .C(reg_file[1044]), .D(
        n25225), .Y(n29786) );
  NAND3X1 U17647 ( .A(n29795), .B(n29796), .C(n29797), .Y(n29784) );
  NOR2X1 U17648 ( .A(n29798), .B(n29799), .Y(n29797) );
  OAI22X1 U17649 ( .A(n25235), .B(n29800), .C(n25245), .D(n29801), .Y(n29799)
         );
  OAI22X1 U17650 ( .A(n25256), .B(n29802), .C(n25266), .D(n29803), .Y(n29798)
         );
  AOI22X1 U17651 ( .A(reg_file[532]), .B(n25277), .C(reg_file[660]), .D(n25288), .Y(n29796) );
  AOI22X1 U17652 ( .A(reg_file[788]), .B(n25298), .C(reg_file[916]), .D(n25309), .Y(n29795) );
  NOR2X1 U17653 ( .A(n29804), .B(n29805), .Y(n29782) );
  NAND3X1 U17654 ( .A(n29806), .B(n29807), .C(n29808), .Y(n29805) );
  NOR2X1 U17655 ( .A(n29809), .B(n29810), .Y(n29808) );
  OAI22X1 U17656 ( .A(n25319), .B(n29811), .C(n25329), .D(n29812), .Y(n29810)
         );
  OAI22X1 U17657 ( .A(n25340), .B(n29813), .C(n25350), .D(n29814), .Y(n29809)
         );
  AOI22X1 U17658 ( .A(reg_file[3476]), .B(n25361), .C(reg_file[3348]), .D(
        n25372), .Y(n29807) );
  AOI22X1 U17659 ( .A(reg_file[3220]), .B(n25382), .C(reg_file[3092]), .D(
        n25393), .Y(n29806) );
  NAND3X1 U17660 ( .A(n29815), .B(n29816), .C(n29817), .Y(n29804) );
  NOR2X1 U17661 ( .A(n29818), .B(n29819), .Y(n29817) );
  OAI22X1 U17662 ( .A(n25403), .B(n29820), .C(n25413), .D(n29821), .Y(n29819)
         );
  OAI22X1 U17663 ( .A(n25424), .B(n29822), .C(n25434), .D(n29823), .Y(n29818)
         );
  AOI22X1 U17664 ( .A(reg_file[2452]), .B(n25445), .C(reg_file[2324]), .D(
        n25456), .Y(n29816) );
  AOI22X1 U17665 ( .A(reg_file[2196]), .B(n25466), .C(reg_file[2068]), .D(
        n25477), .Y(n29815) );
  AOI21X1 U17666 ( .A(n29824), .B(n29825), .C(n25140), .Y(rd2data1040_1_) );
  NOR2X1 U17667 ( .A(n29826), .B(n29827), .Y(n29825) );
  NAND3X1 U17668 ( .A(n29828), .B(n29829), .C(n29830), .Y(n29827) );
  NOR2X1 U17669 ( .A(n29831), .B(n29832), .Y(n29830) );
  OAI22X1 U17670 ( .A(n25151), .B(n29833), .C(n25161), .D(n29834), .Y(n29832)
         );
  OAI22X1 U17671 ( .A(n25172), .B(n29835), .C(n25182), .D(n29836), .Y(n29831)
         );
  AOI22X1 U17672 ( .A(reg_file[1409]), .B(n25193), .C(reg_file[1281]), .D(
        n25204), .Y(n29829) );
  AOI22X1 U17673 ( .A(reg_file[1153]), .B(n25214), .C(reg_file[1025]), .D(
        n25225), .Y(n29828) );
  NAND3X1 U17674 ( .A(n29837), .B(n29838), .C(n29839), .Y(n29826) );
  NOR2X1 U17675 ( .A(n29840), .B(n29841), .Y(n29839) );
  OAI22X1 U17676 ( .A(n25235), .B(n29842), .C(n25245), .D(n29843), .Y(n29841)
         );
  OAI22X1 U17677 ( .A(n25256), .B(n29844), .C(n25266), .D(n29845), .Y(n29840)
         );
  AOI22X1 U17678 ( .A(reg_file[513]), .B(n25277), .C(reg_file[641]), .D(n25288), .Y(n29838) );
  AOI22X1 U17679 ( .A(reg_file[769]), .B(n25298), .C(reg_file[897]), .D(n25309), .Y(n29837) );
  NOR2X1 U17680 ( .A(n29846), .B(n29847), .Y(n29824) );
  NAND3X1 U17681 ( .A(n29848), .B(n29849), .C(n29850), .Y(n29847) );
  NOR2X1 U17682 ( .A(n29851), .B(n29852), .Y(n29850) );
  OAI22X1 U17683 ( .A(n25319), .B(n29853), .C(n25329), .D(n29854), .Y(n29852)
         );
  OAI22X1 U17684 ( .A(n25340), .B(n29855), .C(n25350), .D(n29856), .Y(n29851)
         );
  AOI22X1 U17685 ( .A(reg_file[3457]), .B(n25361), .C(reg_file[3329]), .D(
        n25372), .Y(n29849) );
  AOI22X1 U17686 ( .A(reg_file[3201]), .B(n25382), .C(reg_file[3073]), .D(
        n25393), .Y(n29848) );
  NAND3X1 U17687 ( .A(n29857), .B(n29858), .C(n29859), .Y(n29846) );
  NOR2X1 U17688 ( .A(n29860), .B(n29861), .Y(n29859) );
  OAI22X1 U17689 ( .A(n25403), .B(n29862), .C(n25413), .D(n29863), .Y(n29861)
         );
  OAI22X1 U17690 ( .A(n25424), .B(n29864), .C(n25434), .D(n29865), .Y(n29860)
         );
  AOI22X1 U17691 ( .A(reg_file[2433]), .B(n25445), .C(reg_file[2305]), .D(
        n25456), .Y(n29858) );
  AOI22X1 U17692 ( .A(reg_file[2177]), .B(n25466), .C(reg_file[2049]), .D(
        n25477), .Y(n29857) );
  AOI21X1 U17693 ( .A(n29866), .B(n29867), .C(n25140), .Y(rd2data1040_19_) );
  NOR2X1 U17694 ( .A(n29868), .B(n29869), .Y(n29867) );
  NAND3X1 U17695 ( .A(n29870), .B(n29871), .C(n29872), .Y(n29869) );
  NOR2X1 U17696 ( .A(n29873), .B(n29874), .Y(n29872) );
  OAI22X1 U17697 ( .A(n25150), .B(n29875), .C(n25161), .D(n29876), .Y(n29874)
         );
  OAI22X1 U17698 ( .A(n25171), .B(n29877), .C(n25182), .D(n29878), .Y(n29873)
         );
  AOI22X1 U17699 ( .A(reg_file[1427]), .B(n25193), .C(reg_file[1299]), .D(
        n25203), .Y(n29871) );
  AOI22X1 U17700 ( .A(reg_file[1171]), .B(n25214), .C(reg_file[1043]), .D(
        n25224), .Y(n29870) );
  NAND3X1 U17701 ( .A(n29879), .B(n29880), .C(n29881), .Y(n29868) );
  NOR2X1 U17702 ( .A(n29882), .B(n29883), .Y(n29881) );
  OAI22X1 U17703 ( .A(n25234), .B(n29884), .C(n25245), .D(n29885), .Y(n29883)
         );
  OAI22X1 U17704 ( .A(n25255), .B(n29886), .C(n25266), .D(n29887), .Y(n29882)
         );
  AOI22X1 U17705 ( .A(reg_file[531]), .B(n25277), .C(reg_file[659]), .D(n25287), .Y(n29880) );
  AOI22X1 U17706 ( .A(reg_file[787]), .B(n25298), .C(reg_file[915]), .D(n25308), .Y(n29879) );
  NOR2X1 U17707 ( .A(n29888), .B(n29889), .Y(n29866) );
  NAND3X1 U17708 ( .A(n29890), .B(n29891), .C(n29892), .Y(n29889) );
  NOR2X1 U17709 ( .A(n29893), .B(n29894), .Y(n29892) );
  OAI22X1 U17710 ( .A(n25318), .B(n29895), .C(n25329), .D(n29896), .Y(n29894)
         );
  OAI22X1 U17711 ( .A(n25339), .B(n29897), .C(n25350), .D(n29898), .Y(n29893)
         );
  AOI22X1 U17712 ( .A(reg_file[3475]), .B(n25361), .C(reg_file[3347]), .D(
        n25371), .Y(n29891) );
  AOI22X1 U17713 ( .A(reg_file[3219]), .B(n25382), .C(reg_file[3091]), .D(
        n25392), .Y(n29890) );
  NAND3X1 U17714 ( .A(n29899), .B(n29900), .C(n29901), .Y(n29888) );
  NOR2X1 U17715 ( .A(n29902), .B(n29903), .Y(n29901) );
  OAI22X1 U17716 ( .A(n25402), .B(n29904), .C(n25413), .D(n29905), .Y(n29903)
         );
  OAI22X1 U17717 ( .A(n25423), .B(n29906), .C(n25434), .D(n29907), .Y(n29902)
         );
  AOI22X1 U17718 ( .A(reg_file[2451]), .B(n25445), .C(reg_file[2323]), .D(
        n25455), .Y(n29900) );
  AOI22X1 U17719 ( .A(reg_file[2195]), .B(n25466), .C(reg_file[2067]), .D(
        n25476), .Y(n29899) );
  AOI21X1 U17720 ( .A(n29908), .B(n29909), .C(n25140), .Y(rd2data1040_18_) );
  NOR2X1 U17721 ( .A(n29910), .B(n29911), .Y(n29909) );
  NAND3X1 U17722 ( .A(n29912), .B(n29913), .C(n29914), .Y(n29911) );
  NOR2X1 U17723 ( .A(n29915), .B(n29916), .Y(n29914) );
  OAI22X1 U17724 ( .A(n25150), .B(n29917), .C(n25161), .D(n29918), .Y(n29916)
         );
  OAI22X1 U17725 ( .A(n25171), .B(n29919), .C(n25182), .D(n29920), .Y(n29915)
         );
  AOI22X1 U17726 ( .A(reg_file[1426]), .B(n25193), .C(reg_file[1298]), .D(
        n25203), .Y(n29913) );
  AOI22X1 U17727 ( .A(reg_file[1170]), .B(n25214), .C(reg_file[1042]), .D(
        n25224), .Y(n29912) );
  NAND3X1 U17728 ( .A(n29921), .B(n29922), .C(n29923), .Y(n29910) );
  NOR2X1 U17729 ( .A(n29924), .B(n29925), .Y(n29923) );
  OAI22X1 U17730 ( .A(n25234), .B(n29926), .C(n25245), .D(n29927), .Y(n29925)
         );
  OAI22X1 U17731 ( .A(n25255), .B(n29928), .C(n25266), .D(n29929), .Y(n29924)
         );
  AOI22X1 U17732 ( .A(reg_file[530]), .B(n25277), .C(reg_file[658]), .D(n25287), .Y(n29922) );
  AOI22X1 U17733 ( .A(reg_file[786]), .B(n25298), .C(reg_file[914]), .D(n25308), .Y(n29921) );
  NOR2X1 U17734 ( .A(n29930), .B(n29931), .Y(n29908) );
  NAND3X1 U17735 ( .A(n29932), .B(n29933), .C(n29934), .Y(n29931) );
  NOR2X1 U17736 ( .A(n29935), .B(n29936), .Y(n29934) );
  OAI22X1 U17737 ( .A(n25318), .B(n29937), .C(n25329), .D(n29938), .Y(n29936)
         );
  OAI22X1 U17738 ( .A(n25339), .B(n29939), .C(n25350), .D(n29940), .Y(n29935)
         );
  AOI22X1 U17739 ( .A(reg_file[3474]), .B(n25361), .C(reg_file[3346]), .D(
        n25371), .Y(n29933) );
  AOI22X1 U17740 ( .A(reg_file[3218]), .B(n25382), .C(reg_file[3090]), .D(
        n25392), .Y(n29932) );
  NAND3X1 U17741 ( .A(n29941), .B(n29942), .C(n29943), .Y(n29930) );
  NOR2X1 U17742 ( .A(n29944), .B(n29945), .Y(n29943) );
  OAI22X1 U17743 ( .A(n25402), .B(n29946), .C(n25413), .D(n29947), .Y(n29945)
         );
  OAI22X1 U17744 ( .A(n25423), .B(n29948), .C(n25434), .D(n29949), .Y(n29944)
         );
  AOI22X1 U17745 ( .A(reg_file[2450]), .B(n25445), .C(reg_file[2322]), .D(
        n25455), .Y(n29942) );
  AOI22X1 U17746 ( .A(reg_file[2194]), .B(n25466), .C(reg_file[2066]), .D(
        n25476), .Y(n29941) );
  AOI21X1 U17747 ( .A(n29950), .B(n29951), .C(n25140), .Y(rd2data1040_17_) );
  NOR2X1 U17748 ( .A(n29952), .B(n29953), .Y(n29951) );
  NAND3X1 U17749 ( .A(n29954), .B(n29955), .C(n29956), .Y(n29953) );
  NOR2X1 U17750 ( .A(n29957), .B(n29958), .Y(n29956) );
  OAI22X1 U17751 ( .A(n25150), .B(n29959), .C(n25161), .D(n29960), .Y(n29958)
         );
  OAI22X1 U17752 ( .A(n25171), .B(n29961), .C(n25182), .D(n29962), .Y(n29957)
         );
  AOI22X1 U17753 ( .A(reg_file[1425]), .B(n25193), .C(reg_file[1297]), .D(
        n25203), .Y(n29955) );
  AOI22X1 U17754 ( .A(reg_file[1169]), .B(n25214), .C(reg_file[1041]), .D(
        n25224), .Y(n29954) );
  NAND3X1 U17755 ( .A(n29963), .B(n29964), .C(n29965), .Y(n29952) );
  NOR2X1 U17756 ( .A(n29966), .B(n29967), .Y(n29965) );
  OAI22X1 U17757 ( .A(n25234), .B(n29968), .C(n25245), .D(n29969), .Y(n29967)
         );
  OAI22X1 U17758 ( .A(n25255), .B(n29970), .C(n25266), .D(n29971), .Y(n29966)
         );
  AOI22X1 U17759 ( .A(reg_file[529]), .B(n25277), .C(reg_file[657]), .D(n25287), .Y(n29964) );
  AOI22X1 U17760 ( .A(reg_file[785]), .B(n25298), .C(reg_file[913]), .D(n25308), .Y(n29963) );
  NOR2X1 U17761 ( .A(n29972), .B(n29973), .Y(n29950) );
  NAND3X1 U17762 ( .A(n29974), .B(n29975), .C(n29976), .Y(n29973) );
  NOR2X1 U17763 ( .A(n29977), .B(n29978), .Y(n29976) );
  OAI22X1 U17764 ( .A(n25318), .B(n29979), .C(n25329), .D(n29980), .Y(n29978)
         );
  OAI22X1 U17765 ( .A(n25339), .B(n29981), .C(n25350), .D(n29982), .Y(n29977)
         );
  AOI22X1 U17766 ( .A(reg_file[3473]), .B(n25361), .C(reg_file[3345]), .D(
        n25371), .Y(n29975) );
  AOI22X1 U17767 ( .A(reg_file[3217]), .B(n25382), .C(reg_file[3089]), .D(
        n25392), .Y(n29974) );
  NAND3X1 U17768 ( .A(n29983), .B(n29984), .C(n29985), .Y(n29972) );
  NOR2X1 U17769 ( .A(n29986), .B(n29987), .Y(n29985) );
  OAI22X1 U17770 ( .A(n25402), .B(n29988), .C(n25413), .D(n29989), .Y(n29987)
         );
  OAI22X1 U17771 ( .A(n25423), .B(n29990), .C(n25434), .D(n29991), .Y(n29986)
         );
  AOI22X1 U17772 ( .A(reg_file[2449]), .B(n25445), .C(reg_file[2321]), .D(
        n25455), .Y(n29984) );
  AOI22X1 U17773 ( .A(reg_file[2193]), .B(n25466), .C(reg_file[2065]), .D(
        n25476), .Y(n29983) );
  AOI21X1 U17774 ( .A(n29992), .B(n29993), .C(n25139), .Y(rd2data1040_16_) );
  NOR2X1 U17775 ( .A(n29994), .B(n29995), .Y(n29993) );
  NAND3X1 U17776 ( .A(n29996), .B(n29997), .C(n29998), .Y(n29995) );
  NOR2X1 U17777 ( .A(n29999), .B(n30000), .Y(n29998) );
  OAI22X1 U17778 ( .A(n25150), .B(n30001), .C(n25160), .D(n30002), .Y(n30000)
         );
  OAI22X1 U17779 ( .A(n25171), .B(n30003), .C(n25181), .D(n30004), .Y(n29999)
         );
  AOI22X1 U17780 ( .A(reg_file[1424]), .B(n25192), .C(reg_file[1296]), .D(
        n25203), .Y(n29997) );
  AOI22X1 U17781 ( .A(reg_file[1168]), .B(n25213), .C(reg_file[1040]), .D(
        n25224), .Y(n29996) );
  NAND3X1 U17782 ( .A(n30005), .B(n30006), .C(n30007), .Y(n29994) );
  NOR2X1 U17783 ( .A(n30008), .B(n30009), .Y(n30007) );
  OAI22X1 U17784 ( .A(n25234), .B(n30010), .C(n25244), .D(n30011), .Y(n30009)
         );
  OAI22X1 U17785 ( .A(n25255), .B(n30012), .C(n25265), .D(n30013), .Y(n30008)
         );
  AOI22X1 U17786 ( .A(reg_file[528]), .B(n25276), .C(reg_file[656]), .D(n25287), .Y(n30006) );
  AOI22X1 U17787 ( .A(reg_file[784]), .B(n25297), .C(reg_file[912]), .D(n25308), .Y(n30005) );
  NOR2X1 U17788 ( .A(n30014), .B(n30015), .Y(n29992) );
  NAND3X1 U17789 ( .A(n30016), .B(n30017), .C(n30018), .Y(n30015) );
  NOR2X1 U17790 ( .A(n30019), .B(n30020), .Y(n30018) );
  OAI22X1 U17791 ( .A(n25318), .B(n30021), .C(n25328), .D(n30022), .Y(n30020)
         );
  OAI22X1 U17792 ( .A(n25339), .B(n30023), .C(n25349), .D(n30024), .Y(n30019)
         );
  AOI22X1 U17793 ( .A(reg_file[3472]), .B(n25360), .C(reg_file[3344]), .D(
        n25371), .Y(n30017) );
  AOI22X1 U17794 ( .A(reg_file[3216]), .B(n25381), .C(reg_file[3088]), .D(
        n25392), .Y(n30016) );
  NAND3X1 U17795 ( .A(n30025), .B(n30026), .C(n30027), .Y(n30014) );
  NOR2X1 U17796 ( .A(n30028), .B(n30029), .Y(n30027) );
  OAI22X1 U17797 ( .A(n25402), .B(n30030), .C(n25412), .D(n30031), .Y(n30029)
         );
  OAI22X1 U17798 ( .A(n25423), .B(n30032), .C(n25433), .D(n30033), .Y(n30028)
         );
  AOI22X1 U17799 ( .A(reg_file[2448]), .B(n25444), .C(reg_file[2320]), .D(
        n25455), .Y(n30026) );
  AOI22X1 U17800 ( .A(reg_file[2192]), .B(n25465), .C(reg_file[2064]), .D(
        n25476), .Y(n30025) );
  AOI21X1 U17801 ( .A(n30034), .B(n30035), .C(n25139), .Y(rd2data1040_15_) );
  NOR2X1 U17802 ( .A(n30036), .B(n30037), .Y(n30035) );
  NAND3X1 U17803 ( .A(n30038), .B(n30039), .C(n30040), .Y(n30037) );
  NOR2X1 U17804 ( .A(n30041), .B(n30042), .Y(n30040) );
  OAI22X1 U17805 ( .A(n25150), .B(n30043), .C(n25160), .D(n30044), .Y(n30042)
         );
  OAI22X1 U17806 ( .A(n25171), .B(n30045), .C(n25181), .D(n30046), .Y(n30041)
         );
  AOI22X1 U17807 ( .A(reg_file[1423]), .B(n25192), .C(reg_file[1295]), .D(
        n25203), .Y(n30039) );
  AOI22X1 U17808 ( .A(reg_file[1167]), .B(n25213), .C(reg_file[1039]), .D(
        n25224), .Y(n30038) );
  NAND3X1 U17809 ( .A(n30047), .B(n30048), .C(n30049), .Y(n30036) );
  NOR2X1 U17810 ( .A(n30050), .B(n30051), .Y(n30049) );
  OAI22X1 U17811 ( .A(n25234), .B(n30052), .C(n25244), .D(n30053), .Y(n30051)
         );
  OAI22X1 U17812 ( .A(n25255), .B(n30054), .C(n25265), .D(n30055), .Y(n30050)
         );
  AOI22X1 U17813 ( .A(reg_file[527]), .B(n25276), .C(reg_file[655]), .D(n25287), .Y(n30048) );
  AOI22X1 U17814 ( .A(reg_file[783]), .B(n25297), .C(reg_file[911]), .D(n25308), .Y(n30047) );
  NOR2X1 U17815 ( .A(n30056), .B(n30057), .Y(n30034) );
  NAND3X1 U17816 ( .A(n30058), .B(n30059), .C(n30060), .Y(n30057) );
  NOR2X1 U17817 ( .A(n30061), .B(n30062), .Y(n30060) );
  OAI22X1 U17818 ( .A(n25318), .B(n30063), .C(n25328), .D(n30064), .Y(n30062)
         );
  OAI22X1 U17819 ( .A(n25339), .B(n30065), .C(n25349), .D(n30066), .Y(n30061)
         );
  AOI22X1 U17820 ( .A(reg_file[3471]), .B(n25360), .C(reg_file[3343]), .D(
        n25371), .Y(n30059) );
  AOI22X1 U17821 ( .A(reg_file[3215]), .B(n25381), .C(reg_file[3087]), .D(
        n25392), .Y(n30058) );
  NAND3X1 U17822 ( .A(n30067), .B(n30068), .C(n30069), .Y(n30056) );
  NOR2X1 U17823 ( .A(n30070), .B(n30071), .Y(n30069) );
  OAI22X1 U17824 ( .A(n25402), .B(n30072), .C(n25412), .D(n30073), .Y(n30071)
         );
  OAI22X1 U17825 ( .A(n25423), .B(n30074), .C(n25433), .D(n30075), .Y(n30070)
         );
  AOI22X1 U17826 ( .A(reg_file[2447]), .B(n25444), .C(reg_file[2319]), .D(
        n25455), .Y(n30068) );
  AOI22X1 U17827 ( .A(reg_file[2191]), .B(n25465), .C(reg_file[2063]), .D(
        n25476), .Y(n30067) );
  AOI21X1 U17828 ( .A(n30076), .B(n30077), .C(n25139), .Y(rd2data1040_14_) );
  NOR2X1 U17829 ( .A(n30078), .B(n30079), .Y(n30077) );
  NAND3X1 U17830 ( .A(n30080), .B(n30081), .C(n30082), .Y(n30079) );
  NOR2X1 U17831 ( .A(n30083), .B(n30084), .Y(n30082) );
  OAI22X1 U17832 ( .A(n25150), .B(n30085), .C(n25160), .D(n30086), .Y(n30084)
         );
  OAI22X1 U17833 ( .A(n25171), .B(n30087), .C(n25181), .D(n30088), .Y(n30083)
         );
  AOI22X1 U17834 ( .A(reg_file[1422]), .B(n25192), .C(reg_file[1294]), .D(
        n25203), .Y(n30081) );
  AOI22X1 U17835 ( .A(reg_file[1166]), .B(n25213), .C(reg_file[1038]), .D(
        n25224), .Y(n30080) );
  NAND3X1 U17836 ( .A(n30089), .B(n30090), .C(n30091), .Y(n30078) );
  NOR2X1 U17837 ( .A(n30092), .B(n30093), .Y(n30091) );
  OAI22X1 U17838 ( .A(n25234), .B(n30094), .C(n25244), .D(n30095), .Y(n30093)
         );
  OAI22X1 U17839 ( .A(n25255), .B(n30096), .C(n25265), .D(n30097), .Y(n30092)
         );
  AOI22X1 U17840 ( .A(reg_file[526]), .B(n25276), .C(reg_file[654]), .D(n25287), .Y(n30090) );
  AOI22X1 U17841 ( .A(reg_file[782]), .B(n25297), .C(reg_file[910]), .D(n25308), .Y(n30089) );
  NOR2X1 U17842 ( .A(n30098), .B(n30099), .Y(n30076) );
  NAND3X1 U17843 ( .A(n30100), .B(n30101), .C(n30102), .Y(n30099) );
  NOR2X1 U17844 ( .A(n30103), .B(n30104), .Y(n30102) );
  OAI22X1 U17845 ( .A(n25318), .B(n30105), .C(n25328), .D(n30106), .Y(n30104)
         );
  OAI22X1 U17846 ( .A(n25339), .B(n30107), .C(n25349), .D(n30108), .Y(n30103)
         );
  AOI22X1 U17847 ( .A(reg_file[3470]), .B(n25360), .C(reg_file[3342]), .D(
        n25371), .Y(n30101) );
  AOI22X1 U17848 ( .A(reg_file[3214]), .B(n25381), .C(reg_file[3086]), .D(
        n25392), .Y(n30100) );
  NAND3X1 U17849 ( .A(n30109), .B(n30110), .C(n30111), .Y(n30098) );
  NOR2X1 U17850 ( .A(n30112), .B(n30113), .Y(n30111) );
  OAI22X1 U17851 ( .A(n25402), .B(n30114), .C(n25412), .D(n30115), .Y(n30113)
         );
  OAI22X1 U17852 ( .A(n25423), .B(n30116), .C(n25433), .D(n30117), .Y(n30112)
         );
  AOI22X1 U17853 ( .A(reg_file[2446]), .B(n25444), .C(reg_file[2318]), .D(
        n25455), .Y(n30110) );
  AOI22X1 U17854 ( .A(reg_file[2190]), .B(n25465), .C(reg_file[2062]), .D(
        n25476), .Y(n30109) );
  AOI21X1 U17855 ( .A(n30118), .B(n30119), .C(n25139), .Y(rd2data1040_13_) );
  NOR2X1 U17856 ( .A(n30120), .B(n30121), .Y(n30119) );
  NAND3X1 U17857 ( .A(n30122), .B(n30123), .C(n30124), .Y(n30121) );
  NOR2X1 U17858 ( .A(n30125), .B(n30126), .Y(n30124) );
  OAI22X1 U17859 ( .A(n25150), .B(n30127), .C(n25160), .D(n30128), .Y(n30126)
         );
  OAI22X1 U17860 ( .A(n25171), .B(n30129), .C(n25181), .D(n30130), .Y(n30125)
         );
  AOI22X1 U17861 ( .A(reg_file[1421]), .B(n25192), .C(reg_file[1293]), .D(
        n25203), .Y(n30123) );
  AOI22X1 U17862 ( .A(reg_file[1165]), .B(n25213), .C(reg_file[1037]), .D(
        n25224), .Y(n30122) );
  NAND3X1 U17863 ( .A(n30131), .B(n30132), .C(n30133), .Y(n30120) );
  NOR2X1 U17864 ( .A(n30134), .B(n30135), .Y(n30133) );
  OAI22X1 U17865 ( .A(n25234), .B(n30136), .C(n25244), .D(n30137), .Y(n30135)
         );
  OAI22X1 U17866 ( .A(n25255), .B(n30138), .C(n25265), .D(n30139), .Y(n30134)
         );
  AOI22X1 U17867 ( .A(reg_file[525]), .B(n25276), .C(reg_file[653]), .D(n25287), .Y(n30132) );
  AOI22X1 U17868 ( .A(reg_file[781]), .B(n25297), .C(reg_file[909]), .D(n25308), .Y(n30131) );
  NOR2X1 U17869 ( .A(n30140), .B(n30141), .Y(n30118) );
  NAND3X1 U17870 ( .A(n30142), .B(n30143), .C(n30144), .Y(n30141) );
  NOR2X1 U17871 ( .A(n30145), .B(n30146), .Y(n30144) );
  OAI22X1 U17872 ( .A(n25318), .B(n30147), .C(n25328), .D(n30148), .Y(n30146)
         );
  OAI22X1 U17873 ( .A(n25339), .B(n30149), .C(n25349), .D(n30150), .Y(n30145)
         );
  AOI22X1 U17874 ( .A(reg_file[3469]), .B(n25360), .C(reg_file[3341]), .D(
        n25371), .Y(n30143) );
  AOI22X1 U17875 ( .A(reg_file[3213]), .B(n25381), .C(reg_file[3085]), .D(
        n25392), .Y(n30142) );
  NAND3X1 U17876 ( .A(n30151), .B(n30152), .C(n30153), .Y(n30140) );
  NOR2X1 U17877 ( .A(n30154), .B(n30155), .Y(n30153) );
  OAI22X1 U17878 ( .A(n25402), .B(n30156), .C(n25412), .D(n30157), .Y(n30155)
         );
  OAI22X1 U17879 ( .A(n25423), .B(n30158), .C(n25433), .D(n30159), .Y(n30154)
         );
  AOI22X1 U17880 ( .A(reg_file[2445]), .B(n25444), .C(reg_file[2317]), .D(
        n25455), .Y(n30152) );
  AOI22X1 U17881 ( .A(reg_file[2189]), .B(n25465), .C(reg_file[2061]), .D(
        n25476), .Y(n30151) );
  AOI21X1 U17882 ( .A(n30160), .B(n30161), .C(n25139), .Y(rd2data1040_12_) );
  NOR2X1 U17883 ( .A(n30162), .B(n30163), .Y(n30161) );
  NAND3X1 U17884 ( .A(n30164), .B(n30165), .C(n30166), .Y(n30163) );
  NOR2X1 U17885 ( .A(n30167), .B(n30168), .Y(n30166) );
  OAI22X1 U17886 ( .A(n25150), .B(n30169), .C(n25160), .D(n30170), .Y(n30168)
         );
  OAI22X1 U17887 ( .A(n25171), .B(n30171), .C(n25181), .D(n30172), .Y(n30167)
         );
  AOI22X1 U17888 ( .A(reg_file[1420]), .B(n25192), .C(reg_file[1292]), .D(
        n25203), .Y(n30165) );
  AOI22X1 U17889 ( .A(reg_file[1164]), .B(n25213), .C(reg_file[1036]), .D(
        n25224), .Y(n30164) );
  NAND3X1 U17890 ( .A(n30173), .B(n30174), .C(n30175), .Y(n30162) );
  NOR2X1 U17891 ( .A(n30176), .B(n30177), .Y(n30175) );
  OAI22X1 U17892 ( .A(n25234), .B(n30178), .C(n25244), .D(n30179), .Y(n30177)
         );
  OAI22X1 U17893 ( .A(n25255), .B(n30180), .C(n25265), .D(n30181), .Y(n30176)
         );
  AOI22X1 U17894 ( .A(reg_file[524]), .B(n25276), .C(reg_file[652]), .D(n25287), .Y(n30174) );
  AOI22X1 U17895 ( .A(reg_file[780]), .B(n25297), .C(reg_file[908]), .D(n25308), .Y(n30173) );
  NOR2X1 U17896 ( .A(n30182), .B(n30183), .Y(n30160) );
  NAND3X1 U17897 ( .A(n30184), .B(n30185), .C(n30186), .Y(n30183) );
  NOR2X1 U17898 ( .A(n30187), .B(n30188), .Y(n30186) );
  OAI22X1 U17899 ( .A(n25318), .B(n30189), .C(n25328), .D(n30190), .Y(n30188)
         );
  OAI22X1 U17900 ( .A(n25339), .B(n30191), .C(n25349), .D(n30192), .Y(n30187)
         );
  AOI22X1 U17901 ( .A(reg_file[3468]), .B(n25360), .C(reg_file[3340]), .D(
        n25371), .Y(n30185) );
  AOI22X1 U17902 ( .A(reg_file[3212]), .B(n25381), .C(reg_file[3084]), .D(
        n25392), .Y(n30184) );
  NAND3X1 U17903 ( .A(n30193), .B(n30194), .C(n30195), .Y(n30182) );
  NOR2X1 U17904 ( .A(n30196), .B(n30197), .Y(n30195) );
  OAI22X1 U17905 ( .A(n25402), .B(n30198), .C(n25412), .D(n30199), .Y(n30197)
         );
  OAI22X1 U17906 ( .A(n25423), .B(n30200), .C(n25433), .D(n30201), .Y(n30196)
         );
  AOI22X1 U17907 ( .A(reg_file[2444]), .B(n25444), .C(reg_file[2316]), .D(
        n25455), .Y(n30194) );
  AOI22X1 U17908 ( .A(reg_file[2188]), .B(n25465), .C(reg_file[2060]), .D(
        n25476), .Y(n30193) );
  AOI21X1 U17909 ( .A(n30202), .B(n30203), .C(n25139), .Y(rd2data1040_127_) );
  NOR2X1 U17910 ( .A(n30204), .B(n30205), .Y(n30203) );
  NAND3X1 U17911 ( .A(n30206), .B(n30207), .C(n30208), .Y(n30205) );
  NOR2X1 U17912 ( .A(n30209), .B(n30210), .Y(n30208) );
  OAI22X1 U17913 ( .A(n25150), .B(n30211), .C(n25160), .D(n30212), .Y(n30210)
         );
  OAI22X1 U17914 ( .A(n25171), .B(n30213), .C(n25181), .D(n30214), .Y(n30209)
         );
  AOI22X1 U17915 ( .A(reg_file[1535]), .B(n25192), .C(reg_file[1407]), .D(
        n25203), .Y(n30207) );
  AOI22X1 U17916 ( .A(reg_file[1279]), .B(n25213), .C(reg_file[1151]), .D(
        n25224), .Y(n30206) );
  NAND3X1 U17917 ( .A(n30215), .B(n30216), .C(n30217), .Y(n30204) );
  NOR2X1 U17918 ( .A(n30218), .B(n30219), .Y(n30217) );
  OAI22X1 U17919 ( .A(n25234), .B(n30220), .C(n25244), .D(n30221), .Y(n30219)
         );
  OAI22X1 U17920 ( .A(n25255), .B(n30222), .C(n25265), .D(n30223), .Y(n30218)
         );
  AOI22X1 U17921 ( .A(reg_file[639]), .B(n25276), .C(reg_file[767]), .D(n25287), .Y(n30216) );
  AOI22X1 U17922 ( .A(reg_file[895]), .B(n25297), .C(reg_file[1023]), .D(
        n25308), .Y(n30215) );
  NOR2X1 U17923 ( .A(n30224), .B(n30225), .Y(n30202) );
  NAND3X1 U17924 ( .A(n30226), .B(n30227), .C(n30228), .Y(n30225) );
  NOR2X1 U17925 ( .A(n30229), .B(n30230), .Y(n30228) );
  OAI22X1 U17926 ( .A(n25318), .B(n30231), .C(n25328), .D(n30232), .Y(n30230)
         );
  OAI22X1 U17927 ( .A(n25339), .B(n30233), .C(n25349), .D(n30234), .Y(n30229)
         );
  AOI22X1 U17928 ( .A(reg_file[3583]), .B(n25360), .C(reg_file[3455]), .D(
        n25371), .Y(n30227) );
  AOI22X1 U17929 ( .A(reg_file[3327]), .B(n25381), .C(reg_file[3199]), .D(
        n25392), .Y(n30226) );
  NAND3X1 U17930 ( .A(n30235), .B(n30236), .C(n30237), .Y(n30224) );
  NOR2X1 U17931 ( .A(n30238), .B(n30239), .Y(n30237) );
  OAI22X1 U17932 ( .A(n25402), .B(n30240), .C(n25412), .D(n30241), .Y(n30239)
         );
  OAI22X1 U17933 ( .A(n25423), .B(n30242), .C(n25433), .D(n30243), .Y(n30238)
         );
  AOI22X1 U17934 ( .A(reg_file[2559]), .B(n25444), .C(reg_file[2431]), .D(
        n25455), .Y(n30236) );
  AOI22X1 U17935 ( .A(reg_file[2303]), .B(n25465), .C(reg_file[2175]), .D(
        n25476), .Y(n30235) );
  AOI21X1 U17936 ( .A(n30244), .B(n30245), .C(n25139), .Y(rd2data1040_126_) );
  NOR2X1 U17937 ( .A(n30246), .B(n30247), .Y(n30245) );
  NAND3X1 U17938 ( .A(n30248), .B(n30249), .C(n30250), .Y(n30247) );
  NOR2X1 U17939 ( .A(n30251), .B(n30252), .Y(n30250) );
  OAI22X1 U17940 ( .A(n25150), .B(n30253), .C(n25160), .D(n30254), .Y(n30252)
         );
  OAI22X1 U17941 ( .A(n25171), .B(n30255), .C(n25181), .D(n30256), .Y(n30251)
         );
  AOI22X1 U17942 ( .A(reg_file[1534]), .B(n25192), .C(reg_file[1406]), .D(
        n25203), .Y(n30249) );
  AOI22X1 U17943 ( .A(reg_file[1278]), .B(n25213), .C(reg_file[1150]), .D(
        n25224), .Y(n30248) );
  NAND3X1 U17944 ( .A(n30257), .B(n30258), .C(n30259), .Y(n30246) );
  NOR2X1 U17945 ( .A(n30260), .B(n30261), .Y(n30259) );
  OAI22X1 U17946 ( .A(n25234), .B(n30262), .C(n25244), .D(n30263), .Y(n30261)
         );
  OAI22X1 U17947 ( .A(n25255), .B(n30264), .C(n25265), .D(n30265), .Y(n30260)
         );
  AOI22X1 U17948 ( .A(reg_file[638]), .B(n25276), .C(reg_file[766]), .D(n25287), .Y(n30258) );
  AOI22X1 U17949 ( .A(reg_file[894]), .B(n25297), .C(reg_file[1022]), .D(
        n25308), .Y(n30257) );
  NOR2X1 U17950 ( .A(n30266), .B(n30267), .Y(n30244) );
  NAND3X1 U17951 ( .A(n30268), .B(n30269), .C(n30270), .Y(n30267) );
  NOR2X1 U17952 ( .A(n30271), .B(n30272), .Y(n30270) );
  OAI22X1 U17953 ( .A(n25318), .B(n30273), .C(n25328), .D(n30274), .Y(n30272)
         );
  OAI22X1 U17954 ( .A(n25339), .B(n30275), .C(n25349), .D(n30276), .Y(n30271)
         );
  AOI22X1 U17955 ( .A(reg_file[3582]), .B(n25360), .C(reg_file[3454]), .D(
        n25371), .Y(n30269) );
  AOI22X1 U17956 ( .A(reg_file[3326]), .B(n25381), .C(reg_file[3198]), .D(
        n25392), .Y(n30268) );
  NAND3X1 U17957 ( .A(n30277), .B(n30278), .C(n30279), .Y(n30266) );
  NOR2X1 U17958 ( .A(n30280), .B(n30281), .Y(n30279) );
  OAI22X1 U17959 ( .A(n25402), .B(n30282), .C(n25412), .D(n30283), .Y(n30281)
         );
  OAI22X1 U17960 ( .A(n25423), .B(n30284), .C(n25433), .D(n30285), .Y(n30280)
         );
  AOI22X1 U17961 ( .A(reg_file[2558]), .B(n25444), .C(reg_file[2430]), .D(
        n25455), .Y(n30278) );
  AOI22X1 U17962 ( .A(reg_file[2302]), .B(n25465), .C(reg_file[2174]), .D(
        n25476), .Y(n30277) );
  AOI21X1 U17963 ( .A(n30286), .B(n30287), .C(n25139), .Y(rd2data1040_125_) );
  NOR2X1 U17964 ( .A(n30288), .B(n30289), .Y(n30287) );
  NAND3X1 U17965 ( .A(n30290), .B(n30291), .C(n30292), .Y(n30289) );
  NOR2X1 U17966 ( .A(n30293), .B(n30294), .Y(n30292) );
  OAI22X1 U17967 ( .A(n25150), .B(n30295), .C(n25160), .D(n30296), .Y(n30294)
         );
  OAI22X1 U17968 ( .A(n25171), .B(n30297), .C(n25181), .D(n30298), .Y(n30293)
         );
  AOI22X1 U17969 ( .A(reg_file[1533]), .B(n25192), .C(reg_file[1405]), .D(
        n25203), .Y(n30291) );
  AOI22X1 U17970 ( .A(reg_file[1277]), .B(n25213), .C(reg_file[1149]), .D(
        n25224), .Y(n30290) );
  NAND3X1 U17971 ( .A(n30299), .B(n30300), .C(n30301), .Y(n30288) );
  NOR2X1 U17972 ( .A(n30302), .B(n30303), .Y(n30301) );
  OAI22X1 U17973 ( .A(n25234), .B(n30304), .C(n25244), .D(n30305), .Y(n30303)
         );
  OAI22X1 U17974 ( .A(n25255), .B(n30306), .C(n25265), .D(n30307), .Y(n30302)
         );
  AOI22X1 U17975 ( .A(reg_file[637]), .B(n25276), .C(reg_file[765]), .D(n25287), .Y(n30300) );
  AOI22X1 U17976 ( .A(reg_file[893]), .B(n25297), .C(reg_file[1021]), .D(
        n25308), .Y(n30299) );
  NOR2X1 U17977 ( .A(n30308), .B(n30309), .Y(n30286) );
  NAND3X1 U17978 ( .A(n30310), .B(n30311), .C(n30312), .Y(n30309) );
  NOR2X1 U17979 ( .A(n30313), .B(n30314), .Y(n30312) );
  OAI22X1 U17980 ( .A(n25318), .B(n30315), .C(n25328), .D(n30316), .Y(n30314)
         );
  OAI22X1 U17981 ( .A(n25339), .B(n30317), .C(n25349), .D(n30318), .Y(n30313)
         );
  AOI22X1 U17982 ( .A(reg_file[3581]), .B(n25360), .C(reg_file[3453]), .D(
        n25371), .Y(n30311) );
  AOI22X1 U17983 ( .A(reg_file[3325]), .B(n25381), .C(reg_file[3197]), .D(
        n25392), .Y(n30310) );
  NAND3X1 U17984 ( .A(n30319), .B(n30320), .C(n30321), .Y(n30308) );
  NOR2X1 U17985 ( .A(n30322), .B(n30323), .Y(n30321) );
  OAI22X1 U17986 ( .A(n25402), .B(n30324), .C(n25412), .D(n30325), .Y(n30323)
         );
  OAI22X1 U17987 ( .A(n25423), .B(n30326), .C(n25433), .D(n30327), .Y(n30322)
         );
  AOI22X1 U17988 ( .A(reg_file[2557]), .B(n25444), .C(reg_file[2429]), .D(
        n25455), .Y(n30320) );
  AOI22X1 U17989 ( .A(reg_file[2301]), .B(n25465), .C(reg_file[2173]), .D(
        n25476), .Y(n30319) );
  AOI21X1 U17990 ( .A(n30328), .B(n30329), .C(n25139), .Y(rd2data1040_124_) );
  NOR2X1 U17991 ( .A(n30330), .B(n30331), .Y(n30329) );
  NAND3X1 U17992 ( .A(n30332), .B(n30333), .C(n30334), .Y(n30331) );
  NOR2X1 U17993 ( .A(n30335), .B(n30336), .Y(n30334) );
  OAI22X1 U17994 ( .A(n25150), .B(n30337), .C(n25160), .D(n30338), .Y(n30336)
         );
  OAI22X1 U17995 ( .A(n25171), .B(n30339), .C(n25181), .D(n30340), .Y(n30335)
         );
  AOI22X1 U17996 ( .A(reg_file[1532]), .B(n25192), .C(reg_file[1404]), .D(
        n25203), .Y(n30333) );
  AOI22X1 U17997 ( .A(reg_file[1276]), .B(n25213), .C(reg_file[1148]), .D(
        n25224), .Y(n30332) );
  NAND3X1 U17998 ( .A(n30341), .B(n30342), .C(n30343), .Y(n30330) );
  NOR2X1 U17999 ( .A(n30344), .B(n30345), .Y(n30343) );
  OAI22X1 U18000 ( .A(n25234), .B(n30346), .C(n25244), .D(n30347), .Y(n30345)
         );
  OAI22X1 U18001 ( .A(n25255), .B(n30348), .C(n25265), .D(n30349), .Y(n30344)
         );
  AOI22X1 U18002 ( .A(reg_file[636]), .B(n25276), .C(reg_file[764]), .D(n25287), .Y(n30342) );
  AOI22X1 U18003 ( .A(reg_file[892]), .B(n25297), .C(reg_file[1020]), .D(
        n25308), .Y(n30341) );
  NOR2X1 U18004 ( .A(n30350), .B(n30351), .Y(n30328) );
  NAND3X1 U18005 ( .A(n30352), .B(n30353), .C(n30354), .Y(n30351) );
  NOR2X1 U18006 ( .A(n30355), .B(n30356), .Y(n30354) );
  OAI22X1 U18007 ( .A(n25318), .B(n30357), .C(n25328), .D(n30358), .Y(n30356)
         );
  OAI22X1 U18008 ( .A(n25339), .B(n30359), .C(n25349), .D(n30360), .Y(n30355)
         );
  AOI22X1 U18009 ( .A(reg_file[3580]), .B(n25360), .C(reg_file[3452]), .D(
        n25371), .Y(n30353) );
  AOI22X1 U18010 ( .A(reg_file[3324]), .B(n25381), .C(reg_file[3196]), .D(
        n25392), .Y(n30352) );
  NAND3X1 U18011 ( .A(n30361), .B(n30362), .C(n30363), .Y(n30350) );
  NOR2X1 U18012 ( .A(n30364), .B(n30365), .Y(n30363) );
  OAI22X1 U18013 ( .A(n25402), .B(n30366), .C(n25412), .D(n30367), .Y(n30365)
         );
  OAI22X1 U18014 ( .A(n25423), .B(n30368), .C(n25433), .D(n30369), .Y(n30364)
         );
  AOI22X1 U18015 ( .A(reg_file[2556]), .B(n25444), .C(reg_file[2428]), .D(
        n25455), .Y(n30362) );
  AOI22X1 U18016 ( .A(reg_file[2300]), .B(n25465), .C(reg_file[2172]), .D(
        n25476), .Y(n30361) );
  AOI21X1 U18017 ( .A(n30370), .B(n30371), .C(n25139), .Y(rd2data1040_123_) );
  NOR2X1 U18018 ( .A(n30372), .B(n30373), .Y(n30371) );
  NAND3X1 U18019 ( .A(n30374), .B(n30375), .C(n30376), .Y(n30373) );
  NOR2X1 U18020 ( .A(n30377), .B(n30378), .Y(n30376) );
  OAI22X1 U18021 ( .A(n25150), .B(n30379), .C(n25160), .D(n30380), .Y(n30378)
         );
  OAI22X1 U18022 ( .A(n25171), .B(n30381), .C(n25181), .D(n30382), .Y(n30377)
         );
  AOI22X1 U18023 ( .A(reg_file[1531]), .B(n25192), .C(reg_file[1403]), .D(
        n25203), .Y(n30375) );
  AOI22X1 U18024 ( .A(reg_file[1275]), .B(n25213), .C(reg_file[1147]), .D(
        n25224), .Y(n30374) );
  NAND3X1 U18025 ( .A(n30383), .B(n30384), .C(n30385), .Y(n30372) );
  NOR2X1 U18026 ( .A(n30386), .B(n30387), .Y(n30385) );
  OAI22X1 U18027 ( .A(n25234), .B(n30388), .C(n25244), .D(n30389), .Y(n30387)
         );
  OAI22X1 U18028 ( .A(n25255), .B(n30390), .C(n25265), .D(n30391), .Y(n30386)
         );
  AOI22X1 U18029 ( .A(reg_file[635]), .B(n25276), .C(reg_file[763]), .D(n25287), .Y(n30384) );
  AOI22X1 U18030 ( .A(reg_file[891]), .B(n25297), .C(reg_file[1019]), .D(
        n25308), .Y(n30383) );
  NOR2X1 U18031 ( .A(n30392), .B(n30393), .Y(n30370) );
  NAND3X1 U18032 ( .A(n30394), .B(n30395), .C(n30396), .Y(n30393) );
  NOR2X1 U18033 ( .A(n30397), .B(n30398), .Y(n30396) );
  OAI22X1 U18034 ( .A(n25318), .B(n30399), .C(n25328), .D(n30400), .Y(n30398)
         );
  OAI22X1 U18035 ( .A(n25339), .B(n30401), .C(n25349), .D(n30402), .Y(n30397)
         );
  AOI22X1 U18036 ( .A(reg_file[3579]), .B(n25360), .C(reg_file[3451]), .D(
        n25371), .Y(n30395) );
  AOI22X1 U18037 ( .A(reg_file[3323]), .B(n25381), .C(reg_file[3195]), .D(
        n25392), .Y(n30394) );
  NAND3X1 U18038 ( .A(n30403), .B(n30404), .C(n30405), .Y(n30392) );
  NOR2X1 U18039 ( .A(n30406), .B(n30407), .Y(n30405) );
  OAI22X1 U18040 ( .A(n25402), .B(n30408), .C(n25412), .D(n30409), .Y(n30407)
         );
  OAI22X1 U18041 ( .A(n25423), .B(n30410), .C(n25433), .D(n30411), .Y(n30406)
         );
  AOI22X1 U18042 ( .A(reg_file[2555]), .B(n25444), .C(reg_file[2427]), .D(
        n25455), .Y(n30404) );
  AOI22X1 U18043 ( .A(reg_file[2299]), .B(n25465), .C(reg_file[2171]), .D(
        n25476), .Y(n30403) );
  AOI21X1 U18044 ( .A(n30412), .B(n30413), .C(n25139), .Y(rd2data1040_122_) );
  NOR2X1 U18045 ( .A(n30414), .B(n30415), .Y(n30413) );
  NAND3X1 U18046 ( .A(n30416), .B(n30417), .C(n30418), .Y(n30415) );
  NOR2X1 U18047 ( .A(n30419), .B(n30420), .Y(n30418) );
  OAI22X1 U18048 ( .A(n25149), .B(n30421), .C(n25160), .D(n30422), .Y(n30420)
         );
  OAI22X1 U18049 ( .A(n25170), .B(n30423), .C(n25181), .D(n30424), .Y(n30419)
         );
  AOI22X1 U18050 ( .A(reg_file[1530]), .B(n25192), .C(reg_file[1402]), .D(
        n25202), .Y(n30417) );
  AOI22X1 U18051 ( .A(reg_file[1274]), .B(n25213), .C(reg_file[1146]), .D(
        n25223), .Y(n30416) );
  NAND3X1 U18052 ( .A(n30425), .B(n30426), .C(n30427), .Y(n30414) );
  NOR2X1 U18053 ( .A(n30428), .B(n30429), .Y(n30427) );
  OAI22X1 U18054 ( .A(n25233), .B(n30430), .C(n25244), .D(n30431), .Y(n30429)
         );
  OAI22X1 U18055 ( .A(n25254), .B(n30432), .C(n25265), .D(n30433), .Y(n30428)
         );
  AOI22X1 U18056 ( .A(reg_file[634]), .B(n25276), .C(reg_file[762]), .D(n25286), .Y(n30426) );
  AOI22X1 U18057 ( .A(reg_file[890]), .B(n25297), .C(reg_file[1018]), .D(
        n25307), .Y(n30425) );
  NOR2X1 U18058 ( .A(n30434), .B(n30435), .Y(n30412) );
  NAND3X1 U18059 ( .A(n30436), .B(n30437), .C(n30438), .Y(n30435) );
  NOR2X1 U18060 ( .A(n30439), .B(n30440), .Y(n30438) );
  OAI22X1 U18061 ( .A(n25317), .B(n30441), .C(n25328), .D(n30442), .Y(n30440)
         );
  OAI22X1 U18062 ( .A(n25338), .B(n30443), .C(n25349), .D(n30444), .Y(n30439)
         );
  AOI22X1 U18063 ( .A(reg_file[3578]), .B(n25360), .C(reg_file[3450]), .D(
        n25370), .Y(n30437) );
  AOI22X1 U18064 ( .A(reg_file[3322]), .B(n25381), .C(reg_file[3194]), .D(
        n25391), .Y(n30436) );
  NAND3X1 U18065 ( .A(n30445), .B(n30446), .C(n30447), .Y(n30434) );
  NOR2X1 U18066 ( .A(n30448), .B(n30449), .Y(n30447) );
  OAI22X1 U18067 ( .A(n25401), .B(n30450), .C(n25412), .D(n30451), .Y(n30449)
         );
  OAI22X1 U18068 ( .A(n25422), .B(n30452), .C(n25433), .D(n30453), .Y(n30448)
         );
  AOI22X1 U18069 ( .A(reg_file[2554]), .B(n25444), .C(reg_file[2426]), .D(
        n25454), .Y(n30446) );
  AOI22X1 U18070 ( .A(reg_file[2298]), .B(n25465), .C(reg_file[2170]), .D(
        n25475), .Y(n30445) );
  AOI21X1 U18071 ( .A(n30454), .B(n30455), .C(n25139), .Y(rd2data1040_121_) );
  NOR2X1 U18072 ( .A(n30456), .B(n30457), .Y(n30455) );
  NAND3X1 U18073 ( .A(n30458), .B(n30459), .C(n30460), .Y(n30457) );
  NOR2X1 U18074 ( .A(n30461), .B(n30462), .Y(n30460) );
  OAI22X1 U18075 ( .A(n25149), .B(n30463), .C(n25160), .D(n30464), .Y(n30462)
         );
  OAI22X1 U18076 ( .A(n25170), .B(n30465), .C(n25181), .D(n30466), .Y(n30461)
         );
  AOI22X1 U18077 ( .A(reg_file[1529]), .B(n25192), .C(reg_file[1401]), .D(
        n25202), .Y(n30459) );
  AOI22X1 U18078 ( .A(reg_file[1273]), .B(n25213), .C(reg_file[1145]), .D(
        n25223), .Y(n30458) );
  NAND3X1 U18079 ( .A(n30467), .B(n30468), .C(n30469), .Y(n30456) );
  NOR2X1 U18080 ( .A(n30470), .B(n30471), .Y(n30469) );
  OAI22X1 U18081 ( .A(n25233), .B(n30472), .C(n25244), .D(n30473), .Y(n30471)
         );
  OAI22X1 U18082 ( .A(n25254), .B(n30474), .C(n25265), .D(n30475), .Y(n30470)
         );
  AOI22X1 U18083 ( .A(reg_file[633]), .B(n25276), .C(reg_file[761]), .D(n25286), .Y(n30468) );
  AOI22X1 U18084 ( .A(reg_file[889]), .B(n25297), .C(reg_file[1017]), .D(
        n25307), .Y(n30467) );
  NOR2X1 U18085 ( .A(n30476), .B(n30477), .Y(n30454) );
  NAND3X1 U18086 ( .A(n30478), .B(n30479), .C(n30480), .Y(n30477) );
  NOR2X1 U18087 ( .A(n30481), .B(n30482), .Y(n30480) );
  OAI22X1 U18088 ( .A(n25317), .B(n30483), .C(n25328), .D(n30484), .Y(n30482)
         );
  OAI22X1 U18089 ( .A(n25338), .B(n30485), .C(n25349), .D(n30486), .Y(n30481)
         );
  AOI22X1 U18090 ( .A(reg_file[3577]), .B(n25360), .C(reg_file[3449]), .D(
        n25370), .Y(n30479) );
  AOI22X1 U18091 ( .A(reg_file[3321]), .B(n25381), .C(reg_file[3193]), .D(
        n25391), .Y(n30478) );
  NAND3X1 U18092 ( .A(n30487), .B(n30488), .C(n30489), .Y(n30476) );
  NOR2X1 U18093 ( .A(n30490), .B(n30491), .Y(n30489) );
  OAI22X1 U18094 ( .A(n25401), .B(n30492), .C(n25412), .D(n30493), .Y(n30491)
         );
  OAI22X1 U18095 ( .A(n25422), .B(n30494), .C(n25433), .D(n30495), .Y(n30490)
         );
  AOI22X1 U18096 ( .A(reg_file[2553]), .B(n25444), .C(reg_file[2425]), .D(
        n25454), .Y(n30488) );
  AOI22X1 U18097 ( .A(reg_file[2297]), .B(n25465), .C(reg_file[2169]), .D(
        n25475), .Y(n30487) );
  AOI21X1 U18098 ( .A(n30496), .B(n30497), .C(n25138), .Y(rd2data1040_120_) );
  NOR2X1 U18099 ( .A(n30498), .B(n30499), .Y(n30497) );
  NAND3X1 U18100 ( .A(n30500), .B(n30501), .C(n30502), .Y(n30499) );
  NOR2X1 U18101 ( .A(n30503), .B(n30504), .Y(n30502) );
  OAI22X1 U18102 ( .A(n25149), .B(n30505), .C(n25159), .D(n30506), .Y(n30504)
         );
  OAI22X1 U18103 ( .A(n25170), .B(n30507), .C(n25180), .D(n30508), .Y(n30503)
         );
  AOI22X1 U18104 ( .A(reg_file[1528]), .B(n25191), .C(reg_file[1400]), .D(
        n25202), .Y(n30501) );
  AOI22X1 U18105 ( .A(reg_file[1272]), .B(n25212), .C(reg_file[1144]), .D(
        n25223), .Y(n30500) );
  NAND3X1 U18106 ( .A(n30509), .B(n30510), .C(n30511), .Y(n30498) );
  NOR2X1 U18107 ( .A(n30512), .B(n30513), .Y(n30511) );
  OAI22X1 U18108 ( .A(n25233), .B(n30514), .C(n25243), .D(n30515), .Y(n30513)
         );
  OAI22X1 U18109 ( .A(n25254), .B(n30516), .C(n25264), .D(n30517), .Y(n30512)
         );
  AOI22X1 U18110 ( .A(reg_file[632]), .B(n25275), .C(reg_file[760]), .D(n25286), .Y(n30510) );
  AOI22X1 U18111 ( .A(reg_file[888]), .B(n25296), .C(reg_file[1016]), .D(
        n25307), .Y(n30509) );
  NOR2X1 U18112 ( .A(n30518), .B(n30519), .Y(n30496) );
  NAND3X1 U18113 ( .A(n30520), .B(n30521), .C(n30522), .Y(n30519) );
  NOR2X1 U18114 ( .A(n30523), .B(n30524), .Y(n30522) );
  OAI22X1 U18115 ( .A(n25317), .B(n30525), .C(n25327), .D(n30526), .Y(n30524)
         );
  OAI22X1 U18116 ( .A(n25338), .B(n30527), .C(n25348), .D(n30528), .Y(n30523)
         );
  AOI22X1 U18117 ( .A(reg_file[3576]), .B(n25359), .C(reg_file[3448]), .D(
        n25370), .Y(n30521) );
  AOI22X1 U18118 ( .A(reg_file[3320]), .B(n25380), .C(reg_file[3192]), .D(
        n25391), .Y(n30520) );
  NAND3X1 U18119 ( .A(n30529), .B(n30530), .C(n30531), .Y(n30518) );
  NOR2X1 U18120 ( .A(n30532), .B(n30533), .Y(n30531) );
  OAI22X1 U18121 ( .A(n25401), .B(n30534), .C(n25411), .D(n30535), .Y(n30533)
         );
  OAI22X1 U18122 ( .A(n25422), .B(n30536), .C(n25432), .D(n30537), .Y(n30532)
         );
  AOI22X1 U18123 ( .A(reg_file[2552]), .B(n25443), .C(reg_file[2424]), .D(
        n25454), .Y(n30530) );
  AOI22X1 U18124 ( .A(reg_file[2296]), .B(n25464), .C(reg_file[2168]), .D(
        n25475), .Y(n30529) );
  AOI21X1 U18125 ( .A(n30538), .B(n30539), .C(n25138), .Y(rd2data1040_11_) );
  NOR2X1 U18126 ( .A(n30540), .B(n30541), .Y(n30539) );
  NAND3X1 U18127 ( .A(n30542), .B(n30543), .C(n30544), .Y(n30541) );
  NOR2X1 U18128 ( .A(n30545), .B(n30546), .Y(n30544) );
  OAI22X1 U18129 ( .A(n25149), .B(n30547), .C(n25159), .D(n30548), .Y(n30546)
         );
  OAI22X1 U18130 ( .A(n25170), .B(n30549), .C(n25180), .D(n30550), .Y(n30545)
         );
  AOI22X1 U18131 ( .A(reg_file[1419]), .B(n25191), .C(reg_file[1291]), .D(
        n25202), .Y(n30543) );
  AOI22X1 U18132 ( .A(reg_file[1163]), .B(n25212), .C(reg_file[1035]), .D(
        n25223), .Y(n30542) );
  NAND3X1 U18133 ( .A(n30551), .B(n30552), .C(n30553), .Y(n30540) );
  NOR2X1 U18134 ( .A(n30554), .B(n30555), .Y(n30553) );
  OAI22X1 U18135 ( .A(n25233), .B(n30556), .C(n25243), .D(n30557), .Y(n30555)
         );
  OAI22X1 U18136 ( .A(n25254), .B(n30558), .C(n25264), .D(n30559), .Y(n30554)
         );
  AOI22X1 U18137 ( .A(reg_file[523]), .B(n25275), .C(reg_file[651]), .D(n25286), .Y(n30552) );
  AOI22X1 U18138 ( .A(reg_file[779]), .B(n25296), .C(reg_file[907]), .D(n25307), .Y(n30551) );
  NOR2X1 U18139 ( .A(n30560), .B(n30561), .Y(n30538) );
  NAND3X1 U18140 ( .A(n30562), .B(n30563), .C(n30564), .Y(n30561) );
  NOR2X1 U18141 ( .A(n30565), .B(n30566), .Y(n30564) );
  OAI22X1 U18142 ( .A(n25317), .B(n30567), .C(n25327), .D(n30568), .Y(n30566)
         );
  OAI22X1 U18143 ( .A(n25338), .B(n30569), .C(n25348), .D(n30570), .Y(n30565)
         );
  AOI22X1 U18144 ( .A(reg_file[3467]), .B(n25359), .C(reg_file[3339]), .D(
        n25370), .Y(n30563) );
  AOI22X1 U18145 ( .A(reg_file[3211]), .B(n25380), .C(reg_file[3083]), .D(
        n25391), .Y(n30562) );
  NAND3X1 U18146 ( .A(n30571), .B(n30572), .C(n30573), .Y(n30560) );
  NOR2X1 U18147 ( .A(n30574), .B(n30575), .Y(n30573) );
  OAI22X1 U18148 ( .A(n25401), .B(n30576), .C(n25411), .D(n30577), .Y(n30575)
         );
  OAI22X1 U18149 ( .A(n25422), .B(n30578), .C(n25432), .D(n30579), .Y(n30574)
         );
  AOI22X1 U18150 ( .A(reg_file[2443]), .B(n25443), .C(reg_file[2315]), .D(
        n25454), .Y(n30572) );
  AOI22X1 U18151 ( .A(reg_file[2187]), .B(n25464), .C(reg_file[2059]), .D(
        n25475), .Y(n30571) );
  AOI21X1 U18152 ( .A(n30580), .B(n30581), .C(n25138), .Y(rd2data1040_119_) );
  NOR2X1 U18153 ( .A(n30582), .B(n30583), .Y(n30581) );
  NAND3X1 U18154 ( .A(n30584), .B(n30585), .C(n30586), .Y(n30583) );
  NOR2X1 U18155 ( .A(n30587), .B(n30588), .Y(n30586) );
  OAI22X1 U18156 ( .A(n25149), .B(n30589), .C(n25159), .D(n30590), .Y(n30588)
         );
  OAI22X1 U18157 ( .A(n25170), .B(n30591), .C(n25180), .D(n30592), .Y(n30587)
         );
  AOI22X1 U18158 ( .A(reg_file[1527]), .B(n25191), .C(reg_file[1399]), .D(
        n25202), .Y(n30585) );
  AOI22X1 U18159 ( .A(reg_file[1271]), .B(n25212), .C(reg_file[1143]), .D(
        n25223), .Y(n30584) );
  NAND3X1 U18160 ( .A(n30593), .B(n30594), .C(n30595), .Y(n30582) );
  NOR2X1 U18161 ( .A(n30596), .B(n30597), .Y(n30595) );
  OAI22X1 U18162 ( .A(n25233), .B(n30598), .C(n25243), .D(n30599), .Y(n30597)
         );
  OAI22X1 U18163 ( .A(n25254), .B(n30600), .C(n25264), .D(n30601), .Y(n30596)
         );
  AOI22X1 U18164 ( .A(reg_file[631]), .B(n25275), .C(reg_file[759]), .D(n25286), .Y(n30594) );
  AOI22X1 U18165 ( .A(reg_file[887]), .B(n25296), .C(reg_file[1015]), .D(
        n25307), .Y(n30593) );
  NOR2X1 U18166 ( .A(n30602), .B(n30603), .Y(n30580) );
  NAND3X1 U18167 ( .A(n30604), .B(n30605), .C(n30606), .Y(n30603) );
  NOR2X1 U18168 ( .A(n30607), .B(n30608), .Y(n30606) );
  OAI22X1 U18169 ( .A(n25317), .B(n30609), .C(n25327), .D(n30610), .Y(n30608)
         );
  OAI22X1 U18170 ( .A(n25338), .B(n30611), .C(n25348), .D(n30612), .Y(n30607)
         );
  AOI22X1 U18171 ( .A(reg_file[3575]), .B(n25359), .C(reg_file[3447]), .D(
        n25370), .Y(n30605) );
  AOI22X1 U18172 ( .A(reg_file[3319]), .B(n25380), .C(reg_file[3191]), .D(
        n25391), .Y(n30604) );
  NAND3X1 U18173 ( .A(n30613), .B(n30614), .C(n30615), .Y(n30602) );
  NOR2X1 U18174 ( .A(n30616), .B(n30617), .Y(n30615) );
  OAI22X1 U18175 ( .A(n25401), .B(n30618), .C(n25411), .D(n30619), .Y(n30617)
         );
  OAI22X1 U18176 ( .A(n25422), .B(n30620), .C(n25432), .D(n30621), .Y(n30616)
         );
  AOI22X1 U18177 ( .A(reg_file[2551]), .B(n25443), .C(reg_file[2423]), .D(
        n25454), .Y(n30614) );
  AOI22X1 U18178 ( .A(reg_file[2295]), .B(n25464), .C(reg_file[2167]), .D(
        n25475), .Y(n30613) );
  AOI21X1 U18179 ( .A(n30622), .B(n30623), .C(n25138), .Y(rd2data1040_118_) );
  NOR2X1 U18180 ( .A(n30624), .B(n30625), .Y(n30623) );
  NAND3X1 U18181 ( .A(n30626), .B(n30627), .C(n30628), .Y(n30625) );
  NOR2X1 U18182 ( .A(n30629), .B(n30630), .Y(n30628) );
  OAI22X1 U18183 ( .A(n25149), .B(n30631), .C(n25159), .D(n30632), .Y(n30630)
         );
  OAI22X1 U18184 ( .A(n25170), .B(n30633), .C(n25180), .D(n30634), .Y(n30629)
         );
  AOI22X1 U18185 ( .A(reg_file[1526]), .B(n25191), .C(reg_file[1398]), .D(
        n25202), .Y(n30627) );
  AOI22X1 U18186 ( .A(reg_file[1270]), .B(n25212), .C(reg_file[1142]), .D(
        n25223), .Y(n30626) );
  NAND3X1 U18187 ( .A(n30635), .B(n30636), .C(n30637), .Y(n30624) );
  NOR2X1 U18188 ( .A(n30638), .B(n30639), .Y(n30637) );
  OAI22X1 U18189 ( .A(n25233), .B(n30640), .C(n25243), .D(n30641), .Y(n30639)
         );
  OAI22X1 U18190 ( .A(n25254), .B(n30642), .C(n25264), .D(n30643), .Y(n30638)
         );
  AOI22X1 U18191 ( .A(reg_file[630]), .B(n25275), .C(reg_file[758]), .D(n25286), .Y(n30636) );
  AOI22X1 U18192 ( .A(reg_file[886]), .B(n25296), .C(reg_file[1014]), .D(
        n25307), .Y(n30635) );
  NOR2X1 U18193 ( .A(n30644), .B(n30645), .Y(n30622) );
  NAND3X1 U18194 ( .A(n30646), .B(n30647), .C(n30648), .Y(n30645) );
  NOR2X1 U18195 ( .A(n30649), .B(n30650), .Y(n30648) );
  OAI22X1 U18196 ( .A(n25317), .B(n30651), .C(n25327), .D(n30652), .Y(n30650)
         );
  OAI22X1 U18197 ( .A(n25338), .B(n30653), .C(n25348), .D(n30654), .Y(n30649)
         );
  AOI22X1 U18198 ( .A(reg_file[3574]), .B(n25359), .C(reg_file[3446]), .D(
        n25370), .Y(n30647) );
  AOI22X1 U18199 ( .A(reg_file[3318]), .B(n25380), .C(reg_file[3190]), .D(
        n25391), .Y(n30646) );
  NAND3X1 U18200 ( .A(n30655), .B(n30656), .C(n30657), .Y(n30644) );
  NOR2X1 U18201 ( .A(n30658), .B(n30659), .Y(n30657) );
  OAI22X1 U18202 ( .A(n25401), .B(n30660), .C(n25411), .D(n30661), .Y(n30659)
         );
  OAI22X1 U18203 ( .A(n25422), .B(n30662), .C(n25432), .D(n30663), .Y(n30658)
         );
  AOI22X1 U18204 ( .A(reg_file[2550]), .B(n25443), .C(reg_file[2422]), .D(
        n25454), .Y(n30656) );
  AOI22X1 U18205 ( .A(reg_file[2294]), .B(n25464), .C(reg_file[2166]), .D(
        n25475), .Y(n30655) );
  AOI21X1 U18206 ( .A(n30664), .B(n30665), .C(n25138), .Y(rd2data1040_117_) );
  NOR2X1 U18207 ( .A(n30666), .B(n30667), .Y(n30665) );
  NAND3X1 U18208 ( .A(n30668), .B(n30669), .C(n30670), .Y(n30667) );
  NOR2X1 U18209 ( .A(n30671), .B(n30672), .Y(n30670) );
  OAI22X1 U18210 ( .A(n25149), .B(n30673), .C(n25159), .D(n30674), .Y(n30672)
         );
  OAI22X1 U18211 ( .A(n25170), .B(n30675), .C(n25180), .D(n30676), .Y(n30671)
         );
  AOI22X1 U18212 ( .A(reg_file[1525]), .B(n25191), .C(reg_file[1397]), .D(
        n25202), .Y(n30669) );
  AOI22X1 U18213 ( .A(reg_file[1269]), .B(n25212), .C(reg_file[1141]), .D(
        n25223), .Y(n30668) );
  NAND3X1 U18214 ( .A(n30677), .B(n30678), .C(n30679), .Y(n30666) );
  NOR2X1 U18215 ( .A(n30680), .B(n30681), .Y(n30679) );
  OAI22X1 U18216 ( .A(n25233), .B(n30682), .C(n25243), .D(n30683), .Y(n30681)
         );
  OAI22X1 U18217 ( .A(n25254), .B(n30684), .C(n25264), .D(n30685), .Y(n30680)
         );
  AOI22X1 U18218 ( .A(reg_file[629]), .B(n25275), .C(reg_file[757]), .D(n25286), .Y(n30678) );
  AOI22X1 U18219 ( .A(reg_file[885]), .B(n25296), .C(reg_file[1013]), .D(
        n25307), .Y(n30677) );
  NOR2X1 U18220 ( .A(n30686), .B(n30687), .Y(n30664) );
  NAND3X1 U18221 ( .A(n30688), .B(n30689), .C(n30690), .Y(n30687) );
  NOR2X1 U18222 ( .A(n30691), .B(n30692), .Y(n30690) );
  OAI22X1 U18223 ( .A(n25317), .B(n30693), .C(n25327), .D(n30694), .Y(n30692)
         );
  OAI22X1 U18224 ( .A(n25338), .B(n30695), .C(n25348), .D(n30696), .Y(n30691)
         );
  AOI22X1 U18225 ( .A(reg_file[3573]), .B(n25359), .C(reg_file[3445]), .D(
        n25370), .Y(n30689) );
  AOI22X1 U18226 ( .A(reg_file[3317]), .B(n25380), .C(reg_file[3189]), .D(
        n25391), .Y(n30688) );
  NAND3X1 U18227 ( .A(n30697), .B(n30698), .C(n30699), .Y(n30686) );
  NOR2X1 U18228 ( .A(n30700), .B(n30701), .Y(n30699) );
  OAI22X1 U18229 ( .A(n25401), .B(n30702), .C(n25411), .D(n30703), .Y(n30701)
         );
  OAI22X1 U18230 ( .A(n25422), .B(n30704), .C(n25432), .D(n30705), .Y(n30700)
         );
  AOI22X1 U18231 ( .A(reg_file[2549]), .B(n25443), .C(reg_file[2421]), .D(
        n25454), .Y(n30698) );
  AOI22X1 U18232 ( .A(reg_file[2293]), .B(n25464), .C(reg_file[2165]), .D(
        n25475), .Y(n30697) );
  AOI21X1 U18233 ( .A(n30706), .B(n30707), .C(n25138), .Y(rd2data1040_116_) );
  NOR2X1 U18234 ( .A(n30708), .B(n30709), .Y(n30707) );
  NAND3X1 U18235 ( .A(n30710), .B(n30711), .C(n30712), .Y(n30709) );
  NOR2X1 U18236 ( .A(n30713), .B(n30714), .Y(n30712) );
  OAI22X1 U18237 ( .A(n25149), .B(n30715), .C(n25159), .D(n30716), .Y(n30714)
         );
  OAI22X1 U18238 ( .A(n25170), .B(n30717), .C(n25180), .D(n30718), .Y(n30713)
         );
  AOI22X1 U18239 ( .A(reg_file[1524]), .B(n25191), .C(reg_file[1396]), .D(
        n25202), .Y(n30711) );
  AOI22X1 U18240 ( .A(reg_file[1268]), .B(n25212), .C(reg_file[1140]), .D(
        n25223), .Y(n30710) );
  NAND3X1 U18241 ( .A(n30719), .B(n30720), .C(n30721), .Y(n30708) );
  NOR2X1 U18242 ( .A(n30722), .B(n30723), .Y(n30721) );
  OAI22X1 U18243 ( .A(n25233), .B(n30724), .C(n25243), .D(n30725), .Y(n30723)
         );
  OAI22X1 U18244 ( .A(n25254), .B(n30726), .C(n25264), .D(n30727), .Y(n30722)
         );
  AOI22X1 U18245 ( .A(reg_file[628]), .B(n25275), .C(reg_file[756]), .D(n25286), .Y(n30720) );
  AOI22X1 U18246 ( .A(reg_file[884]), .B(n25296), .C(reg_file[1012]), .D(
        n25307), .Y(n30719) );
  NOR2X1 U18247 ( .A(n30728), .B(n30729), .Y(n30706) );
  NAND3X1 U18248 ( .A(n30730), .B(n30731), .C(n30732), .Y(n30729) );
  NOR2X1 U18249 ( .A(n30733), .B(n30734), .Y(n30732) );
  OAI22X1 U18250 ( .A(n25317), .B(n30735), .C(n25327), .D(n30736), .Y(n30734)
         );
  OAI22X1 U18251 ( .A(n25338), .B(n30737), .C(n25348), .D(n30738), .Y(n30733)
         );
  AOI22X1 U18252 ( .A(reg_file[3572]), .B(n25359), .C(reg_file[3444]), .D(
        n25370), .Y(n30731) );
  AOI22X1 U18253 ( .A(reg_file[3316]), .B(n25380), .C(reg_file[3188]), .D(
        n25391), .Y(n30730) );
  NAND3X1 U18254 ( .A(n30739), .B(n30740), .C(n30741), .Y(n30728) );
  NOR2X1 U18255 ( .A(n30742), .B(n30743), .Y(n30741) );
  OAI22X1 U18256 ( .A(n25401), .B(n30744), .C(n25411), .D(n30745), .Y(n30743)
         );
  OAI22X1 U18257 ( .A(n25422), .B(n30746), .C(n25432), .D(n30747), .Y(n30742)
         );
  AOI22X1 U18258 ( .A(reg_file[2548]), .B(n25443), .C(reg_file[2420]), .D(
        n25454), .Y(n30740) );
  AOI22X1 U18259 ( .A(reg_file[2292]), .B(n25464), .C(reg_file[2164]), .D(
        n25475), .Y(n30739) );
  AOI21X1 U18260 ( .A(n30748), .B(n30749), .C(n25138), .Y(rd2data1040_115_) );
  NOR2X1 U18261 ( .A(n30750), .B(n30751), .Y(n30749) );
  NAND3X1 U18262 ( .A(n30752), .B(n30753), .C(n30754), .Y(n30751) );
  NOR2X1 U18263 ( .A(n30755), .B(n30756), .Y(n30754) );
  OAI22X1 U18264 ( .A(n25149), .B(n30757), .C(n25159), .D(n30758), .Y(n30756)
         );
  OAI22X1 U18265 ( .A(n25170), .B(n30759), .C(n25180), .D(n30760), .Y(n30755)
         );
  AOI22X1 U18266 ( .A(reg_file[1523]), .B(n25191), .C(reg_file[1395]), .D(
        n25202), .Y(n30753) );
  AOI22X1 U18267 ( .A(reg_file[1267]), .B(n25212), .C(reg_file[1139]), .D(
        n25223), .Y(n30752) );
  NAND3X1 U18268 ( .A(n30761), .B(n30762), .C(n30763), .Y(n30750) );
  NOR2X1 U18269 ( .A(n30764), .B(n30765), .Y(n30763) );
  OAI22X1 U18270 ( .A(n25233), .B(n30766), .C(n25243), .D(n30767), .Y(n30765)
         );
  OAI22X1 U18271 ( .A(n25254), .B(n30768), .C(n25264), .D(n30769), .Y(n30764)
         );
  AOI22X1 U18272 ( .A(reg_file[627]), .B(n25275), .C(reg_file[755]), .D(n25286), .Y(n30762) );
  AOI22X1 U18273 ( .A(reg_file[883]), .B(n25296), .C(reg_file[1011]), .D(
        n25307), .Y(n30761) );
  NOR2X1 U18274 ( .A(n30770), .B(n30771), .Y(n30748) );
  NAND3X1 U18275 ( .A(n30772), .B(n30773), .C(n30774), .Y(n30771) );
  NOR2X1 U18276 ( .A(n30775), .B(n30776), .Y(n30774) );
  OAI22X1 U18277 ( .A(n25317), .B(n30777), .C(n25327), .D(n30778), .Y(n30776)
         );
  OAI22X1 U18278 ( .A(n25338), .B(n30779), .C(n25348), .D(n30780), .Y(n30775)
         );
  AOI22X1 U18279 ( .A(reg_file[3571]), .B(n25359), .C(reg_file[3443]), .D(
        n25370), .Y(n30773) );
  AOI22X1 U18280 ( .A(reg_file[3315]), .B(n25380), .C(reg_file[3187]), .D(
        n25391), .Y(n30772) );
  NAND3X1 U18281 ( .A(n30781), .B(n30782), .C(n30783), .Y(n30770) );
  NOR2X1 U18282 ( .A(n30784), .B(n30785), .Y(n30783) );
  OAI22X1 U18283 ( .A(n25401), .B(n30786), .C(n25411), .D(n30787), .Y(n30785)
         );
  OAI22X1 U18284 ( .A(n25422), .B(n30788), .C(n25432), .D(n30789), .Y(n30784)
         );
  AOI22X1 U18285 ( .A(reg_file[2547]), .B(n25443), .C(reg_file[2419]), .D(
        n25454), .Y(n30782) );
  AOI22X1 U18286 ( .A(reg_file[2291]), .B(n25464), .C(reg_file[2163]), .D(
        n25475), .Y(n30781) );
  AOI21X1 U18287 ( .A(n30790), .B(n30791), .C(n25138), .Y(rd2data1040_114_) );
  NOR2X1 U18288 ( .A(n30792), .B(n30793), .Y(n30791) );
  NAND3X1 U18289 ( .A(n30794), .B(n30795), .C(n30796), .Y(n30793) );
  NOR2X1 U18290 ( .A(n30797), .B(n30798), .Y(n30796) );
  OAI22X1 U18291 ( .A(n25149), .B(n30799), .C(n25159), .D(n30800), .Y(n30798)
         );
  OAI22X1 U18292 ( .A(n25170), .B(n30801), .C(n25180), .D(n30802), .Y(n30797)
         );
  AOI22X1 U18293 ( .A(reg_file[1522]), .B(n25191), .C(reg_file[1394]), .D(
        n25202), .Y(n30795) );
  AOI22X1 U18294 ( .A(reg_file[1266]), .B(n25212), .C(reg_file[1138]), .D(
        n25223), .Y(n30794) );
  NAND3X1 U18295 ( .A(n30803), .B(n30804), .C(n30805), .Y(n30792) );
  NOR2X1 U18296 ( .A(n30806), .B(n30807), .Y(n30805) );
  OAI22X1 U18297 ( .A(n25233), .B(n30808), .C(n25243), .D(n30809), .Y(n30807)
         );
  OAI22X1 U18298 ( .A(n25254), .B(n30810), .C(n25264), .D(n30811), .Y(n30806)
         );
  AOI22X1 U18299 ( .A(reg_file[626]), .B(n25275), .C(reg_file[754]), .D(n25286), .Y(n30804) );
  AOI22X1 U18300 ( .A(reg_file[882]), .B(n25296), .C(reg_file[1010]), .D(
        n25307), .Y(n30803) );
  NOR2X1 U18301 ( .A(n30812), .B(n30813), .Y(n30790) );
  NAND3X1 U18302 ( .A(n30814), .B(n30815), .C(n30816), .Y(n30813) );
  NOR2X1 U18303 ( .A(n30817), .B(n30818), .Y(n30816) );
  OAI22X1 U18304 ( .A(n25317), .B(n30819), .C(n25327), .D(n30820), .Y(n30818)
         );
  OAI22X1 U18305 ( .A(n25338), .B(n30821), .C(n25348), .D(n30822), .Y(n30817)
         );
  AOI22X1 U18306 ( .A(reg_file[3570]), .B(n25359), .C(reg_file[3442]), .D(
        n25370), .Y(n30815) );
  AOI22X1 U18307 ( .A(reg_file[3314]), .B(n25380), .C(reg_file[3186]), .D(
        n25391), .Y(n30814) );
  NAND3X1 U18308 ( .A(n30823), .B(n30824), .C(n30825), .Y(n30812) );
  NOR2X1 U18309 ( .A(n30826), .B(n30827), .Y(n30825) );
  OAI22X1 U18310 ( .A(n25401), .B(n30828), .C(n25411), .D(n30829), .Y(n30827)
         );
  OAI22X1 U18311 ( .A(n25422), .B(n30830), .C(n25432), .D(n30831), .Y(n30826)
         );
  AOI22X1 U18312 ( .A(reg_file[2546]), .B(n25443), .C(reg_file[2418]), .D(
        n25454), .Y(n30824) );
  AOI22X1 U18313 ( .A(reg_file[2290]), .B(n25464), .C(reg_file[2162]), .D(
        n25475), .Y(n30823) );
  AOI21X1 U18314 ( .A(n30832), .B(n30833), .C(n25138), .Y(rd2data1040_113_) );
  NOR2X1 U18315 ( .A(n30834), .B(n30835), .Y(n30833) );
  NAND3X1 U18316 ( .A(n30836), .B(n30837), .C(n30838), .Y(n30835) );
  NOR2X1 U18317 ( .A(n30839), .B(n30840), .Y(n30838) );
  OAI22X1 U18318 ( .A(n25149), .B(n30841), .C(n25159), .D(n30842), .Y(n30840)
         );
  OAI22X1 U18319 ( .A(n25170), .B(n30843), .C(n25180), .D(n30844), .Y(n30839)
         );
  AOI22X1 U18320 ( .A(reg_file[1521]), .B(n25191), .C(reg_file[1393]), .D(
        n25202), .Y(n30837) );
  AOI22X1 U18321 ( .A(reg_file[1265]), .B(n25212), .C(reg_file[1137]), .D(
        n25223), .Y(n30836) );
  NAND3X1 U18322 ( .A(n30845), .B(n30846), .C(n30847), .Y(n30834) );
  NOR2X1 U18323 ( .A(n30848), .B(n30849), .Y(n30847) );
  OAI22X1 U18324 ( .A(n25233), .B(n30850), .C(n25243), .D(n30851), .Y(n30849)
         );
  OAI22X1 U18325 ( .A(n25254), .B(n30852), .C(n25264), .D(n30853), .Y(n30848)
         );
  AOI22X1 U18326 ( .A(reg_file[625]), .B(n25275), .C(reg_file[753]), .D(n25286), .Y(n30846) );
  AOI22X1 U18327 ( .A(reg_file[881]), .B(n25296), .C(reg_file[1009]), .D(
        n25307), .Y(n30845) );
  NOR2X1 U18328 ( .A(n30854), .B(n30855), .Y(n30832) );
  NAND3X1 U18329 ( .A(n30856), .B(n30857), .C(n30858), .Y(n30855) );
  NOR2X1 U18330 ( .A(n30859), .B(n30860), .Y(n30858) );
  OAI22X1 U18331 ( .A(n25317), .B(n30861), .C(n25327), .D(n30862), .Y(n30860)
         );
  OAI22X1 U18332 ( .A(n25338), .B(n30863), .C(n25348), .D(n30864), .Y(n30859)
         );
  AOI22X1 U18333 ( .A(reg_file[3569]), .B(n25359), .C(reg_file[3441]), .D(
        n25370), .Y(n30857) );
  AOI22X1 U18334 ( .A(reg_file[3313]), .B(n25380), .C(reg_file[3185]), .D(
        n25391), .Y(n30856) );
  NAND3X1 U18335 ( .A(n30865), .B(n30866), .C(n30867), .Y(n30854) );
  NOR2X1 U18336 ( .A(n30868), .B(n30869), .Y(n30867) );
  OAI22X1 U18337 ( .A(n25401), .B(n30870), .C(n25411), .D(n30871), .Y(n30869)
         );
  OAI22X1 U18338 ( .A(n25422), .B(n30872), .C(n25432), .D(n30873), .Y(n30868)
         );
  AOI22X1 U18339 ( .A(reg_file[2545]), .B(n25443), .C(reg_file[2417]), .D(
        n25454), .Y(n30866) );
  AOI22X1 U18340 ( .A(reg_file[2289]), .B(n25464), .C(reg_file[2161]), .D(
        n25475), .Y(n30865) );
  AOI21X1 U18341 ( .A(n30874), .B(n30875), .C(n25138), .Y(rd2data1040_112_) );
  NOR2X1 U18342 ( .A(n30876), .B(n30877), .Y(n30875) );
  NAND3X1 U18343 ( .A(n30878), .B(n30879), .C(n30880), .Y(n30877) );
  NOR2X1 U18344 ( .A(n30881), .B(n30882), .Y(n30880) );
  OAI22X1 U18345 ( .A(n25149), .B(n30883), .C(n25159), .D(n30884), .Y(n30882)
         );
  OAI22X1 U18346 ( .A(n25170), .B(n30885), .C(n25180), .D(n30886), .Y(n30881)
         );
  AOI22X1 U18347 ( .A(reg_file[1520]), .B(n25191), .C(reg_file[1392]), .D(
        n25202), .Y(n30879) );
  AOI22X1 U18348 ( .A(reg_file[1264]), .B(n25212), .C(reg_file[1136]), .D(
        n25223), .Y(n30878) );
  NAND3X1 U18349 ( .A(n30887), .B(n30888), .C(n30889), .Y(n30876) );
  NOR2X1 U18350 ( .A(n30890), .B(n30891), .Y(n30889) );
  OAI22X1 U18351 ( .A(n25233), .B(n30892), .C(n25243), .D(n30893), .Y(n30891)
         );
  OAI22X1 U18352 ( .A(n25254), .B(n30894), .C(n25264), .D(n30895), .Y(n30890)
         );
  AOI22X1 U18353 ( .A(reg_file[624]), .B(n25275), .C(reg_file[752]), .D(n25286), .Y(n30888) );
  AOI22X1 U18354 ( .A(reg_file[880]), .B(n25296), .C(reg_file[1008]), .D(
        n25307), .Y(n30887) );
  NOR2X1 U18355 ( .A(n30896), .B(n30897), .Y(n30874) );
  NAND3X1 U18356 ( .A(n30898), .B(n30899), .C(n30900), .Y(n30897) );
  NOR2X1 U18357 ( .A(n30901), .B(n30902), .Y(n30900) );
  OAI22X1 U18358 ( .A(n25317), .B(n30903), .C(n25327), .D(n30904), .Y(n30902)
         );
  OAI22X1 U18359 ( .A(n25338), .B(n30905), .C(n25348), .D(n30906), .Y(n30901)
         );
  AOI22X1 U18360 ( .A(reg_file[3568]), .B(n25359), .C(reg_file[3440]), .D(
        n25370), .Y(n30899) );
  AOI22X1 U18361 ( .A(reg_file[3312]), .B(n25380), .C(reg_file[3184]), .D(
        n25391), .Y(n30898) );
  NAND3X1 U18362 ( .A(n30907), .B(n30908), .C(n30909), .Y(n30896) );
  NOR2X1 U18363 ( .A(n30910), .B(n30911), .Y(n30909) );
  OAI22X1 U18364 ( .A(n25401), .B(n30912), .C(n25411), .D(n30913), .Y(n30911)
         );
  OAI22X1 U18365 ( .A(n25422), .B(n30914), .C(n25432), .D(n30915), .Y(n30910)
         );
  AOI22X1 U18366 ( .A(reg_file[2544]), .B(n25443), .C(reg_file[2416]), .D(
        n25454), .Y(n30908) );
  AOI22X1 U18367 ( .A(reg_file[2288]), .B(n25464), .C(reg_file[2160]), .D(
        n25475), .Y(n30907) );
  AOI21X1 U18368 ( .A(n30916), .B(n30917), .C(n25138), .Y(rd2data1040_111_) );
  NOR2X1 U18369 ( .A(n30918), .B(n30919), .Y(n30917) );
  NAND3X1 U18370 ( .A(n30920), .B(n30921), .C(n30922), .Y(n30919) );
  NOR2X1 U18371 ( .A(n30923), .B(n30924), .Y(n30922) );
  OAI22X1 U18372 ( .A(n25149), .B(n30925), .C(n25159), .D(n30926), .Y(n30924)
         );
  OAI22X1 U18373 ( .A(n25170), .B(n30927), .C(n25180), .D(n30928), .Y(n30923)
         );
  AOI22X1 U18374 ( .A(reg_file[1519]), .B(n25191), .C(reg_file[1391]), .D(
        n25202), .Y(n30921) );
  AOI22X1 U18375 ( .A(reg_file[1263]), .B(n25212), .C(reg_file[1135]), .D(
        n25223), .Y(n30920) );
  NAND3X1 U18376 ( .A(n30929), .B(n30930), .C(n30931), .Y(n30918) );
  NOR2X1 U18377 ( .A(n30932), .B(n30933), .Y(n30931) );
  OAI22X1 U18378 ( .A(n25233), .B(n30934), .C(n25243), .D(n30935), .Y(n30933)
         );
  OAI22X1 U18379 ( .A(n25254), .B(n30936), .C(n25264), .D(n30937), .Y(n30932)
         );
  AOI22X1 U18380 ( .A(reg_file[623]), .B(n25275), .C(reg_file[751]), .D(n25286), .Y(n30930) );
  AOI22X1 U18381 ( .A(reg_file[879]), .B(n25296), .C(reg_file[1007]), .D(
        n25307), .Y(n30929) );
  NOR2X1 U18382 ( .A(n30938), .B(n30939), .Y(n30916) );
  NAND3X1 U18383 ( .A(n30940), .B(n30941), .C(n30942), .Y(n30939) );
  NOR2X1 U18384 ( .A(n30943), .B(n30944), .Y(n30942) );
  OAI22X1 U18385 ( .A(n25317), .B(n30945), .C(n25327), .D(n30946), .Y(n30944)
         );
  OAI22X1 U18386 ( .A(n25338), .B(n30947), .C(n25348), .D(n30948), .Y(n30943)
         );
  AOI22X1 U18387 ( .A(reg_file[3567]), .B(n25359), .C(reg_file[3439]), .D(
        n25370), .Y(n30941) );
  AOI22X1 U18388 ( .A(reg_file[3311]), .B(n25380), .C(reg_file[3183]), .D(
        n25391), .Y(n30940) );
  NAND3X1 U18389 ( .A(n30949), .B(n30950), .C(n30951), .Y(n30938) );
  NOR2X1 U18390 ( .A(n30952), .B(n30953), .Y(n30951) );
  OAI22X1 U18391 ( .A(n25401), .B(n30954), .C(n25411), .D(n30955), .Y(n30953)
         );
  OAI22X1 U18392 ( .A(n25422), .B(n30956), .C(n25432), .D(n30957), .Y(n30952)
         );
  AOI22X1 U18393 ( .A(reg_file[2543]), .B(n25443), .C(reg_file[2415]), .D(
        n25454), .Y(n30950) );
  AOI22X1 U18394 ( .A(reg_file[2287]), .B(n25464), .C(reg_file[2159]), .D(
        n25475), .Y(n30949) );
  AOI21X1 U18395 ( .A(n30958), .B(n30959), .C(n25138), .Y(rd2data1040_110_) );
  NOR2X1 U18396 ( .A(n30960), .B(n30961), .Y(n30959) );
  NAND3X1 U18397 ( .A(n30962), .B(n30963), .C(n30964), .Y(n30961) );
  NOR2X1 U18398 ( .A(n30965), .B(n30966), .Y(n30964) );
  OAI22X1 U18399 ( .A(n25148), .B(n30967), .C(n25159), .D(n30968), .Y(n30966)
         );
  OAI22X1 U18400 ( .A(n25169), .B(n30969), .C(n25180), .D(n30970), .Y(n30965)
         );
  AOI22X1 U18401 ( .A(reg_file[1518]), .B(n25191), .C(reg_file[1390]), .D(
        n25201), .Y(n30963) );
  AOI22X1 U18402 ( .A(reg_file[1262]), .B(n25212), .C(reg_file[1134]), .D(
        n25222), .Y(n30962) );
  NAND3X1 U18403 ( .A(n30971), .B(n30972), .C(n30973), .Y(n30960) );
  NOR2X1 U18404 ( .A(n30974), .B(n30975), .Y(n30973) );
  OAI22X1 U18405 ( .A(n25232), .B(n30976), .C(n25243), .D(n30977), .Y(n30975)
         );
  OAI22X1 U18406 ( .A(n25253), .B(n30978), .C(n25264), .D(n30979), .Y(n30974)
         );
  AOI22X1 U18407 ( .A(reg_file[622]), .B(n25275), .C(reg_file[750]), .D(n25285), .Y(n30972) );
  AOI22X1 U18408 ( .A(reg_file[878]), .B(n25296), .C(reg_file[1006]), .D(
        n25306), .Y(n30971) );
  NOR2X1 U18409 ( .A(n30980), .B(n30981), .Y(n30958) );
  NAND3X1 U18410 ( .A(n30982), .B(n30983), .C(n30984), .Y(n30981) );
  NOR2X1 U18411 ( .A(n30985), .B(n30986), .Y(n30984) );
  OAI22X1 U18412 ( .A(n25316), .B(n30987), .C(n25327), .D(n30988), .Y(n30986)
         );
  OAI22X1 U18413 ( .A(n25337), .B(n30989), .C(n25348), .D(n30990), .Y(n30985)
         );
  AOI22X1 U18414 ( .A(reg_file[3566]), .B(n25359), .C(reg_file[3438]), .D(
        n25369), .Y(n30983) );
  AOI22X1 U18415 ( .A(reg_file[3310]), .B(n25380), .C(reg_file[3182]), .D(
        n25390), .Y(n30982) );
  NAND3X1 U18416 ( .A(n30991), .B(n30992), .C(n30993), .Y(n30980) );
  NOR2X1 U18417 ( .A(n30994), .B(n30995), .Y(n30993) );
  OAI22X1 U18418 ( .A(n25400), .B(n30996), .C(n25411), .D(n30997), .Y(n30995)
         );
  OAI22X1 U18419 ( .A(n25421), .B(n30998), .C(n25432), .D(n30999), .Y(n30994)
         );
  AOI22X1 U18420 ( .A(reg_file[2542]), .B(n25443), .C(reg_file[2414]), .D(
        n25453), .Y(n30992) );
  AOI22X1 U18421 ( .A(reg_file[2286]), .B(n25464), .C(reg_file[2158]), .D(
        n25474), .Y(n30991) );
  AOI21X1 U18422 ( .A(n31000), .B(n31001), .C(n25137), .Y(rd2data1040_10_) );
  NOR2X1 U18423 ( .A(n31002), .B(n31003), .Y(n31001) );
  NAND3X1 U18424 ( .A(n31004), .B(n31005), .C(n31006), .Y(n31003) );
  NOR2X1 U18425 ( .A(n31007), .B(n31008), .Y(n31006) );
  OAI22X1 U18426 ( .A(n25148), .B(n31009), .C(n25158), .D(n31010), .Y(n31008)
         );
  OAI22X1 U18427 ( .A(n25169), .B(n31011), .C(n25179), .D(n31012), .Y(n31007)
         );
  AOI22X1 U18428 ( .A(reg_file[1418]), .B(n25190), .C(reg_file[1290]), .D(
        n25201), .Y(n31005) );
  AOI22X1 U18429 ( .A(reg_file[1162]), .B(n25211), .C(reg_file[1034]), .D(
        n25222), .Y(n31004) );
  NAND3X1 U18430 ( .A(n31013), .B(n31014), .C(n31015), .Y(n31002) );
  NOR2X1 U18431 ( .A(n31016), .B(n31017), .Y(n31015) );
  OAI22X1 U18432 ( .A(n25232), .B(n31018), .C(n25242), .D(n31019), .Y(n31017)
         );
  OAI22X1 U18433 ( .A(n25253), .B(n31020), .C(n25263), .D(n31021), .Y(n31016)
         );
  AOI22X1 U18434 ( .A(reg_file[522]), .B(n25274), .C(reg_file[650]), .D(n25285), .Y(n31014) );
  AOI22X1 U18435 ( .A(reg_file[778]), .B(n25295), .C(reg_file[906]), .D(n25306), .Y(n31013) );
  NOR2X1 U18436 ( .A(n31022), .B(n31023), .Y(n31000) );
  NAND3X1 U18437 ( .A(n31024), .B(n31025), .C(n31026), .Y(n31023) );
  NOR2X1 U18438 ( .A(n31027), .B(n31028), .Y(n31026) );
  OAI22X1 U18439 ( .A(n25316), .B(n31029), .C(n25326), .D(n31030), .Y(n31028)
         );
  OAI22X1 U18440 ( .A(n25337), .B(n31031), .C(n25347), .D(n31032), .Y(n31027)
         );
  AOI22X1 U18441 ( .A(reg_file[3466]), .B(n25358), .C(reg_file[3338]), .D(
        n25369), .Y(n31025) );
  AOI22X1 U18442 ( .A(reg_file[3210]), .B(n25379), .C(reg_file[3082]), .D(
        n25390), .Y(n31024) );
  NAND3X1 U18443 ( .A(n31033), .B(n31034), .C(n31035), .Y(n31022) );
  NOR2X1 U18444 ( .A(n31036), .B(n31037), .Y(n31035) );
  OAI22X1 U18445 ( .A(n25400), .B(n31038), .C(n25410), .D(n31039), .Y(n31037)
         );
  OAI22X1 U18446 ( .A(n25421), .B(n31040), .C(n25431), .D(n31041), .Y(n31036)
         );
  AOI22X1 U18447 ( .A(reg_file[2442]), .B(n25442), .C(reg_file[2314]), .D(
        n25453), .Y(n31034) );
  AOI22X1 U18448 ( .A(reg_file[2186]), .B(n25463), .C(reg_file[2058]), .D(
        n25474), .Y(n31033) );
  AOI21X1 U18449 ( .A(n31042), .B(n31043), .C(n25137), .Y(rd2data1040_109_) );
  NOR2X1 U18450 ( .A(n31044), .B(n31045), .Y(n31043) );
  NAND3X1 U18451 ( .A(n31046), .B(n31047), .C(n31048), .Y(n31045) );
  NOR2X1 U18452 ( .A(n31049), .B(n31050), .Y(n31048) );
  OAI22X1 U18453 ( .A(n25148), .B(n31051), .C(n25158), .D(n31052), .Y(n31050)
         );
  OAI22X1 U18454 ( .A(n25169), .B(n31053), .C(n25179), .D(n31054), .Y(n31049)
         );
  AOI22X1 U18455 ( .A(reg_file[1517]), .B(n25190), .C(reg_file[1389]), .D(
        n25201), .Y(n31047) );
  AOI22X1 U18456 ( .A(reg_file[1261]), .B(n25211), .C(reg_file[1133]), .D(
        n25222), .Y(n31046) );
  NAND3X1 U18457 ( .A(n31055), .B(n31056), .C(n31057), .Y(n31044) );
  NOR2X1 U18458 ( .A(n31058), .B(n31059), .Y(n31057) );
  OAI22X1 U18459 ( .A(n25232), .B(n31060), .C(n25242), .D(n31061), .Y(n31059)
         );
  OAI22X1 U18460 ( .A(n25253), .B(n31062), .C(n25263), .D(n31063), .Y(n31058)
         );
  AOI22X1 U18461 ( .A(reg_file[621]), .B(n25274), .C(reg_file[749]), .D(n25285), .Y(n31056) );
  AOI22X1 U18462 ( .A(reg_file[877]), .B(n25295), .C(reg_file[1005]), .D(
        n25306), .Y(n31055) );
  NOR2X1 U18463 ( .A(n31064), .B(n31065), .Y(n31042) );
  NAND3X1 U18464 ( .A(n31066), .B(n31067), .C(n31068), .Y(n31065) );
  NOR2X1 U18465 ( .A(n31069), .B(n31070), .Y(n31068) );
  OAI22X1 U18466 ( .A(n25316), .B(n31071), .C(n25326), .D(n31072), .Y(n31070)
         );
  OAI22X1 U18467 ( .A(n25337), .B(n31073), .C(n25347), .D(n31074), .Y(n31069)
         );
  AOI22X1 U18468 ( .A(reg_file[3565]), .B(n25358), .C(reg_file[3437]), .D(
        n25369), .Y(n31067) );
  AOI22X1 U18469 ( .A(reg_file[3309]), .B(n25379), .C(reg_file[3181]), .D(
        n25390), .Y(n31066) );
  NAND3X1 U18470 ( .A(n31075), .B(n31076), .C(n31077), .Y(n31064) );
  NOR2X1 U18471 ( .A(n31078), .B(n31079), .Y(n31077) );
  OAI22X1 U18472 ( .A(n25400), .B(n31080), .C(n25410), .D(n31081), .Y(n31079)
         );
  OAI22X1 U18473 ( .A(n25421), .B(n31082), .C(n25431), .D(n31083), .Y(n31078)
         );
  AOI22X1 U18474 ( .A(reg_file[2541]), .B(n25442), .C(reg_file[2413]), .D(
        n25453), .Y(n31076) );
  AOI22X1 U18475 ( .A(reg_file[2285]), .B(n25463), .C(reg_file[2157]), .D(
        n25474), .Y(n31075) );
  AOI21X1 U18476 ( .A(n31084), .B(n31085), .C(n25137), .Y(rd2data1040_108_) );
  NOR2X1 U18477 ( .A(n31086), .B(n31087), .Y(n31085) );
  NAND3X1 U18478 ( .A(n31088), .B(n31089), .C(n31090), .Y(n31087) );
  NOR2X1 U18479 ( .A(n31091), .B(n31092), .Y(n31090) );
  OAI22X1 U18480 ( .A(n25148), .B(n31093), .C(n25158), .D(n31094), .Y(n31092)
         );
  OAI22X1 U18481 ( .A(n25169), .B(n31095), .C(n25179), .D(n31096), .Y(n31091)
         );
  AOI22X1 U18482 ( .A(reg_file[1516]), .B(n25190), .C(reg_file[1388]), .D(
        n25201), .Y(n31089) );
  AOI22X1 U18483 ( .A(reg_file[1260]), .B(n25211), .C(reg_file[1132]), .D(
        n25222), .Y(n31088) );
  NAND3X1 U18484 ( .A(n31097), .B(n31098), .C(n31099), .Y(n31086) );
  NOR2X1 U18485 ( .A(n31100), .B(n31101), .Y(n31099) );
  OAI22X1 U18486 ( .A(n25232), .B(n31102), .C(n25242), .D(n31103), .Y(n31101)
         );
  OAI22X1 U18487 ( .A(n25253), .B(n31104), .C(n25263), .D(n31105), .Y(n31100)
         );
  AOI22X1 U18488 ( .A(reg_file[620]), .B(n25274), .C(reg_file[748]), .D(n25285), .Y(n31098) );
  AOI22X1 U18489 ( .A(reg_file[876]), .B(n25295), .C(reg_file[1004]), .D(
        n25306), .Y(n31097) );
  NOR2X1 U18490 ( .A(n31106), .B(n31107), .Y(n31084) );
  NAND3X1 U18491 ( .A(n31108), .B(n31109), .C(n31110), .Y(n31107) );
  NOR2X1 U18492 ( .A(n31111), .B(n31112), .Y(n31110) );
  OAI22X1 U18493 ( .A(n25316), .B(n31113), .C(n25326), .D(n31114), .Y(n31112)
         );
  OAI22X1 U18494 ( .A(n25337), .B(n31115), .C(n25347), .D(n31116), .Y(n31111)
         );
  AOI22X1 U18495 ( .A(reg_file[3564]), .B(n25358), .C(reg_file[3436]), .D(
        n25369), .Y(n31109) );
  AOI22X1 U18496 ( .A(reg_file[3308]), .B(n25379), .C(reg_file[3180]), .D(
        n25390), .Y(n31108) );
  NAND3X1 U18497 ( .A(n31117), .B(n31118), .C(n31119), .Y(n31106) );
  NOR2X1 U18498 ( .A(n31120), .B(n31121), .Y(n31119) );
  OAI22X1 U18499 ( .A(n25400), .B(n31122), .C(n25410), .D(n31123), .Y(n31121)
         );
  OAI22X1 U18500 ( .A(n25421), .B(n31124), .C(n25431), .D(n31125), .Y(n31120)
         );
  AOI22X1 U18501 ( .A(reg_file[2540]), .B(n25442), .C(reg_file[2412]), .D(
        n25453), .Y(n31118) );
  AOI22X1 U18502 ( .A(reg_file[2284]), .B(n25463), .C(reg_file[2156]), .D(
        n25474), .Y(n31117) );
  AOI21X1 U18503 ( .A(n31126), .B(n31127), .C(n25137), .Y(rd2data1040_107_) );
  NOR2X1 U18504 ( .A(n31128), .B(n31129), .Y(n31127) );
  NAND3X1 U18505 ( .A(n31130), .B(n31131), .C(n31132), .Y(n31129) );
  NOR2X1 U18506 ( .A(n31133), .B(n31134), .Y(n31132) );
  OAI22X1 U18507 ( .A(n25148), .B(n31135), .C(n25158), .D(n31136), .Y(n31134)
         );
  OAI22X1 U18508 ( .A(n25169), .B(n31137), .C(n25179), .D(n31138), .Y(n31133)
         );
  AOI22X1 U18509 ( .A(reg_file[1515]), .B(n25190), .C(reg_file[1387]), .D(
        n25201), .Y(n31131) );
  AOI22X1 U18510 ( .A(reg_file[1259]), .B(n25211), .C(reg_file[1131]), .D(
        n25222), .Y(n31130) );
  NAND3X1 U18511 ( .A(n31139), .B(n31140), .C(n31141), .Y(n31128) );
  NOR2X1 U18512 ( .A(n31142), .B(n31143), .Y(n31141) );
  OAI22X1 U18513 ( .A(n25232), .B(n31144), .C(n25242), .D(n31145), .Y(n31143)
         );
  OAI22X1 U18514 ( .A(n25253), .B(n31146), .C(n25263), .D(n31147), .Y(n31142)
         );
  AOI22X1 U18515 ( .A(reg_file[619]), .B(n25274), .C(reg_file[747]), .D(n25285), .Y(n31140) );
  AOI22X1 U18516 ( .A(reg_file[875]), .B(n25295), .C(reg_file[1003]), .D(
        n25306), .Y(n31139) );
  NOR2X1 U18517 ( .A(n31148), .B(n31149), .Y(n31126) );
  NAND3X1 U18518 ( .A(n31150), .B(n31151), .C(n31152), .Y(n31149) );
  NOR2X1 U18519 ( .A(n31153), .B(n31154), .Y(n31152) );
  OAI22X1 U18520 ( .A(n25316), .B(n31155), .C(n25326), .D(n31156), .Y(n31154)
         );
  OAI22X1 U18521 ( .A(n25337), .B(n31157), .C(n25347), .D(n31158), .Y(n31153)
         );
  AOI22X1 U18522 ( .A(reg_file[3563]), .B(n25358), .C(reg_file[3435]), .D(
        n25369), .Y(n31151) );
  AOI22X1 U18523 ( .A(reg_file[3307]), .B(n25379), .C(reg_file[3179]), .D(
        n25390), .Y(n31150) );
  NAND3X1 U18524 ( .A(n31159), .B(n31160), .C(n31161), .Y(n31148) );
  NOR2X1 U18525 ( .A(n31162), .B(n31163), .Y(n31161) );
  OAI22X1 U18526 ( .A(n25400), .B(n31164), .C(n25410), .D(n31165), .Y(n31163)
         );
  OAI22X1 U18527 ( .A(n25421), .B(n31166), .C(n25431), .D(n31167), .Y(n31162)
         );
  AOI22X1 U18528 ( .A(reg_file[2539]), .B(n25442), .C(reg_file[2411]), .D(
        n25453), .Y(n31160) );
  AOI22X1 U18529 ( .A(reg_file[2283]), .B(n25463), .C(reg_file[2155]), .D(
        n25474), .Y(n31159) );
  AOI21X1 U18530 ( .A(n31168), .B(n31169), .C(n25137), .Y(rd2data1040_106_) );
  NOR2X1 U18531 ( .A(n31170), .B(n31171), .Y(n31169) );
  NAND3X1 U18532 ( .A(n31172), .B(n31173), .C(n31174), .Y(n31171) );
  NOR2X1 U18533 ( .A(n31175), .B(n31176), .Y(n31174) );
  OAI22X1 U18534 ( .A(n25148), .B(n31177), .C(n25158), .D(n31178), .Y(n31176)
         );
  OAI22X1 U18535 ( .A(n25169), .B(n31179), .C(n25179), .D(n31180), .Y(n31175)
         );
  AOI22X1 U18536 ( .A(reg_file[1514]), .B(n25190), .C(reg_file[1386]), .D(
        n25201), .Y(n31173) );
  AOI22X1 U18537 ( .A(reg_file[1258]), .B(n25211), .C(reg_file[1130]), .D(
        n25222), .Y(n31172) );
  NAND3X1 U18538 ( .A(n31181), .B(n31182), .C(n31183), .Y(n31170) );
  NOR2X1 U18539 ( .A(n31184), .B(n31185), .Y(n31183) );
  OAI22X1 U18540 ( .A(n25232), .B(n31186), .C(n25242), .D(n31187), .Y(n31185)
         );
  OAI22X1 U18541 ( .A(n25253), .B(n31188), .C(n25263), .D(n31189), .Y(n31184)
         );
  AOI22X1 U18542 ( .A(reg_file[618]), .B(n25274), .C(reg_file[746]), .D(n25285), .Y(n31182) );
  AOI22X1 U18543 ( .A(reg_file[874]), .B(n25295), .C(reg_file[1002]), .D(
        n25306), .Y(n31181) );
  NOR2X1 U18544 ( .A(n31190), .B(n31191), .Y(n31168) );
  NAND3X1 U18545 ( .A(n31192), .B(n31193), .C(n31194), .Y(n31191) );
  NOR2X1 U18546 ( .A(n31195), .B(n31196), .Y(n31194) );
  OAI22X1 U18547 ( .A(n25316), .B(n31197), .C(n25326), .D(n31198), .Y(n31196)
         );
  OAI22X1 U18548 ( .A(n25337), .B(n31199), .C(n25347), .D(n31200), .Y(n31195)
         );
  AOI22X1 U18549 ( .A(reg_file[3562]), .B(n25358), .C(reg_file[3434]), .D(
        n25369), .Y(n31193) );
  AOI22X1 U18550 ( .A(reg_file[3306]), .B(n25379), .C(reg_file[3178]), .D(
        n25390), .Y(n31192) );
  NAND3X1 U18551 ( .A(n31201), .B(n31202), .C(n31203), .Y(n31190) );
  NOR2X1 U18552 ( .A(n31204), .B(n31205), .Y(n31203) );
  OAI22X1 U18553 ( .A(n25400), .B(n31206), .C(n25410), .D(n31207), .Y(n31205)
         );
  OAI22X1 U18554 ( .A(n25421), .B(n31208), .C(n25431), .D(n31209), .Y(n31204)
         );
  AOI22X1 U18555 ( .A(reg_file[2538]), .B(n25442), .C(reg_file[2410]), .D(
        n25453), .Y(n31202) );
  AOI22X1 U18556 ( .A(reg_file[2282]), .B(n25463), .C(reg_file[2154]), .D(
        n25474), .Y(n31201) );
  AOI21X1 U18557 ( .A(n31210), .B(n31211), .C(n25137), .Y(rd2data1040_105_) );
  NOR2X1 U18558 ( .A(n31212), .B(n31213), .Y(n31211) );
  NAND3X1 U18559 ( .A(n31214), .B(n31215), .C(n31216), .Y(n31213) );
  NOR2X1 U18560 ( .A(n31217), .B(n31218), .Y(n31216) );
  OAI22X1 U18561 ( .A(n25148), .B(n31219), .C(n25158), .D(n31220), .Y(n31218)
         );
  OAI22X1 U18562 ( .A(n25169), .B(n31221), .C(n25179), .D(n31222), .Y(n31217)
         );
  AOI22X1 U18563 ( .A(reg_file[1513]), .B(n25190), .C(reg_file[1385]), .D(
        n25201), .Y(n31215) );
  AOI22X1 U18564 ( .A(reg_file[1257]), .B(n25211), .C(reg_file[1129]), .D(
        n25222), .Y(n31214) );
  NAND3X1 U18565 ( .A(n31223), .B(n31224), .C(n31225), .Y(n31212) );
  NOR2X1 U18566 ( .A(n31226), .B(n31227), .Y(n31225) );
  OAI22X1 U18567 ( .A(n25232), .B(n31228), .C(n25242), .D(n31229), .Y(n31227)
         );
  OAI22X1 U18568 ( .A(n25253), .B(n31230), .C(n25263), .D(n31231), .Y(n31226)
         );
  AOI22X1 U18569 ( .A(reg_file[617]), .B(n25274), .C(reg_file[745]), .D(n25285), .Y(n31224) );
  AOI22X1 U18570 ( .A(reg_file[873]), .B(n25295), .C(reg_file[1001]), .D(
        n25306), .Y(n31223) );
  NOR2X1 U18571 ( .A(n31232), .B(n31233), .Y(n31210) );
  NAND3X1 U18572 ( .A(n31234), .B(n31235), .C(n31236), .Y(n31233) );
  NOR2X1 U18573 ( .A(n31237), .B(n31238), .Y(n31236) );
  OAI22X1 U18574 ( .A(n25316), .B(n31239), .C(n25326), .D(n31240), .Y(n31238)
         );
  OAI22X1 U18575 ( .A(n25337), .B(n31241), .C(n25347), .D(n31242), .Y(n31237)
         );
  AOI22X1 U18576 ( .A(reg_file[3561]), .B(n25358), .C(reg_file[3433]), .D(
        n25369), .Y(n31235) );
  AOI22X1 U18577 ( .A(reg_file[3305]), .B(n25379), .C(reg_file[3177]), .D(
        n25390), .Y(n31234) );
  NAND3X1 U18578 ( .A(n31243), .B(n31244), .C(n31245), .Y(n31232) );
  NOR2X1 U18579 ( .A(n31246), .B(n31247), .Y(n31245) );
  OAI22X1 U18580 ( .A(n25400), .B(n31248), .C(n25410), .D(n31249), .Y(n31247)
         );
  OAI22X1 U18581 ( .A(n25421), .B(n31250), .C(n25431), .D(n31251), .Y(n31246)
         );
  AOI22X1 U18582 ( .A(reg_file[2537]), .B(n25442), .C(reg_file[2409]), .D(
        n25453), .Y(n31244) );
  AOI22X1 U18583 ( .A(reg_file[2281]), .B(n25463), .C(reg_file[2153]), .D(
        n25474), .Y(n31243) );
  AOI21X1 U18584 ( .A(n31252), .B(n31253), .C(n25137), .Y(rd2data1040_104_) );
  NOR2X1 U18585 ( .A(n31254), .B(n31255), .Y(n31253) );
  NAND3X1 U18586 ( .A(n31256), .B(n31257), .C(n31258), .Y(n31255) );
  NOR2X1 U18587 ( .A(n31259), .B(n31260), .Y(n31258) );
  OAI22X1 U18588 ( .A(n25148), .B(n31261), .C(n25158), .D(n31262), .Y(n31260)
         );
  OAI22X1 U18589 ( .A(n25169), .B(n31263), .C(n25179), .D(n31264), .Y(n31259)
         );
  AOI22X1 U18590 ( .A(reg_file[1512]), .B(n25190), .C(reg_file[1384]), .D(
        n25201), .Y(n31257) );
  AOI22X1 U18591 ( .A(reg_file[1256]), .B(n25211), .C(reg_file[1128]), .D(
        n25222), .Y(n31256) );
  NAND3X1 U18592 ( .A(n31265), .B(n31266), .C(n31267), .Y(n31254) );
  NOR2X1 U18593 ( .A(n31268), .B(n31269), .Y(n31267) );
  OAI22X1 U18594 ( .A(n25232), .B(n31270), .C(n25242), .D(n31271), .Y(n31269)
         );
  OAI22X1 U18595 ( .A(n25253), .B(n31272), .C(n25263), .D(n31273), .Y(n31268)
         );
  AOI22X1 U18596 ( .A(reg_file[616]), .B(n25274), .C(reg_file[744]), .D(n25285), .Y(n31266) );
  AOI22X1 U18597 ( .A(reg_file[872]), .B(n25295), .C(reg_file[1000]), .D(
        n25306), .Y(n31265) );
  NOR2X1 U18598 ( .A(n31274), .B(n31275), .Y(n31252) );
  NAND3X1 U18599 ( .A(n31276), .B(n31277), .C(n31278), .Y(n31275) );
  NOR2X1 U18600 ( .A(n31279), .B(n31280), .Y(n31278) );
  OAI22X1 U18601 ( .A(n25316), .B(n31281), .C(n25326), .D(n31282), .Y(n31280)
         );
  OAI22X1 U18602 ( .A(n25337), .B(n31283), .C(n25347), .D(n31284), .Y(n31279)
         );
  AOI22X1 U18603 ( .A(reg_file[3560]), .B(n25358), .C(reg_file[3432]), .D(
        n25369), .Y(n31277) );
  AOI22X1 U18604 ( .A(reg_file[3304]), .B(n25379), .C(reg_file[3176]), .D(
        n25390), .Y(n31276) );
  NAND3X1 U18605 ( .A(n31285), .B(n31286), .C(n31287), .Y(n31274) );
  NOR2X1 U18606 ( .A(n31288), .B(n31289), .Y(n31287) );
  OAI22X1 U18607 ( .A(n25400), .B(n31290), .C(n25410), .D(n31291), .Y(n31289)
         );
  OAI22X1 U18608 ( .A(n25421), .B(n31292), .C(n25431), .D(n31293), .Y(n31288)
         );
  AOI22X1 U18609 ( .A(reg_file[2536]), .B(n25442), .C(reg_file[2408]), .D(
        n25453), .Y(n31286) );
  AOI22X1 U18610 ( .A(reg_file[2280]), .B(n25463), .C(reg_file[2152]), .D(
        n25474), .Y(n31285) );
  AOI21X1 U18611 ( .A(n31294), .B(n31295), .C(n25137), .Y(rd2data1040_103_) );
  NOR2X1 U18612 ( .A(n31296), .B(n31297), .Y(n31295) );
  NAND3X1 U18613 ( .A(n31298), .B(n31299), .C(n31300), .Y(n31297) );
  NOR2X1 U18614 ( .A(n31301), .B(n31302), .Y(n31300) );
  OAI22X1 U18615 ( .A(n25148), .B(n31303), .C(n25158), .D(n31304), .Y(n31302)
         );
  OAI22X1 U18616 ( .A(n25169), .B(n31305), .C(n25179), .D(n31306), .Y(n31301)
         );
  AOI22X1 U18617 ( .A(reg_file[1511]), .B(n25190), .C(reg_file[1383]), .D(
        n25201), .Y(n31299) );
  AOI22X1 U18618 ( .A(reg_file[1255]), .B(n25211), .C(reg_file[1127]), .D(
        n25222), .Y(n31298) );
  NAND3X1 U18619 ( .A(n31307), .B(n31308), .C(n31309), .Y(n31296) );
  NOR2X1 U18620 ( .A(n31310), .B(n31311), .Y(n31309) );
  OAI22X1 U18621 ( .A(n25232), .B(n31312), .C(n25242), .D(n31313), .Y(n31311)
         );
  OAI22X1 U18622 ( .A(n25253), .B(n31314), .C(n25263), .D(n31315), .Y(n31310)
         );
  AOI22X1 U18623 ( .A(reg_file[615]), .B(n25274), .C(reg_file[743]), .D(n25285), .Y(n31308) );
  AOI22X1 U18624 ( .A(reg_file[871]), .B(n25295), .C(reg_file[999]), .D(n25306), .Y(n31307) );
  NOR2X1 U18625 ( .A(n31316), .B(n31317), .Y(n31294) );
  NAND3X1 U18626 ( .A(n31318), .B(n31319), .C(n31320), .Y(n31317) );
  NOR2X1 U18627 ( .A(n31321), .B(n31322), .Y(n31320) );
  OAI22X1 U18628 ( .A(n25316), .B(n31323), .C(n25326), .D(n31324), .Y(n31322)
         );
  OAI22X1 U18629 ( .A(n25337), .B(n31325), .C(n25347), .D(n31326), .Y(n31321)
         );
  AOI22X1 U18630 ( .A(reg_file[3559]), .B(n25358), .C(reg_file[3431]), .D(
        n25369), .Y(n31319) );
  AOI22X1 U18631 ( .A(reg_file[3303]), .B(n25379), .C(reg_file[3175]), .D(
        n25390), .Y(n31318) );
  NAND3X1 U18632 ( .A(n31327), .B(n31328), .C(n31329), .Y(n31316) );
  NOR2X1 U18633 ( .A(n31330), .B(n31331), .Y(n31329) );
  OAI22X1 U18634 ( .A(n25400), .B(n31332), .C(n25410), .D(n31333), .Y(n31331)
         );
  OAI22X1 U18635 ( .A(n25421), .B(n31334), .C(n25431), .D(n31335), .Y(n31330)
         );
  AOI22X1 U18636 ( .A(reg_file[2535]), .B(n25442), .C(reg_file[2407]), .D(
        n25453), .Y(n31328) );
  AOI22X1 U18637 ( .A(reg_file[2279]), .B(n25463), .C(reg_file[2151]), .D(
        n25474), .Y(n31327) );
  AOI21X1 U18638 ( .A(n31336), .B(n31337), .C(n25137), .Y(rd2data1040_102_) );
  NOR2X1 U18639 ( .A(n31338), .B(n31339), .Y(n31337) );
  NAND3X1 U18640 ( .A(n31340), .B(n31341), .C(n31342), .Y(n31339) );
  NOR2X1 U18641 ( .A(n31343), .B(n31344), .Y(n31342) );
  OAI22X1 U18642 ( .A(n25148), .B(n31345), .C(n25158), .D(n31346), .Y(n31344)
         );
  OAI22X1 U18643 ( .A(n25169), .B(n31347), .C(n25179), .D(n31348), .Y(n31343)
         );
  AOI22X1 U18644 ( .A(reg_file[1510]), .B(n25190), .C(reg_file[1382]), .D(
        n25201), .Y(n31341) );
  AOI22X1 U18645 ( .A(reg_file[1254]), .B(n25211), .C(reg_file[1126]), .D(
        n25222), .Y(n31340) );
  NAND3X1 U18646 ( .A(n31349), .B(n31350), .C(n31351), .Y(n31338) );
  NOR2X1 U18647 ( .A(n31352), .B(n31353), .Y(n31351) );
  OAI22X1 U18648 ( .A(n25232), .B(n31354), .C(n25242), .D(n31355), .Y(n31353)
         );
  OAI22X1 U18649 ( .A(n25253), .B(n31356), .C(n25263), .D(n31357), .Y(n31352)
         );
  AOI22X1 U18650 ( .A(reg_file[614]), .B(n25274), .C(reg_file[742]), .D(n25285), .Y(n31350) );
  AOI22X1 U18651 ( .A(reg_file[870]), .B(n25295), .C(reg_file[998]), .D(n25306), .Y(n31349) );
  NOR2X1 U18652 ( .A(n31358), .B(n31359), .Y(n31336) );
  NAND3X1 U18653 ( .A(n31360), .B(n31361), .C(n31362), .Y(n31359) );
  NOR2X1 U18654 ( .A(n31363), .B(n31364), .Y(n31362) );
  OAI22X1 U18655 ( .A(n25316), .B(n31365), .C(n25326), .D(n31366), .Y(n31364)
         );
  OAI22X1 U18656 ( .A(n25337), .B(n31367), .C(n25347), .D(n31368), .Y(n31363)
         );
  AOI22X1 U18657 ( .A(reg_file[3558]), .B(n25358), .C(reg_file[3430]), .D(
        n25369), .Y(n31361) );
  AOI22X1 U18658 ( .A(reg_file[3302]), .B(n25379), .C(reg_file[3174]), .D(
        n25390), .Y(n31360) );
  NAND3X1 U18659 ( .A(n31369), .B(n31370), .C(n31371), .Y(n31358) );
  NOR2X1 U18660 ( .A(n31372), .B(n31373), .Y(n31371) );
  OAI22X1 U18661 ( .A(n25400), .B(n31374), .C(n25410), .D(n31375), .Y(n31373)
         );
  OAI22X1 U18662 ( .A(n25421), .B(n31376), .C(n25431), .D(n31377), .Y(n31372)
         );
  AOI22X1 U18663 ( .A(reg_file[2534]), .B(n25442), .C(reg_file[2406]), .D(
        n25453), .Y(n31370) );
  AOI22X1 U18664 ( .A(reg_file[2278]), .B(n25463), .C(reg_file[2150]), .D(
        n25474), .Y(n31369) );
  AOI21X1 U18665 ( .A(n31378), .B(n31379), .C(n25137), .Y(rd2data1040_101_) );
  NOR2X1 U18666 ( .A(n31380), .B(n31381), .Y(n31379) );
  NAND3X1 U18667 ( .A(n31382), .B(n31383), .C(n31384), .Y(n31381) );
  NOR2X1 U18668 ( .A(n31385), .B(n31386), .Y(n31384) );
  OAI22X1 U18669 ( .A(n25148), .B(n31387), .C(n25158), .D(n31388), .Y(n31386)
         );
  OAI22X1 U18670 ( .A(n25169), .B(n31389), .C(n25179), .D(n31390), .Y(n31385)
         );
  AOI22X1 U18671 ( .A(reg_file[1509]), .B(n25190), .C(reg_file[1381]), .D(
        n25201), .Y(n31383) );
  AOI22X1 U18672 ( .A(reg_file[1253]), .B(n25211), .C(reg_file[1125]), .D(
        n25222), .Y(n31382) );
  NAND3X1 U18673 ( .A(n31391), .B(n31392), .C(n31393), .Y(n31380) );
  NOR2X1 U18674 ( .A(n31394), .B(n31395), .Y(n31393) );
  OAI22X1 U18675 ( .A(n25232), .B(n31396), .C(n25242), .D(n31397), .Y(n31395)
         );
  OAI22X1 U18676 ( .A(n25253), .B(n31398), .C(n25263), .D(n31399), .Y(n31394)
         );
  AOI22X1 U18677 ( .A(reg_file[613]), .B(n25274), .C(reg_file[741]), .D(n25285), .Y(n31392) );
  AOI22X1 U18678 ( .A(reg_file[869]), .B(n25295), .C(reg_file[997]), .D(n25306), .Y(n31391) );
  NOR2X1 U18679 ( .A(n31400), .B(n31401), .Y(n31378) );
  NAND3X1 U18680 ( .A(n31402), .B(n31403), .C(n31404), .Y(n31401) );
  NOR2X1 U18681 ( .A(n31405), .B(n31406), .Y(n31404) );
  OAI22X1 U18682 ( .A(n25316), .B(n31407), .C(n25326), .D(n31408), .Y(n31406)
         );
  OAI22X1 U18683 ( .A(n25337), .B(n31409), .C(n25347), .D(n31410), .Y(n31405)
         );
  AOI22X1 U18684 ( .A(reg_file[3557]), .B(n25358), .C(reg_file[3429]), .D(
        n25369), .Y(n31403) );
  AOI22X1 U18685 ( .A(reg_file[3301]), .B(n25379), .C(reg_file[3173]), .D(
        n25390), .Y(n31402) );
  NAND3X1 U18686 ( .A(n31411), .B(n31412), .C(n31413), .Y(n31400) );
  NOR2X1 U18687 ( .A(n31414), .B(n31415), .Y(n31413) );
  OAI22X1 U18688 ( .A(n25400), .B(n31416), .C(n25410), .D(n31417), .Y(n31415)
         );
  OAI22X1 U18689 ( .A(n25421), .B(n31418), .C(n25431), .D(n31419), .Y(n31414)
         );
  AOI22X1 U18690 ( .A(reg_file[2533]), .B(n25442), .C(reg_file[2405]), .D(
        n25453), .Y(n31412) );
  AOI22X1 U18691 ( .A(reg_file[2277]), .B(n25463), .C(reg_file[2149]), .D(
        n25474), .Y(n31411) );
  AOI21X1 U18692 ( .A(n31420), .B(n31421), .C(n25137), .Y(rd2data1040_100_) );
  NOR2X1 U18693 ( .A(n31422), .B(n31423), .Y(n31421) );
  NAND3X1 U18694 ( .A(n31424), .B(n31425), .C(n31426), .Y(n31423) );
  NOR2X1 U18695 ( .A(n31427), .B(n31428), .Y(n31426) );
  OAI22X1 U18696 ( .A(n25148), .B(n31429), .C(n25158), .D(n31430), .Y(n31428)
         );
  OAI22X1 U18697 ( .A(n25169), .B(n31431), .C(n25179), .D(n31432), .Y(n31427)
         );
  AOI22X1 U18698 ( .A(reg_file[1508]), .B(n25190), .C(reg_file[1380]), .D(
        n25201), .Y(n31425) );
  AOI22X1 U18699 ( .A(reg_file[1252]), .B(n25211), .C(reg_file[1124]), .D(
        n25222), .Y(n31424) );
  NAND3X1 U18700 ( .A(n31433), .B(n31434), .C(n31435), .Y(n31422) );
  NOR2X1 U18701 ( .A(n31436), .B(n31437), .Y(n31435) );
  OAI22X1 U18702 ( .A(n25232), .B(n31438), .C(n25242), .D(n31439), .Y(n31437)
         );
  OAI22X1 U18703 ( .A(n25253), .B(n31440), .C(n25263), .D(n31441), .Y(n31436)
         );
  AOI22X1 U18704 ( .A(reg_file[612]), .B(n25274), .C(reg_file[740]), .D(n25285), .Y(n31434) );
  AOI22X1 U18705 ( .A(reg_file[868]), .B(n25295), .C(reg_file[996]), .D(n25306), .Y(n31433) );
  NOR2X1 U18706 ( .A(n31442), .B(n31443), .Y(n31420) );
  NAND3X1 U18707 ( .A(n31444), .B(n31445), .C(n31446), .Y(n31443) );
  NOR2X1 U18708 ( .A(n31447), .B(n31448), .Y(n31446) );
  OAI22X1 U18709 ( .A(n25316), .B(n31449), .C(n25326), .D(n31450), .Y(n31448)
         );
  OAI22X1 U18710 ( .A(n25337), .B(n31451), .C(n25347), .D(n31452), .Y(n31447)
         );
  AOI22X1 U18711 ( .A(reg_file[3556]), .B(n25358), .C(reg_file[3428]), .D(
        n25369), .Y(n31445) );
  AOI22X1 U18712 ( .A(reg_file[3300]), .B(n25379), .C(reg_file[3172]), .D(
        n25390), .Y(n31444) );
  NAND3X1 U18713 ( .A(n31453), .B(n31454), .C(n31455), .Y(n31442) );
  NOR2X1 U18714 ( .A(n31456), .B(n31457), .Y(n31455) );
  OAI22X1 U18715 ( .A(n25400), .B(n31458), .C(n25410), .D(n31459), .Y(n31457)
         );
  OAI22X1 U18716 ( .A(n25421), .B(n31460), .C(n25431), .D(n31461), .Y(n31456)
         );
  AOI22X1 U18717 ( .A(reg_file[2532]), .B(n25442), .C(reg_file[2404]), .D(
        n25453), .Y(n31454) );
  AOI22X1 U18718 ( .A(reg_file[2276]), .B(n25463), .C(reg_file[2148]), .D(
        n25474), .Y(n31453) );
  AOI21X1 U18719 ( .A(n31462), .B(n31463), .C(n25137), .Y(rd2data1040_0_) );
  INVX1 U18720 ( .A(rd2en), .Y(n26097) );
  NOR2X1 U18721 ( .A(n31464), .B(n31465), .Y(n31463) );
  NAND3X1 U18722 ( .A(n31466), .B(n31467), .C(n31468), .Y(n31465) );
  NOR2X1 U18723 ( .A(n31469), .B(n31470), .Y(n31468) );
  OAI22X1 U18724 ( .A(n25148), .B(n31471), .C(n25158), .D(n31472), .Y(n31470)
         );
  NAND2X1 U18725 ( .A(n31473), .B(n31474), .Y(n26107) );
  NAND2X1 U18726 ( .A(n31475), .B(n31474), .Y(n26105) );
  OAI22X1 U18727 ( .A(n25169), .B(n31476), .C(n25179), .D(n31477), .Y(n31469)
         );
  NAND2X1 U18728 ( .A(n31473), .B(n31478), .Y(n26111) );
  NAND2X1 U18729 ( .A(n31475), .B(n31478), .Y(n26109) );
  AOI22X1 U18730 ( .A(reg_file[1408]), .B(n25190), .C(reg_file[1280]), .D(
        n25201), .Y(n31467) );
  AND2X1 U18731 ( .A(n31475), .B(n31479), .Y(n26114) );
  AND2X1 U18732 ( .A(n31473), .B(n31479), .Y(n26113) );
  AOI22X1 U18733 ( .A(reg_file[1152]), .B(n25211), .C(reg_file[1024]), .D(
        n25222), .Y(n31466) );
  AND2X1 U18734 ( .A(n31475), .B(n31480), .Y(n26116) );
  INVX1 U18735 ( .A(n31481), .Y(n31475) );
  NAND3X1 U18736 ( .A(n31482), .B(n31483), .C(rd2addr[3]), .Y(n31481) );
  AND2X1 U18737 ( .A(n31473), .B(n31480), .Y(n26115) );
  INVX1 U18738 ( .A(n31484), .Y(n31473) );
  NAND3X1 U18739 ( .A(rd2addr[0]), .B(n31483), .C(rd2addr[3]), .Y(n31484) );
  NAND3X1 U18740 ( .A(n31485), .B(n31486), .C(n31487), .Y(n31464) );
  NOR2X1 U18741 ( .A(n31488), .B(n31489), .Y(n31487) );
  OAI22X1 U18742 ( .A(n25232), .B(n31490), .C(n25242), .D(n31491), .Y(n31489)
         );
  NAND2X1 U18743 ( .A(n31479), .B(n31492), .Y(n26124) );
  NAND2X1 U18744 ( .A(n31479), .B(n31493), .Y(n26122) );
  OAI22X1 U18745 ( .A(n25253), .B(n31494), .C(n25263), .D(n31495), .Y(n31488)
         );
  NAND2X1 U18746 ( .A(n31480), .B(n31492), .Y(n26128) );
  NAND2X1 U18747 ( .A(n31493), .B(n31480), .Y(n26126) );
  AOI22X1 U18748 ( .A(reg_file[512]), .B(n25274), .C(reg_file[640]), .D(n25285), .Y(n31486) );
  AND2X1 U18749 ( .A(n31474), .B(n31493), .Y(n26131) );
  AND2X1 U18750 ( .A(n31474), .B(n31492), .Y(n26130) );
  AOI22X1 U18751 ( .A(reg_file[768]), .B(n25295), .C(reg_file[896]), .D(n25306), .Y(n31485) );
  AND2X1 U18752 ( .A(n31478), .B(n31493), .Y(n26133) );
  INVX1 U18753 ( .A(n31496), .Y(n31493) );
  NAND3X1 U18754 ( .A(n31497), .B(n31483), .C(rd2addr[0]), .Y(n31496) );
  AND2X1 U18755 ( .A(n31478), .B(n31492), .Y(n26132) );
  INVX1 U18756 ( .A(n31498), .Y(n31492) );
  NAND3X1 U18757 ( .A(n31497), .B(n31483), .C(n31482), .Y(n31498) );
  INVX1 U18758 ( .A(rd2addr[4]), .Y(n31483) );
  NOR2X1 U18759 ( .A(n31499), .B(n31500), .Y(n31462) );
  NAND3X1 U18760 ( .A(n31501), .B(n31502), .C(n31503), .Y(n31500) );
  NOR2X1 U18761 ( .A(n31504), .B(n31505), .Y(n31503) );
  OAI22X1 U18762 ( .A(n25316), .B(n31506), .C(n25326), .D(n31507), .Y(n31505)
         );
  NAND2X1 U18763 ( .A(n31508), .B(n31474), .Y(n26143) );
  NAND2X1 U18764 ( .A(n31509), .B(n31474), .Y(n26141) );
  OAI22X1 U18765 ( .A(n25337), .B(n31510), .C(n25347), .D(n31511), .Y(n31504)
         );
  NAND2X1 U18766 ( .A(n31508), .B(n31478), .Y(n26147) );
  NAND2X1 U18767 ( .A(n31509), .B(n31478), .Y(n26145) );
  AOI22X1 U18768 ( .A(reg_file[3456]), .B(n25358), .C(reg_file[3328]), .D(
        n25369), .Y(n31502) );
  AND2X1 U18769 ( .A(n31509), .B(n31479), .Y(n26150) );
  AND2X1 U18770 ( .A(n31508), .B(n31479), .Y(n26149) );
  AOI22X1 U18771 ( .A(reg_file[3200]), .B(n25379), .C(reg_file[3072]), .D(
        n25390), .Y(n31501) );
  AND2X1 U18772 ( .A(n31509), .B(n31480), .Y(n26152) );
  INVX1 U18773 ( .A(n31512), .Y(n31509) );
  NAND3X1 U18774 ( .A(rd2addr[3]), .B(n31482), .C(rd2addr[4]), .Y(n31512) );
  AND2X1 U18775 ( .A(n31508), .B(n31480), .Y(n26151) );
  INVX1 U18776 ( .A(n31513), .Y(n31508) );
  NAND3X1 U18777 ( .A(rd2addr[3]), .B(rd2addr[0]), .C(rd2addr[4]), .Y(n31513)
         );
  NAND3X1 U18778 ( .A(n31514), .B(n31515), .C(n31516), .Y(n31499) );
  NOR2X1 U18779 ( .A(n31517), .B(n31518), .Y(n31516) );
  OAI22X1 U18780 ( .A(n25400), .B(n31519), .C(n25410), .D(n31520), .Y(n31518)
         );
  NAND2X1 U18781 ( .A(n31521), .B(n31474), .Y(n26160) );
  NAND2X1 U18782 ( .A(n31522), .B(n31474), .Y(n26158) );
  AND2X1 U18783 ( .A(rd2addr[2]), .B(n31523), .Y(n31474) );
  OAI22X1 U18784 ( .A(n25421), .B(n31524), .C(n25431), .D(n31525), .Y(n31517)
         );
  NAND2X1 U18785 ( .A(n31521), .B(n31478), .Y(n26164) );
  NAND2X1 U18786 ( .A(n31522), .B(n31478), .Y(n26162) );
  AND2X1 U18787 ( .A(rd2addr[2]), .B(rd2addr[1]), .Y(n31478) );
  AOI22X1 U18788 ( .A(reg_file[2432]), .B(n25442), .C(reg_file[2304]), .D(
        n25453), .Y(n31515) );
  AND2X1 U18789 ( .A(n31522), .B(n31479), .Y(n26167) );
  AND2X1 U18790 ( .A(n31521), .B(n31479), .Y(n26166) );
  NOR2X1 U18791 ( .A(n31523), .B(rd2addr[2]), .Y(n31479) );
  INVX1 U18792 ( .A(rd2addr[1]), .Y(n31523) );
  AOI22X1 U18793 ( .A(reg_file[2176]), .B(n25463), .C(reg_file[2048]), .D(
        n25474), .Y(n31514) );
  AND2X1 U18794 ( .A(n31522), .B(n31480), .Y(n26169) );
  INVX1 U18795 ( .A(n31526), .Y(n31522) );
  NAND3X1 U18796 ( .A(n31482), .B(n31497), .C(rd2addr[4]), .Y(n31526) );
  INVX1 U18797 ( .A(rd2addr[0]), .Y(n31482) );
  AND2X1 U18798 ( .A(n31521), .B(n31480), .Y(n26168) );
  NOR2X1 U18799 ( .A(rd2addr[1]), .B(rd2addr[2]), .Y(n31480) );
  INVX1 U18800 ( .A(n31527), .Y(n31521) );
  NAND3X1 U18801 ( .A(rd2addr[0]), .B(n31497), .C(rd2addr[4]), .Y(n31527) );
  INVX1 U18802 ( .A(rd2addr[3]), .Y(n31497) );
  AOI21X1 U18803 ( .A(n31528), .B(n31529), .C(n25494), .Y(rd1data1033_9_) );
  NOR2X1 U18804 ( .A(n31531), .B(n31532), .Y(n31529) );
  NAND3X1 U18805 ( .A(n31533), .B(n31534), .C(n31535), .Y(n31532) );
  NOR2X1 U18806 ( .A(n31536), .B(n31537), .Y(n31535) );
  OAI22X1 U18807 ( .A(n26106), .B(n25505), .C(n26108), .D(n25515), .Y(n31537)
         );
  OAI22X1 U18808 ( .A(n26110), .B(n25526), .C(n26112), .D(n25536), .Y(n31536)
         );
  AOI22X1 U18809 ( .A(n25547), .B(reg_file[1417]), .C(n25558), .D(
        reg_file[1289]), .Y(n31534) );
  AOI22X1 U18810 ( .A(n25569), .B(reg_file[1161]), .C(n25580), .D(
        reg_file[1033]), .Y(n31533) );
  NAND3X1 U18811 ( .A(n31546), .B(n31547), .C(n31548), .Y(n31531) );
  NOR2X1 U18812 ( .A(n31549), .B(n31550), .Y(n31548) );
  OAI22X1 U18813 ( .A(n26123), .B(n25591), .C(n26125), .D(n25601), .Y(n31550)
         );
  OAI22X1 U18814 ( .A(n26127), .B(n25612), .C(n26129), .D(n25622), .Y(n31549)
         );
  AOI22X1 U18815 ( .A(n25633), .B(reg_file[521]), .C(n25644), .D(reg_file[649]), .Y(n31547) );
  AOI22X1 U18816 ( .A(n25655), .B(reg_file[777]), .C(n25666), .D(reg_file[905]), .Y(n31546) );
  NOR2X1 U18817 ( .A(n31559), .B(n31560), .Y(n31528) );
  NAND3X1 U18818 ( .A(n31561), .B(n31562), .C(n31563), .Y(n31560) );
  NOR2X1 U18819 ( .A(n31564), .B(n31565), .Y(n31563) );
  OAI22X1 U18820 ( .A(n26142), .B(n25677), .C(n26144), .D(n25687), .Y(n31565)
         );
  OAI22X1 U18821 ( .A(n26146), .B(n25698), .C(n26148), .D(n25708), .Y(n31564)
         );
  AOI22X1 U18822 ( .A(n25719), .B(reg_file[3465]), .C(n25730), .D(
        reg_file[3337]), .Y(n31562) );
  AOI22X1 U18823 ( .A(n25741), .B(reg_file[3209]), .C(n25752), .D(
        reg_file[3081]), .Y(n31561) );
  NAND3X1 U18824 ( .A(n31574), .B(n31575), .C(n31576), .Y(n31559) );
  NOR2X1 U18825 ( .A(n31577), .B(n31578), .Y(n31576) );
  OAI22X1 U18826 ( .A(n26159), .B(n25763), .C(n26161), .D(n25773), .Y(n31578)
         );
  OAI22X1 U18827 ( .A(n26163), .B(n25784), .C(n26165), .D(n25794), .Y(n31577)
         );
  AOI22X1 U18828 ( .A(n25805), .B(reg_file[2441]), .C(n25816), .D(
        reg_file[2313]), .Y(n31575) );
  AOI22X1 U18829 ( .A(n25827), .B(reg_file[2185]), .C(n25838), .D(
        reg_file[2057]), .Y(n31574) );
  AOI21X1 U18830 ( .A(n31587), .B(n31588), .C(n25494), .Y(rd1data1033_99_) );
  NOR2X1 U18831 ( .A(n31589), .B(n31590), .Y(n31588) );
  NAND3X1 U18832 ( .A(n31591), .B(n31592), .C(n31593), .Y(n31590) );
  NOR2X1 U18833 ( .A(n31594), .B(n31595), .Y(n31593) );
  OAI22X1 U18834 ( .A(n26179), .B(n25505), .C(n26180), .D(n25515), .Y(n31595)
         );
  OAI22X1 U18835 ( .A(n26181), .B(n25526), .C(n26182), .D(n25536), .Y(n31594)
         );
  AOI22X1 U18836 ( .A(n25547), .B(reg_file[1507]), .C(n25558), .D(
        reg_file[1379]), .Y(n31592) );
  AOI22X1 U18837 ( .A(n25569), .B(reg_file[1251]), .C(n25580), .D(
        reg_file[1123]), .Y(n31591) );
  NAND3X1 U18838 ( .A(n31596), .B(n31597), .C(n31598), .Y(n31589) );
  NOR2X1 U18839 ( .A(n31599), .B(n31600), .Y(n31598) );
  OAI22X1 U18840 ( .A(n26188), .B(n25591), .C(n26189), .D(n25601), .Y(n31600)
         );
  OAI22X1 U18841 ( .A(n26190), .B(n25612), .C(n26191), .D(n25622), .Y(n31599)
         );
  AOI22X1 U18842 ( .A(n25633), .B(reg_file[611]), .C(n25644), .D(reg_file[739]), .Y(n31597) );
  AOI22X1 U18843 ( .A(n25655), .B(reg_file[867]), .C(n25666), .D(reg_file[995]), .Y(n31596) );
  NOR2X1 U18844 ( .A(n31601), .B(n31602), .Y(n31587) );
  NAND3X1 U18845 ( .A(n31603), .B(n31604), .C(n31605), .Y(n31602) );
  NOR2X1 U18846 ( .A(n31606), .B(n31607), .Y(n31605) );
  OAI22X1 U18847 ( .A(n26199), .B(n25677), .C(n26200), .D(n25687), .Y(n31607)
         );
  OAI22X1 U18848 ( .A(n26201), .B(n25698), .C(n26202), .D(n25708), .Y(n31606)
         );
  AOI22X1 U18849 ( .A(n25719), .B(reg_file[3555]), .C(n25730), .D(
        reg_file[3427]), .Y(n31604) );
  AOI22X1 U18850 ( .A(n25741), .B(reg_file[3299]), .C(n25752), .D(
        reg_file[3171]), .Y(n31603) );
  NAND3X1 U18851 ( .A(n31608), .B(n31609), .C(n31610), .Y(n31601) );
  NOR2X1 U18852 ( .A(n31611), .B(n31612), .Y(n31610) );
  OAI22X1 U18853 ( .A(n26208), .B(n25763), .C(n26209), .D(n25773), .Y(n31612)
         );
  OAI22X1 U18854 ( .A(n26210), .B(n25784), .C(n26211), .D(n25794), .Y(n31611)
         );
  AOI22X1 U18855 ( .A(n25805), .B(reg_file[2531]), .C(n25816), .D(
        reg_file[2403]), .Y(n31609) );
  AOI22X1 U18856 ( .A(n25827), .B(reg_file[2275]), .C(n25838), .D(
        reg_file[2147]), .Y(n31608) );
  AOI21X1 U18857 ( .A(n31613), .B(n31614), .C(n25494), .Y(rd1data1033_98_) );
  NOR2X1 U18858 ( .A(n31615), .B(n31616), .Y(n31614) );
  NAND3X1 U18859 ( .A(n31617), .B(n31618), .C(n31619), .Y(n31616) );
  NOR2X1 U18860 ( .A(n31620), .B(n31621), .Y(n31619) );
  OAI22X1 U18861 ( .A(n26221), .B(n25505), .C(n26222), .D(n25515), .Y(n31621)
         );
  OAI22X1 U18862 ( .A(n26223), .B(n25526), .C(n26224), .D(n25536), .Y(n31620)
         );
  AOI22X1 U18863 ( .A(n25547), .B(reg_file[1506]), .C(n25558), .D(
        reg_file[1378]), .Y(n31618) );
  AOI22X1 U18864 ( .A(n25569), .B(reg_file[1250]), .C(n25580), .D(
        reg_file[1122]), .Y(n31617) );
  NAND3X1 U18865 ( .A(n31622), .B(n31623), .C(n31624), .Y(n31615) );
  NOR2X1 U18866 ( .A(n31625), .B(n31626), .Y(n31624) );
  OAI22X1 U18867 ( .A(n26230), .B(n25591), .C(n26231), .D(n25601), .Y(n31626)
         );
  OAI22X1 U18868 ( .A(n26232), .B(n25612), .C(n26233), .D(n25622), .Y(n31625)
         );
  AOI22X1 U18869 ( .A(n25633), .B(reg_file[610]), .C(n25644), .D(reg_file[738]), .Y(n31623) );
  AOI22X1 U18870 ( .A(n25655), .B(reg_file[866]), .C(n25666), .D(reg_file[994]), .Y(n31622) );
  NOR2X1 U18871 ( .A(n31627), .B(n31628), .Y(n31613) );
  NAND3X1 U18872 ( .A(n31629), .B(n31630), .C(n31631), .Y(n31628) );
  NOR2X1 U18873 ( .A(n31632), .B(n31633), .Y(n31631) );
  OAI22X1 U18874 ( .A(n26241), .B(n25677), .C(n26242), .D(n25687), .Y(n31633)
         );
  OAI22X1 U18875 ( .A(n26243), .B(n25698), .C(n26244), .D(n25708), .Y(n31632)
         );
  AOI22X1 U18876 ( .A(n25719), .B(reg_file[3554]), .C(n25730), .D(
        reg_file[3426]), .Y(n31630) );
  AOI22X1 U18877 ( .A(n25741), .B(reg_file[3298]), .C(n25752), .D(
        reg_file[3170]), .Y(n31629) );
  NAND3X1 U18878 ( .A(n31634), .B(n31635), .C(n31636), .Y(n31627) );
  NOR2X1 U18879 ( .A(n31637), .B(n31638), .Y(n31636) );
  OAI22X1 U18880 ( .A(n26250), .B(n25763), .C(n26251), .D(n25773), .Y(n31638)
         );
  OAI22X1 U18881 ( .A(n26252), .B(n25784), .C(n26253), .D(n25794), .Y(n31637)
         );
  AOI22X1 U18882 ( .A(n25805), .B(reg_file[2530]), .C(n25816), .D(
        reg_file[2402]), .Y(n31635) );
  AOI22X1 U18883 ( .A(n25827), .B(reg_file[2274]), .C(n25838), .D(
        reg_file[2146]), .Y(n31634) );
  AOI21X1 U18884 ( .A(n31639), .B(n31640), .C(n25494), .Y(rd1data1033_97_) );
  NOR2X1 U18885 ( .A(n31641), .B(n31642), .Y(n31640) );
  NAND3X1 U18886 ( .A(n31643), .B(n31644), .C(n31645), .Y(n31642) );
  NOR2X1 U18887 ( .A(n31646), .B(n31647), .Y(n31645) );
  OAI22X1 U18888 ( .A(n26263), .B(n25505), .C(n26264), .D(n25515), .Y(n31647)
         );
  OAI22X1 U18889 ( .A(n26265), .B(n25526), .C(n26266), .D(n25536), .Y(n31646)
         );
  AOI22X1 U18890 ( .A(n25547), .B(reg_file[1505]), .C(n25558), .D(
        reg_file[1377]), .Y(n31644) );
  AOI22X1 U18891 ( .A(n25569), .B(reg_file[1249]), .C(n25580), .D(
        reg_file[1121]), .Y(n31643) );
  NAND3X1 U18892 ( .A(n31648), .B(n31649), .C(n31650), .Y(n31641) );
  NOR2X1 U18893 ( .A(n31651), .B(n31652), .Y(n31650) );
  OAI22X1 U18894 ( .A(n26272), .B(n25591), .C(n26273), .D(n25601), .Y(n31652)
         );
  OAI22X1 U18895 ( .A(n26274), .B(n25612), .C(n26275), .D(n25622), .Y(n31651)
         );
  AOI22X1 U18896 ( .A(n25633), .B(reg_file[609]), .C(n25644), .D(reg_file[737]), .Y(n31649) );
  AOI22X1 U18897 ( .A(n25655), .B(reg_file[865]), .C(n25666), .D(reg_file[993]), .Y(n31648) );
  NOR2X1 U18898 ( .A(n31653), .B(n31654), .Y(n31639) );
  NAND3X1 U18899 ( .A(n31655), .B(n31656), .C(n31657), .Y(n31654) );
  NOR2X1 U18900 ( .A(n31658), .B(n31659), .Y(n31657) );
  OAI22X1 U18901 ( .A(n26283), .B(n25677), .C(n26284), .D(n25687), .Y(n31659)
         );
  OAI22X1 U18902 ( .A(n26285), .B(n25698), .C(n26286), .D(n25708), .Y(n31658)
         );
  AOI22X1 U18903 ( .A(n25719), .B(reg_file[3553]), .C(n25730), .D(
        reg_file[3425]), .Y(n31656) );
  AOI22X1 U18904 ( .A(n25741), .B(reg_file[3297]), .C(n25752), .D(
        reg_file[3169]), .Y(n31655) );
  NAND3X1 U18905 ( .A(n31660), .B(n31661), .C(n31662), .Y(n31653) );
  NOR2X1 U18906 ( .A(n31663), .B(n31664), .Y(n31662) );
  OAI22X1 U18907 ( .A(n26292), .B(n25763), .C(n26293), .D(n25773), .Y(n31664)
         );
  OAI22X1 U18908 ( .A(n26294), .B(n25784), .C(n26295), .D(n25794), .Y(n31663)
         );
  AOI22X1 U18909 ( .A(n25805), .B(reg_file[2529]), .C(n25816), .D(
        reg_file[2401]), .Y(n31661) );
  AOI22X1 U18910 ( .A(n25827), .B(reg_file[2273]), .C(n25838), .D(
        reg_file[2145]), .Y(n31660) );
  AOI21X1 U18911 ( .A(n31665), .B(n31666), .C(n25494), .Y(rd1data1033_96_) );
  NOR2X1 U18912 ( .A(n31667), .B(n31668), .Y(n31666) );
  NAND3X1 U18913 ( .A(n31669), .B(n31670), .C(n31671), .Y(n31668) );
  NOR2X1 U18914 ( .A(n31672), .B(n31673), .Y(n31671) );
  OAI22X1 U18915 ( .A(n26305), .B(n25505), .C(n26306), .D(n25515), .Y(n31673)
         );
  OAI22X1 U18916 ( .A(n26307), .B(n25526), .C(n26308), .D(n25536), .Y(n31672)
         );
  AOI22X1 U18917 ( .A(n25547), .B(reg_file[1504]), .C(n25558), .D(
        reg_file[1376]), .Y(n31670) );
  AOI22X1 U18918 ( .A(n25569), .B(reg_file[1248]), .C(n25580), .D(
        reg_file[1120]), .Y(n31669) );
  NAND3X1 U18919 ( .A(n31674), .B(n31675), .C(n31676), .Y(n31667) );
  NOR2X1 U18920 ( .A(n31677), .B(n31678), .Y(n31676) );
  OAI22X1 U18921 ( .A(n26314), .B(n25591), .C(n26315), .D(n25601), .Y(n31678)
         );
  OAI22X1 U18922 ( .A(n26316), .B(n25612), .C(n26317), .D(n25622), .Y(n31677)
         );
  AOI22X1 U18923 ( .A(n25633), .B(reg_file[608]), .C(n25644), .D(reg_file[736]), .Y(n31675) );
  AOI22X1 U18924 ( .A(n25655), .B(reg_file[864]), .C(n25666), .D(reg_file[992]), .Y(n31674) );
  NOR2X1 U18925 ( .A(n31679), .B(n31680), .Y(n31665) );
  NAND3X1 U18926 ( .A(n31681), .B(n31682), .C(n31683), .Y(n31680) );
  NOR2X1 U18927 ( .A(n31684), .B(n31685), .Y(n31683) );
  OAI22X1 U18928 ( .A(n26325), .B(n25677), .C(n26326), .D(n25687), .Y(n31685)
         );
  OAI22X1 U18929 ( .A(n26327), .B(n25698), .C(n26328), .D(n25708), .Y(n31684)
         );
  AOI22X1 U18930 ( .A(n25719), .B(reg_file[3552]), .C(n25730), .D(
        reg_file[3424]), .Y(n31682) );
  AOI22X1 U18931 ( .A(n25741), .B(reg_file[3296]), .C(n25752), .D(
        reg_file[3168]), .Y(n31681) );
  NAND3X1 U18932 ( .A(n31686), .B(n31687), .C(n31688), .Y(n31679) );
  NOR2X1 U18933 ( .A(n31689), .B(n31690), .Y(n31688) );
  OAI22X1 U18934 ( .A(n26334), .B(n25763), .C(n26335), .D(n25773), .Y(n31690)
         );
  OAI22X1 U18935 ( .A(n26336), .B(n25784), .C(n26337), .D(n25794), .Y(n31689)
         );
  AOI22X1 U18936 ( .A(n25805), .B(reg_file[2528]), .C(n25816), .D(
        reg_file[2400]), .Y(n31687) );
  AOI22X1 U18937 ( .A(n25827), .B(reg_file[2272]), .C(n25838), .D(
        reg_file[2144]), .Y(n31686) );
  AOI21X1 U18938 ( .A(n31691), .B(n31692), .C(n25494), .Y(rd1data1033_95_) );
  NOR2X1 U18939 ( .A(n31693), .B(n31694), .Y(n31692) );
  NAND3X1 U18940 ( .A(n31695), .B(n31696), .C(n31697), .Y(n31694) );
  NOR2X1 U18941 ( .A(n31698), .B(n31699), .Y(n31697) );
  OAI22X1 U18942 ( .A(n26347), .B(n25505), .C(n26348), .D(n25515), .Y(n31699)
         );
  OAI22X1 U18943 ( .A(n26349), .B(n25526), .C(n26350), .D(n25536), .Y(n31698)
         );
  AOI22X1 U18944 ( .A(n25547), .B(reg_file[1503]), .C(n25558), .D(
        reg_file[1375]), .Y(n31696) );
  AOI22X1 U18945 ( .A(n25569), .B(reg_file[1247]), .C(n25580), .D(
        reg_file[1119]), .Y(n31695) );
  NAND3X1 U18946 ( .A(n31700), .B(n31701), .C(n31702), .Y(n31693) );
  NOR2X1 U18947 ( .A(n31703), .B(n31704), .Y(n31702) );
  OAI22X1 U18948 ( .A(n26356), .B(n25591), .C(n26357), .D(n25601), .Y(n31704)
         );
  OAI22X1 U18949 ( .A(n26358), .B(n25612), .C(n26359), .D(n25622), .Y(n31703)
         );
  AOI22X1 U18950 ( .A(n25633), .B(reg_file[607]), .C(n25644), .D(reg_file[735]), .Y(n31701) );
  AOI22X1 U18951 ( .A(n25655), .B(reg_file[863]), .C(n25666), .D(reg_file[991]), .Y(n31700) );
  NOR2X1 U18952 ( .A(n31705), .B(n31706), .Y(n31691) );
  NAND3X1 U18953 ( .A(n31707), .B(n31708), .C(n31709), .Y(n31706) );
  NOR2X1 U18954 ( .A(n31710), .B(n31711), .Y(n31709) );
  OAI22X1 U18955 ( .A(n26367), .B(n25677), .C(n26368), .D(n25687), .Y(n31711)
         );
  OAI22X1 U18956 ( .A(n26369), .B(n25698), .C(n26370), .D(n25708), .Y(n31710)
         );
  AOI22X1 U18957 ( .A(n25719), .B(reg_file[3551]), .C(n25730), .D(
        reg_file[3423]), .Y(n31708) );
  AOI22X1 U18958 ( .A(n25741), .B(reg_file[3295]), .C(n25752), .D(
        reg_file[3167]), .Y(n31707) );
  NAND3X1 U18959 ( .A(n31712), .B(n31713), .C(n31714), .Y(n31705) );
  NOR2X1 U18960 ( .A(n31715), .B(n31716), .Y(n31714) );
  OAI22X1 U18961 ( .A(n26376), .B(n25763), .C(n26377), .D(n25773), .Y(n31716)
         );
  OAI22X1 U18962 ( .A(n26378), .B(n25784), .C(n26379), .D(n25794), .Y(n31715)
         );
  AOI22X1 U18963 ( .A(n25805), .B(reg_file[2527]), .C(n25816), .D(
        reg_file[2399]), .Y(n31713) );
  AOI22X1 U18964 ( .A(n25827), .B(reg_file[2271]), .C(n25838), .D(
        reg_file[2143]), .Y(n31712) );
  AOI21X1 U18965 ( .A(n31717), .B(n31718), .C(n25494), .Y(rd1data1033_94_) );
  NOR2X1 U18966 ( .A(n31719), .B(n31720), .Y(n31718) );
  NAND3X1 U18967 ( .A(n31721), .B(n31722), .C(n31723), .Y(n31720) );
  NOR2X1 U18968 ( .A(n31724), .B(n31725), .Y(n31723) );
  OAI22X1 U18969 ( .A(n26389), .B(n25505), .C(n26390), .D(n25515), .Y(n31725)
         );
  OAI22X1 U18970 ( .A(n26391), .B(n25526), .C(n26392), .D(n25536), .Y(n31724)
         );
  AOI22X1 U18971 ( .A(n25547), .B(reg_file[1502]), .C(n25558), .D(
        reg_file[1374]), .Y(n31722) );
  AOI22X1 U18972 ( .A(n25569), .B(reg_file[1246]), .C(n25580), .D(
        reg_file[1118]), .Y(n31721) );
  NAND3X1 U18973 ( .A(n31726), .B(n31727), .C(n31728), .Y(n31719) );
  NOR2X1 U18974 ( .A(n31729), .B(n31730), .Y(n31728) );
  OAI22X1 U18975 ( .A(n26398), .B(n25591), .C(n26399), .D(n25601), .Y(n31730)
         );
  OAI22X1 U18976 ( .A(n26400), .B(n25612), .C(n26401), .D(n25622), .Y(n31729)
         );
  AOI22X1 U18977 ( .A(n25633), .B(reg_file[606]), .C(n25644), .D(reg_file[734]), .Y(n31727) );
  AOI22X1 U18978 ( .A(n25655), .B(reg_file[862]), .C(n25666), .D(reg_file[990]), .Y(n31726) );
  NOR2X1 U18979 ( .A(n31731), .B(n31732), .Y(n31717) );
  NAND3X1 U18980 ( .A(n31733), .B(n31734), .C(n31735), .Y(n31732) );
  NOR2X1 U18981 ( .A(n31736), .B(n31737), .Y(n31735) );
  OAI22X1 U18982 ( .A(n26409), .B(n25677), .C(n26410), .D(n25687), .Y(n31737)
         );
  OAI22X1 U18983 ( .A(n26411), .B(n25698), .C(n26412), .D(n25708), .Y(n31736)
         );
  AOI22X1 U18984 ( .A(n25719), .B(reg_file[3550]), .C(n25730), .D(
        reg_file[3422]), .Y(n31734) );
  AOI22X1 U18985 ( .A(n25741), .B(reg_file[3294]), .C(n25752), .D(
        reg_file[3166]), .Y(n31733) );
  NAND3X1 U18986 ( .A(n31738), .B(n31739), .C(n31740), .Y(n31731) );
  NOR2X1 U18987 ( .A(n31741), .B(n31742), .Y(n31740) );
  OAI22X1 U18988 ( .A(n26418), .B(n25763), .C(n26419), .D(n25773), .Y(n31742)
         );
  OAI22X1 U18989 ( .A(n26420), .B(n25784), .C(n26421), .D(n25794), .Y(n31741)
         );
  AOI22X1 U18990 ( .A(n25805), .B(reg_file[2526]), .C(n25816), .D(
        reg_file[2398]), .Y(n31739) );
  AOI22X1 U18991 ( .A(n25827), .B(reg_file[2270]), .C(n25838), .D(
        reg_file[2142]), .Y(n31738) );
  AOI21X1 U18992 ( .A(n31743), .B(n31744), .C(n25494), .Y(rd1data1033_93_) );
  NOR2X1 U18993 ( .A(n31745), .B(n31746), .Y(n31744) );
  NAND3X1 U18994 ( .A(n31747), .B(n31748), .C(n31749), .Y(n31746) );
  NOR2X1 U18995 ( .A(n31750), .B(n31751), .Y(n31749) );
  OAI22X1 U18996 ( .A(n26431), .B(n25505), .C(n26432), .D(n25515), .Y(n31751)
         );
  OAI22X1 U18997 ( .A(n26433), .B(n25526), .C(n26434), .D(n25536), .Y(n31750)
         );
  AOI22X1 U18998 ( .A(n25547), .B(reg_file[1501]), .C(n25558), .D(
        reg_file[1373]), .Y(n31748) );
  AOI22X1 U18999 ( .A(n25569), .B(reg_file[1245]), .C(n25580), .D(
        reg_file[1117]), .Y(n31747) );
  NAND3X1 U19000 ( .A(n31752), .B(n31753), .C(n31754), .Y(n31745) );
  NOR2X1 U19001 ( .A(n31755), .B(n31756), .Y(n31754) );
  OAI22X1 U19002 ( .A(n26440), .B(n25591), .C(n26441), .D(n25601), .Y(n31756)
         );
  OAI22X1 U19003 ( .A(n26442), .B(n25612), .C(n26443), .D(n25622), .Y(n31755)
         );
  AOI22X1 U19004 ( .A(n25633), .B(reg_file[605]), .C(n25644), .D(reg_file[733]), .Y(n31753) );
  AOI22X1 U19005 ( .A(n25655), .B(reg_file[861]), .C(n25666), .D(reg_file[989]), .Y(n31752) );
  NOR2X1 U19006 ( .A(n31757), .B(n31758), .Y(n31743) );
  NAND3X1 U19007 ( .A(n31759), .B(n31760), .C(n31761), .Y(n31758) );
  NOR2X1 U19008 ( .A(n31762), .B(n31763), .Y(n31761) );
  OAI22X1 U19009 ( .A(n26451), .B(n25677), .C(n26452), .D(n25687), .Y(n31763)
         );
  OAI22X1 U19010 ( .A(n26453), .B(n25698), .C(n26454), .D(n25708), .Y(n31762)
         );
  AOI22X1 U19011 ( .A(n25719), .B(reg_file[3549]), .C(n25730), .D(
        reg_file[3421]), .Y(n31760) );
  AOI22X1 U19012 ( .A(n25741), .B(reg_file[3293]), .C(n25752), .D(
        reg_file[3165]), .Y(n31759) );
  NAND3X1 U19013 ( .A(n31764), .B(n31765), .C(n31766), .Y(n31757) );
  NOR2X1 U19014 ( .A(n31767), .B(n31768), .Y(n31766) );
  OAI22X1 U19015 ( .A(n26460), .B(n25763), .C(n26461), .D(n25773), .Y(n31768)
         );
  OAI22X1 U19016 ( .A(n26462), .B(n25784), .C(n26463), .D(n25794), .Y(n31767)
         );
  AOI22X1 U19017 ( .A(n25805), .B(reg_file[2525]), .C(n25816), .D(
        reg_file[2397]), .Y(n31765) );
  AOI22X1 U19018 ( .A(n25827), .B(reg_file[2269]), .C(n25838), .D(
        reg_file[2141]), .Y(n31764) );
  AOI21X1 U19019 ( .A(n31769), .B(n31770), .C(n25493), .Y(rd1data1033_92_) );
  NOR2X1 U19020 ( .A(n31771), .B(n31772), .Y(n31770) );
  NAND3X1 U19021 ( .A(n31773), .B(n31774), .C(n31775), .Y(n31772) );
  NOR2X1 U19022 ( .A(n31776), .B(n31777), .Y(n31775) );
  OAI22X1 U19023 ( .A(n26473), .B(n25504), .C(n26474), .D(n25515), .Y(n31777)
         );
  OAI22X1 U19024 ( .A(n26475), .B(n25525), .C(n26476), .D(n25536), .Y(n31776)
         );
  AOI22X1 U19025 ( .A(n25546), .B(reg_file[1500]), .C(n25557), .D(
        reg_file[1372]), .Y(n31774) );
  AOI22X1 U19026 ( .A(n25568), .B(reg_file[1244]), .C(n25579), .D(
        reg_file[1116]), .Y(n31773) );
  NAND3X1 U19027 ( .A(n31778), .B(n31779), .C(n31780), .Y(n31771) );
  NOR2X1 U19028 ( .A(n31781), .B(n31782), .Y(n31780) );
  OAI22X1 U19029 ( .A(n26482), .B(n25590), .C(n26483), .D(n25601), .Y(n31782)
         );
  OAI22X1 U19030 ( .A(n26484), .B(n25611), .C(n26485), .D(n25622), .Y(n31781)
         );
  AOI22X1 U19031 ( .A(n25632), .B(reg_file[604]), .C(n25643), .D(reg_file[732]), .Y(n31779) );
  AOI22X1 U19032 ( .A(n25654), .B(reg_file[860]), .C(n25665), .D(reg_file[988]), .Y(n31778) );
  NOR2X1 U19033 ( .A(n31783), .B(n31784), .Y(n31769) );
  NAND3X1 U19034 ( .A(n31785), .B(n31786), .C(n31787), .Y(n31784) );
  NOR2X1 U19035 ( .A(n31788), .B(n31789), .Y(n31787) );
  OAI22X1 U19036 ( .A(n26493), .B(n25676), .C(n26494), .D(n25687), .Y(n31789)
         );
  OAI22X1 U19037 ( .A(n26495), .B(n25697), .C(n26496), .D(n25708), .Y(n31788)
         );
  AOI22X1 U19038 ( .A(n25718), .B(reg_file[3548]), .C(n25729), .D(
        reg_file[3420]), .Y(n31786) );
  AOI22X1 U19039 ( .A(n25740), .B(reg_file[3292]), .C(n25751), .D(
        reg_file[3164]), .Y(n31785) );
  NAND3X1 U19040 ( .A(n31790), .B(n31791), .C(n31792), .Y(n31783) );
  NOR2X1 U19041 ( .A(n31793), .B(n31794), .Y(n31792) );
  OAI22X1 U19042 ( .A(n26502), .B(n25762), .C(n26503), .D(n25773), .Y(n31794)
         );
  OAI22X1 U19043 ( .A(n26504), .B(n25783), .C(n26505), .D(n25794), .Y(n31793)
         );
  AOI22X1 U19044 ( .A(n25804), .B(reg_file[2524]), .C(n25815), .D(
        reg_file[2396]), .Y(n31791) );
  AOI22X1 U19045 ( .A(n25826), .B(reg_file[2268]), .C(n25837), .D(
        reg_file[2140]), .Y(n31790) );
  AOI21X1 U19046 ( .A(n31795), .B(n31796), .C(n25493), .Y(rd1data1033_91_) );
  NOR2X1 U19047 ( .A(n31797), .B(n31798), .Y(n31796) );
  NAND3X1 U19048 ( .A(n31799), .B(n31800), .C(n31801), .Y(n31798) );
  NOR2X1 U19049 ( .A(n31802), .B(n31803), .Y(n31801) );
  OAI22X1 U19050 ( .A(n26515), .B(n25504), .C(n26516), .D(n25515), .Y(n31803)
         );
  OAI22X1 U19051 ( .A(n26517), .B(n25525), .C(n26518), .D(n25536), .Y(n31802)
         );
  AOI22X1 U19052 ( .A(n25546), .B(reg_file[1499]), .C(n25557), .D(
        reg_file[1371]), .Y(n31800) );
  AOI22X1 U19053 ( .A(n25568), .B(reg_file[1243]), .C(n25579), .D(
        reg_file[1115]), .Y(n31799) );
  NAND3X1 U19054 ( .A(n31804), .B(n31805), .C(n31806), .Y(n31797) );
  NOR2X1 U19055 ( .A(n31807), .B(n31808), .Y(n31806) );
  OAI22X1 U19056 ( .A(n26524), .B(n25590), .C(n26525), .D(n25601), .Y(n31808)
         );
  OAI22X1 U19057 ( .A(n26526), .B(n25611), .C(n26527), .D(n25622), .Y(n31807)
         );
  AOI22X1 U19058 ( .A(n25632), .B(reg_file[603]), .C(n25643), .D(reg_file[731]), .Y(n31805) );
  AOI22X1 U19059 ( .A(n25654), .B(reg_file[859]), .C(n25665), .D(reg_file[987]), .Y(n31804) );
  NOR2X1 U19060 ( .A(n31809), .B(n31810), .Y(n31795) );
  NAND3X1 U19061 ( .A(n31811), .B(n31812), .C(n31813), .Y(n31810) );
  NOR2X1 U19062 ( .A(n31814), .B(n31815), .Y(n31813) );
  OAI22X1 U19063 ( .A(n26535), .B(n25676), .C(n26536), .D(n25687), .Y(n31815)
         );
  OAI22X1 U19064 ( .A(n26537), .B(n25697), .C(n26538), .D(n25708), .Y(n31814)
         );
  AOI22X1 U19065 ( .A(n25718), .B(reg_file[3547]), .C(n25729), .D(
        reg_file[3419]), .Y(n31812) );
  AOI22X1 U19066 ( .A(n25740), .B(reg_file[3291]), .C(n25751), .D(
        reg_file[3163]), .Y(n31811) );
  NAND3X1 U19067 ( .A(n31816), .B(n31817), .C(n31818), .Y(n31809) );
  NOR2X1 U19068 ( .A(n31819), .B(n31820), .Y(n31818) );
  OAI22X1 U19069 ( .A(n26544), .B(n25762), .C(n26545), .D(n25773), .Y(n31820)
         );
  OAI22X1 U19070 ( .A(n26546), .B(n25783), .C(n26547), .D(n25794), .Y(n31819)
         );
  AOI22X1 U19071 ( .A(n25804), .B(reg_file[2523]), .C(n25815), .D(
        reg_file[2395]), .Y(n31817) );
  AOI22X1 U19072 ( .A(n25826), .B(reg_file[2267]), .C(n25837), .D(
        reg_file[2139]), .Y(n31816) );
  AOI21X1 U19073 ( .A(n31821), .B(n31822), .C(n25493), .Y(rd1data1033_90_) );
  NOR2X1 U19074 ( .A(n31823), .B(n31824), .Y(n31822) );
  NAND3X1 U19075 ( .A(n31825), .B(n31826), .C(n31827), .Y(n31824) );
  NOR2X1 U19076 ( .A(n31828), .B(n31829), .Y(n31827) );
  OAI22X1 U19077 ( .A(n26557), .B(n25504), .C(n26558), .D(n25515), .Y(n31829)
         );
  OAI22X1 U19078 ( .A(n26559), .B(n25525), .C(n26560), .D(n25536), .Y(n31828)
         );
  AOI22X1 U19079 ( .A(n25546), .B(reg_file[1498]), .C(n25557), .D(
        reg_file[1370]), .Y(n31826) );
  AOI22X1 U19080 ( .A(n25568), .B(reg_file[1242]), .C(n25579), .D(
        reg_file[1114]), .Y(n31825) );
  NAND3X1 U19081 ( .A(n31830), .B(n31831), .C(n31832), .Y(n31823) );
  NOR2X1 U19082 ( .A(n31833), .B(n31834), .Y(n31832) );
  OAI22X1 U19083 ( .A(n26566), .B(n25590), .C(n26567), .D(n25601), .Y(n31834)
         );
  OAI22X1 U19084 ( .A(n26568), .B(n25611), .C(n26569), .D(n25622), .Y(n31833)
         );
  AOI22X1 U19085 ( .A(n25632), .B(reg_file[602]), .C(n25643), .D(reg_file[730]), .Y(n31831) );
  AOI22X1 U19086 ( .A(n25654), .B(reg_file[858]), .C(n25665), .D(reg_file[986]), .Y(n31830) );
  NOR2X1 U19087 ( .A(n31835), .B(n31836), .Y(n31821) );
  NAND3X1 U19088 ( .A(n31837), .B(n31838), .C(n31839), .Y(n31836) );
  NOR2X1 U19089 ( .A(n31840), .B(n31841), .Y(n31839) );
  OAI22X1 U19090 ( .A(n26577), .B(n25676), .C(n26578), .D(n25687), .Y(n31841)
         );
  OAI22X1 U19091 ( .A(n26579), .B(n25697), .C(n26580), .D(n25708), .Y(n31840)
         );
  AOI22X1 U19092 ( .A(n25718), .B(reg_file[3546]), .C(n25729), .D(
        reg_file[3418]), .Y(n31838) );
  AOI22X1 U19093 ( .A(n25740), .B(reg_file[3290]), .C(n25751), .D(
        reg_file[3162]), .Y(n31837) );
  NAND3X1 U19094 ( .A(n31842), .B(n31843), .C(n31844), .Y(n31835) );
  NOR2X1 U19095 ( .A(n31845), .B(n31846), .Y(n31844) );
  OAI22X1 U19096 ( .A(n26586), .B(n25762), .C(n26587), .D(n25773), .Y(n31846)
         );
  OAI22X1 U19097 ( .A(n26588), .B(n25783), .C(n26589), .D(n25794), .Y(n31845)
         );
  AOI22X1 U19098 ( .A(n25804), .B(reg_file[2522]), .C(n25815), .D(
        reg_file[2394]), .Y(n31843) );
  AOI22X1 U19099 ( .A(n25826), .B(reg_file[2266]), .C(n25837), .D(
        reg_file[2138]), .Y(n31842) );
  AOI21X1 U19100 ( .A(n31847), .B(n31848), .C(n25493), .Y(rd1data1033_8_) );
  NOR2X1 U19101 ( .A(n31849), .B(n31850), .Y(n31848) );
  NAND3X1 U19102 ( .A(n31851), .B(n31852), .C(n31853), .Y(n31850) );
  NOR2X1 U19103 ( .A(n31854), .B(n31855), .Y(n31853) );
  OAI22X1 U19104 ( .A(n26599), .B(n25504), .C(n26600), .D(n25514), .Y(n31855)
         );
  OAI22X1 U19105 ( .A(n26601), .B(n25525), .C(n26602), .D(n25535), .Y(n31854)
         );
  AOI22X1 U19106 ( .A(n25546), .B(reg_file[1416]), .C(n25557), .D(
        reg_file[1288]), .Y(n31852) );
  AOI22X1 U19107 ( .A(n25568), .B(reg_file[1160]), .C(n25579), .D(
        reg_file[1032]), .Y(n31851) );
  NAND3X1 U19108 ( .A(n31856), .B(n31857), .C(n31858), .Y(n31849) );
  NOR2X1 U19109 ( .A(n31859), .B(n31860), .Y(n31858) );
  OAI22X1 U19110 ( .A(n26608), .B(n25590), .C(n26609), .D(n25600), .Y(n31860)
         );
  OAI22X1 U19111 ( .A(n26610), .B(n25611), .C(n26611), .D(n25621), .Y(n31859)
         );
  AOI22X1 U19112 ( .A(n25632), .B(reg_file[520]), .C(n25643), .D(reg_file[648]), .Y(n31857) );
  AOI22X1 U19113 ( .A(n25654), .B(reg_file[776]), .C(n25665), .D(reg_file[904]), .Y(n31856) );
  NOR2X1 U19114 ( .A(n31861), .B(n31862), .Y(n31847) );
  NAND3X1 U19115 ( .A(n31863), .B(n31864), .C(n31865), .Y(n31862) );
  NOR2X1 U19116 ( .A(n31866), .B(n31867), .Y(n31865) );
  OAI22X1 U19117 ( .A(n26619), .B(n25676), .C(n26620), .D(n25686), .Y(n31867)
         );
  OAI22X1 U19118 ( .A(n26621), .B(n25697), .C(n26622), .D(n25707), .Y(n31866)
         );
  AOI22X1 U19119 ( .A(n25718), .B(reg_file[3464]), .C(n25729), .D(
        reg_file[3336]), .Y(n31864) );
  AOI22X1 U19120 ( .A(n25740), .B(reg_file[3208]), .C(n25751), .D(
        reg_file[3080]), .Y(n31863) );
  NAND3X1 U19121 ( .A(n31868), .B(n31869), .C(n31870), .Y(n31861) );
  NOR2X1 U19122 ( .A(n31871), .B(n31872), .Y(n31870) );
  OAI22X1 U19123 ( .A(n26628), .B(n25762), .C(n26629), .D(n25772), .Y(n31872)
         );
  OAI22X1 U19124 ( .A(n26630), .B(n25783), .C(n26631), .D(n25793), .Y(n31871)
         );
  AOI22X1 U19125 ( .A(n25804), .B(reg_file[2440]), .C(n25815), .D(
        reg_file[2312]), .Y(n31869) );
  AOI22X1 U19126 ( .A(n25826), .B(reg_file[2184]), .C(n25837), .D(
        reg_file[2056]), .Y(n31868) );
  AOI21X1 U19127 ( .A(n31873), .B(n31874), .C(n25493), .Y(rd1data1033_89_) );
  NOR2X1 U19128 ( .A(n31875), .B(n31876), .Y(n31874) );
  NAND3X1 U19129 ( .A(n31877), .B(n31878), .C(n31879), .Y(n31876) );
  NOR2X1 U19130 ( .A(n31880), .B(n31881), .Y(n31879) );
  OAI22X1 U19131 ( .A(n26641), .B(n25504), .C(n26642), .D(n25514), .Y(n31881)
         );
  OAI22X1 U19132 ( .A(n26643), .B(n25525), .C(n26644), .D(n25535), .Y(n31880)
         );
  AOI22X1 U19133 ( .A(n25546), .B(reg_file[1497]), .C(n25557), .D(
        reg_file[1369]), .Y(n31878) );
  AOI22X1 U19134 ( .A(n25568), .B(reg_file[1241]), .C(n25579), .D(
        reg_file[1113]), .Y(n31877) );
  NAND3X1 U19135 ( .A(n31882), .B(n31883), .C(n31884), .Y(n31875) );
  NOR2X1 U19136 ( .A(n31885), .B(n31886), .Y(n31884) );
  OAI22X1 U19137 ( .A(n26650), .B(n25590), .C(n26651), .D(n25600), .Y(n31886)
         );
  OAI22X1 U19138 ( .A(n26652), .B(n25611), .C(n26653), .D(n25621), .Y(n31885)
         );
  AOI22X1 U19139 ( .A(n25632), .B(reg_file[601]), .C(n25643), .D(reg_file[729]), .Y(n31883) );
  AOI22X1 U19140 ( .A(n25654), .B(reg_file[857]), .C(n25665), .D(reg_file[985]), .Y(n31882) );
  NOR2X1 U19141 ( .A(n31887), .B(n31888), .Y(n31873) );
  NAND3X1 U19142 ( .A(n31889), .B(n31890), .C(n31891), .Y(n31888) );
  NOR2X1 U19143 ( .A(n31892), .B(n31893), .Y(n31891) );
  OAI22X1 U19144 ( .A(n26661), .B(n25676), .C(n26662), .D(n25686), .Y(n31893)
         );
  OAI22X1 U19145 ( .A(n26663), .B(n25697), .C(n26664), .D(n25707), .Y(n31892)
         );
  AOI22X1 U19146 ( .A(n25718), .B(reg_file[3545]), .C(n25729), .D(
        reg_file[3417]), .Y(n31890) );
  AOI22X1 U19147 ( .A(n25740), .B(reg_file[3289]), .C(n25751), .D(
        reg_file[3161]), .Y(n31889) );
  NAND3X1 U19148 ( .A(n31894), .B(n31895), .C(n31896), .Y(n31887) );
  NOR2X1 U19149 ( .A(n31897), .B(n31898), .Y(n31896) );
  OAI22X1 U19150 ( .A(n26670), .B(n25762), .C(n26671), .D(n25772), .Y(n31898)
         );
  OAI22X1 U19151 ( .A(n26672), .B(n25783), .C(n26673), .D(n25793), .Y(n31897)
         );
  AOI22X1 U19152 ( .A(n25804), .B(reg_file[2521]), .C(n25815), .D(
        reg_file[2393]), .Y(n31895) );
  AOI22X1 U19153 ( .A(n25826), .B(reg_file[2265]), .C(n25837), .D(
        reg_file[2137]), .Y(n31894) );
  AOI21X1 U19154 ( .A(n31899), .B(n31900), .C(n25493), .Y(rd1data1033_88_) );
  NOR2X1 U19155 ( .A(n31901), .B(n31902), .Y(n31900) );
  NAND3X1 U19156 ( .A(n31903), .B(n31904), .C(n31905), .Y(n31902) );
  NOR2X1 U19157 ( .A(n31906), .B(n31907), .Y(n31905) );
  OAI22X1 U19158 ( .A(n26683), .B(n25504), .C(n26684), .D(n25514), .Y(n31907)
         );
  OAI22X1 U19159 ( .A(n26685), .B(n25525), .C(n26686), .D(n25535), .Y(n31906)
         );
  AOI22X1 U19160 ( .A(n25546), .B(reg_file[1496]), .C(n25557), .D(
        reg_file[1368]), .Y(n31904) );
  AOI22X1 U19161 ( .A(n25568), .B(reg_file[1240]), .C(n25579), .D(
        reg_file[1112]), .Y(n31903) );
  NAND3X1 U19162 ( .A(n31908), .B(n31909), .C(n31910), .Y(n31901) );
  NOR2X1 U19163 ( .A(n31911), .B(n31912), .Y(n31910) );
  OAI22X1 U19164 ( .A(n26692), .B(n25590), .C(n26693), .D(n25600), .Y(n31912)
         );
  OAI22X1 U19165 ( .A(n26694), .B(n25611), .C(n26695), .D(n25621), .Y(n31911)
         );
  AOI22X1 U19166 ( .A(n25632), .B(reg_file[600]), .C(n25643), .D(reg_file[728]), .Y(n31909) );
  AOI22X1 U19167 ( .A(n25654), .B(reg_file[856]), .C(n25665), .D(reg_file[984]), .Y(n31908) );
  NOR2X1 U19168 ( .A(n31913), .B(n31914), .Y(n31899) );
  NAND3X1 U19169 ( .A(n31915), .B(n31916), .C(n31917), .Y(n31914) );
  NOR2X1 U19170 ( .A(n31918), .B(n31919), .Y(n31917) );
  OAI22X1 U19171 ( .A(n26703), .B(n25676), .C(n26704), .D(n25686), .Y(n31919)
         );
  OAI22X1 U19172 ( .A(n26705), .B(n25697), .C(n26706), .D(n25707), .Y(n31918)
         );
  AOI22X1 U19173 ( .A(n25718), .B(reg_file[3544]), .C(n25729), .D(
        reg_file[3416]), .Y(n31916) );
  AOI22X1 U19174 ( .A(n25740), .B(reg_file[3288]), .C(n25751), .D(
        reg_file[3160]), .Y(n31915) );
  NAND3X1 U19175 ( .A(n31920), .B(n31921), .C(n31922), .Y(n31913) );
  NOR2X1 U19176 ( .A(n31923), .B(n31924), .Y(n31922) );
  OAI22X1 U19177 ( .A(n26712), .B(n25762), .C(n26713), .D(n25772), .Y(n31924)
         );
  OAI22X1 U19178 ( .A(n26714), .B(n25783), .C(n26715), .D(n25793), .Y(n31923)
         );
  AOI22X1 U19179 ( .A(n25804), .B(reg_file[2520]), .C(n25815), .D(
        reg_file[2392]), .Y(n31921) );
  AOI22X1 U19180 ( .A(n25826), .B(reg_file[2264]), .C(n25837), .D(
        reg_file[2136]), .Y(n31920) );
  AOI21X1 U19181 ( .A(n31925), .B(n31926), .C(n25493), .Y(rd1data1033_87_) );
  NOR2X1 U19182 ( .A(n31927), .B(n31928), .Y(n31926) );
  NAND3X1 U19183 ( .A(n31929), .B(n31930), .C(n31931), .Y(n31928) );
  NOR2X1 U19184 ( .A(n31932), .B(n31933), .Y(n31931) );
  OAI22X1 U19185 ( .A(n26725), .B(n25504), .C(n26726), .D(n25514), .Y(n31933)
         );
  OAI22X1 U19186 ( .A(n26727), .B(n25525), .C(n26728), .D(n25535), .Y(n31932)
         );
  AOI22X1 U19187 ( .A(n25546), .B(reg_file[1495]), .C(n25557), .D(
        reg_file[1367]), .Y(n31930) );
  AOI22X1 U19188 ( .A(n25568), .B(reg_file[1239]), .C(n25579), .D(
        reg_file[1111]), .Y(n31929) );
  NAND3X1 U19189 ( .A(n31934), .B(n31935), .C(n31936), .Y(n31927) );
  NOR2X1 U19190 ( .A(n31937), .B(n31938), .Y(n31936) );
  OAI22X1 U19191 ( .A(n26734), .B(n25590), .C(n26735), .D(n25600), .Y(n31938)
         );
  OAI22X1 U19192 ( .A(n26736), .B(n25611), .C(n26737), .D(n25621), .Y(n31937)
         );
  AOI22X1 U19193 ( .A(n25632), .B(reg_file[599]), .C(n25643), .D(reg_file[727]), .Y(n31935) );
  AOI22X1 U19194 ( .A(n25654), .B(reg_file[855]), .C(n25665), .D(reg_file[983]), .Y(n31934) );
  NOR2X1 U19195 ( .A(n31939), .B(n31940), .Y(n31925) );
  NAND3X1 U19196 ( .A(n31941), .B(n31942), .C(n31943), .Y(n31940) );
  NOR2X1 U19197 ( .A(n31944), .B(n31945), .Y(n31943) );
  OAI22X1 U19198 ( .A(n26745), .B(n25676), .C(n26746), .D(n25686), .Y(n31945)
         );
  OAI22X1 U19199 ( .A(n26747), .B(n25697), .C(n26748), .D(n25707), .Y(n31944)
         );
  AOI22X1 U19200 ( .A(n25718), .B(reg_file[3543]), .C(n25729), .D(
        reg_file[3415]), .Y(n31942) );
  AOI22X1 U19201 ( .A(n25740), .B(reg_file[3287]), .C(n25751), .D(
        reg_file[3159]), .Y(n31941) );
  NAND3X1 U19202 ( .A(n31946), .B(n31947), .C(n31948), .Y(n31939) );
  NOR2X1 U19203 ( .A(n31949), .B(n31950), .Y(n31948) );
  OAI22X1 U19204 ( .A(n26754), .B(n25762), .C(n26755), .D(n25772), .Y(n31950)
         );
  OAI22X1 U19205 ( .A(n26756), .B(n25783), .C(n26757), .D(n25793), .Y(n31949)
         );
  AOI22X1 U19206 ( .A(n25804), .B(reg_file[2519]), .C(n25815), .D(
        reg_file[2391]), .Y(n31947) );
  AOI22X1 U19207 ( .A(n25826), .B(reg_file[2263]), .C(n25837), .D(
        reg_file[2135]), .Y(n31946) );
  AOI21X1 U19208 ( .A(n31951), .B(n31952), .C(n25493), .Y(rd1data1033_86_) );
  NOR2X1 U19209 ( .A(n31953), .B(n31954), .Y(n31952) );
  NAND3X1 U19210 ( .A(n31955), .B(n31956), .C(n31957), .Y(n31954) );
  NOR2X1 U19211 ( .A(n31958), .B(n31959), .Y(n31957) );
  OAI22X1 U19212 ( .A(n26767), .B(n25504), .C(n26768), .D(n25514), .Y(n31959)
         );
  OAI22X1 U19213 ( .A(n26769), .B(n25525), .C(n26770), .D(n25535), .Y(n31958)
         );
  AOI22X1 U19214 ( .A(n25546), .B(reg_file[1494]), .C(n25557), .D(
        reg_file[1366]), .Y(n31956) );
  AOI22X1 U19215 ( .A(n25568), .B(reg_file[1238]), .C(n25579), .D(
        reg_file[1110]), .Y(n31955) );
  NAND3X1 U19216 ( .A(n31960), .B(n31961), .C(n31962), .Y(n31953) );
  NOR2X1 U19217 ( .A(n31963), .B(n31964), .Y(n31962) );
  OAI22X1 U19218 ( .A(n26776), .B(n25590), .C(n26777), .D(n25600), .Y(n31964)
         );
  OAI22X1 U19219 ( .A(n26778), .B(n25611), .C(n26779), .D(n25621), .Y(n31963)
         );
  AOI22X1 U19220 ( .A(n25632), .B(reg_file[598]), .C(n25643), .D(reg_file[726]), .Y(n31961) );
  AOI22X1 U19221 ( .A(n25654), .B(reg_file[854]), .C(n25665), .D(reg_file[982]), .Y(n31960) );
  NOR2X1 U19222 ( .A(n31965), .B(n31966), .Y(n31951) );
  NAND3X1 U19223 ( .A(n31967), .B(n31968), .C(n31969), .Y(n31966) );
  NOR2X1 U19224 ( .A(n31970), .B(n31971), .Y(n31969) );
  OAI22X1 U19225 ( .A(n26787), .B(n25676), .C(n26788), .D(n25686), .Y(n31971)
         );
  OAI22X1 U19226 ( .A(n26789), .B(n25697), .C(n26790), .D(n25707), .Y(n31970)
         );
  AOI22X1 U19227 ( .A(n25718), .B(reg_file[3542]), .C(n25729), .D(
        reg_file[3414]), .Y(n31968) );
  AOI22X1 U19228 ( .A(n25740), .B(reg_file[3286]), .C(n25751), .D(
        reg_file[3158]), .Y(n31967) );
  NAND3X1 U19229 ( .A(n31972), .B(n31973), .C(n31974), .Y(n31965) );
  NOR2X1 U19230 ( .A(n31975), .B(n31976), .Y(n31974) );
  OAI22X1 U19231 ( .A(n26796), .B(n25762), .C(n26797), .D(n25772), .Y(n31976)
         );
  OAI22X1 U19232 ( .A(n26798), .B(n25783), .C(n26799), .D(n25793), .Y(n31975)
         );
  AOI22X1 U19233 ( .A(n25804), .B(reg_file[2518]), .C(n25815), .D(
        reg_file[2390]), .Y(n31973) );
  AOI22X1 U19234 ( .A(n25826), .B(reg_file[2262]), .C(n25837), .D(
        reg_file[2134]), .Y(n31972) );
  AOI21X1 U19235 ( .A(n31977), .B(n31978), .C(n25493), .Y(rd1data1033_85_) );
  NOR2X1 U19236 ( .A(n31979), .B(n31980), .Y(n31978) );
  NAND3X1 U19237 ( .A(n31981), .B(n31982), .C(n31983), .Y(n31980) );
  NOR2X1 U19238 ( .A(n31984), .B(n31985), .Y(n31983) );
  OAI22X1 U19239 ( .A(n26809), .B(n25504), .C(n26810), .D(n25514), .Y(n31985)
         );
  OAI22X1 U19240 ( .A(n26811), .B(n25525), .C(n26812), .D(n25535), .Y(n31984)
         );
  AOI22X1 U19241 ( .A(n25546), .B(reg_file[1493]), .C(n25557), .D(
        reg_file[1365]), .Y(n31982) );
  AOI22X1 U19242 ( .A(n25568), .B(reg_file[1237]), .C(n25579), .D(
        reg_file[1109]), .Y(n31981) );
  NAND3X1 U19243 ( .A(n31986), .B(n31987), .C(n31988), .Y(n31979) );
  NOR2X1 U19244 ( .A(n31989), .B(n31990), .Y(n31988) );
  OAI22X1 U19245 ( .A(n26818), .B(n25590), .C(n26819), .D(n25600), .Y(n31990)
         );
  OAI22X1 U19246 ( .A(n26820), .B(n25611), .C(n26821), .D(n25621), .Y(n31989)
         );
  AOI22X1 U19247 ( .A(n25632), .B(reg_file[597]), .C(n25643), .D(reg_file[725]), .Y(n31987) );
  AOI22X1 U19248 ( .A(n25654), .B(reg_file[853]), .C(n25665), .D(reg_file[981]), .Y(n31986) );
  NOR2X1 U19249 ( .A(n31991), .B(n31992), .Y(n31977) );
  NAND3X1 U19250 ( .A(n31993), .B(n31994), .C(n31995), .Y(n31992) );
  NOR2X1 U19251 ( .A(n31996), .B(n31997), .Y(n31995) );
  OAI22X1 U19252 ( .A(n26829), .B(n25676), .C(n26830), .D(n25686), .Y(n31997)
         );
  OAI22X1 U19253 ( .A(n26831), .B(n25697), .C(n26832), .D(n25707), .Y(n31996)
         );
  AOI22X1 U19254 ( .A(n25718), .B(reg_file[3541]), .C(n25729), .D(
        reg_file[3413]), .Y(n31994) );
  AOI22X1 U19255 ( .A(n25740), .B(reg_file[3285]), .C(n25751), .D(
        reg_file[3157]), .Y(n31993) );
  NAND3X1 U19256 ( .A(n31998), .B(n31999), .C(n32000), .Y(n31991) );
  NOR2X1 U19257 ( .A(n32001), .B(n32002), .Y(n32000) );
  OAI22X1 U19258 ( .A(n26838), .B(n25762), .C(n26839), .D(n25772), .Y(n32002)
         );
  OAI22X1 U19259 ( .A(n26840), .B(n25783), .C(n26841), .D(n25793), .Y(n32001)
         );
  AOI22X1 U19260 ( .A(n25804), .B(reg_file[2517]), .C(n25815), .D(
        reg_file[2389]), .Y(n31999) );
  AOI22X1 U19261 ( .A(n25826), .B(reg_file[2261]), .C(n25837), .D(
        reg_file[2133]), .Y(n31998) );
  AOI21X1 U19262 ( .A(n32003), .B(n32004), .C(n25493), .Y(rd1data1033_84_) );
  NOR2X1 U19263 ( .A(n32005), .B(n32006), .Y(n32004) );
  NAND3X1 U19264 ( .A(n32007), .B(n32008), .C(n32009), .Y(n32006) );
  NOR2X1 U19265 ( .A(n32010), .B(n32011), .Y(n32009) );
  OAI22X1 U19266 ( .A(n26851), .B(n25504), .C(n26852), .D(n25514), .Y(n32011)
         );
  OAI22X1 U19267 ( .A(n26853), .B(n25525), .C(n26854), .D(n25535), .Y(n32010)
         );
  AOI22X1 U19268 ( .A(n25546), .B(reg_file[1492]), .C(n25557), .D(
        reg_file[1364]), .Y(n32008) );
  AOI22X1 U19269 ( .A(n25568), .B(reg_file[1236]), .C(n25579), .D(
        reg_file[1108]), .Y(n32007) );
  NAND3X1 U19270 ( .A(n32012), .B(n32013), .C(n32014), .Y(n32005) );
  NOR2X1 U19271 ( .A(n32015), .B(n32016), .Y(n32014) );
  OAI22X1 U19272 ( .A(n26860), .B(n25590), .C(n26861), .D(n25600), .Y(n32016)
         );
  OAI22X1 U19273 ( .A(n26862), .B(n25611), .C(n26863), .D(n25621), .Y(n32015)
         );
  AOI22X1 U19274 ( .A(n25632), .B(reg_file[596]), .C(n25643), .D(reg_file[724]), .Y(n32013) );
  AOI22X1 U19275 ( .A(n25654), .B(reg_file[852]), .C(n25665), .D(reg_file[980]), .Y(n32012) );
  NOR2X1 U19276 ( .A(n32017), .B(n32018), .Y(n32003) );
  NAND3X1 U19277 ( .A(n32019), .B(n32020), .C(n32021), .Y(n32018) );
  NOR2X1 U19278 ( .A(n32022), .B(n32023), .Y(n32021) );
  OAI22X1 U19279 ( .A(n26871), .B(n25676), .C(n26872), .D(n25686), .Y(n32023)
         );
  OAI22X1 U19280 ( .A(n26873), .B(n25697), .C(n26874), .D(n25707), .Y(n32022)
         );
  AOI22X1 U19281 ( .A(n25718), .B(reg_file[3540]), .C(n25729), .D(
        reg_file[3412]), .Y(n32020) );
  AOI22X1 U19282 ( .A(n25740), .B(reg_file[3284]), .C(n25751), .D(
        reg_file[3156]), .Y(n32019) );
  NAND3X1 U19283 ( .A(n32024), .B(n32025), .C(n32026), .Y(n32017) );
  NOR2X1 U19284 ( .A(n32027), .B(n32028), .Y(n32026) );
  OAI22X1 U19285 ( .A(n26880), .B(n25762), .C(n26881), .D(n25772), .Y(n32028)
         );
  OAI22X1 U19286 ( .A(n26882), .B(n25783), .C(n26883), .D(n25793), .Y(n32027)
         );
  AOI22X1 U19287 ( .A(n25804), .B(reg_file[2516]), .C(n25815), .D(
        reg_file[2388]), .Y(n32025) );
  AOI22X1 U19288 ( .A(n25826), .B(reg_file[2260]), .C(n25837), .D(
        reg_file[2132]), .Y(n32024) );
  AOI21X1 U19289 ( .A(n32029), .B(n32030), .C(n25493), .Y(rd1data1033_83_) );
  NOR2X1 U19290 ( .A(n32031), .B(n32032), .Y(n32030) );
  NAND3X1 U19291 ( .A(n32033), .B(n32034), .C(n32035), .Y(n32032) );
  NOR2X1 U19292 ( .A(n32036), .B(n32037), .Y(n32035) );
  OAI22X1 U19293 ( .A(n26893), .B(n25504), .C(n26894), .D(n25514), .Y(n32037)
         );
  OAI22X1 U19294 ( .A(n26895), .B(n25525), .C(n26896), .D(n25535), .Y(n32036)
         );
  AOI22X1 U19295 ( .A(n25546), .B(reg_file[1491]), .C(n25557), .D(
        reg_file[1363]), .Y(n32034) );
  AOI22X1 U19296 ( .A(n25568), .B(reg_file[1235]), .C(n25579), .D(
        reg_file[1107]), .Y(n32033) );
  NAND3X1 U19297 ( .A(n32038), .B(n32039), .C(n32040), .Y(n32031) );
  NOR2X1 U19298 ( .A(n32041), .B(n32042), .Y(n32040) );
  OAI22X1 U19299 ( .A(n26902), .B(n25590), .C(n26903), .D(n25600), .Y(n32042)
         );
  OAI22X1 U19300 ( .A(n26904), .B(n25611), .C(n26905), .D(n25621), .Y(n32041)
         );
  AOI22X1 U19301 ( .A(n25632), .B(reg_file[595]), .C(n25643), .D(reg_file[723]), .Y(n32039) );
  AOI22X1 U19302 ( .A(n25654), .B(reg_file[851]), .C(n25665), .D(reg_file[979]), .Y(n32038) );
  NOR2X1 U19303 ( .A(n32043), .B(n32044), .Y(n32029) );
  NAND3X1 U19304 ( .A(n32045), .B(n32046), .C(n32047), .Y(n32044) );
  NOR2X1 U19305 ( .A(n32048), .B(n32049), .Y(n32047) );
  OAI22X1 U19306 ( .A(n26913), .B(n25676), .C(n26914), .D(n25686), .Y(n32049)
         );
  OAI22X1 U19307 ( .A(n26915), .B(n25697), .C(n26916), .D(n25707), .Y(n32048)
         );
  AOI22X1 U19308 ( .A(n25718), .B(reg_file[3539]), .C(n25729), .D(
        reg_file[3411]), .Y(n32046) );
  AOI22X1 U19309 ( .A(n25740), .B(reg_file[3283]), .C(n25751), .D(
        reg_file[3155]), .Y(n32045) );
  NAND3X1 U19310 ( .A(n32050), .B(n32051), .C(n32052), .Y(n32043) );
  NOR2X1 U19311 ( .A(n32053), .B(n32054), .Y(n32052) );
  OAI22X1 U19312 ( .A(n26922), .B(n25762), .C(n26923), .D(n25772), .Y(n32054)
         );
  OAI22X1 U19313 ( .A(n26924), .B(n25783), .C(n26925), .D(n25793), .Y(n32053)
         );
  AOI22X1 U19314 ( .A(n25804), .B(reg_file[2515]), .C(n25815), .D(
        reg_file[2387]), .Y(n32051) );
  AOI22X1 U19315 ( .A(n25826), .B(reg_file[2259]), .C(n25837), .D(
        reg_file[2131]), .Y(n32050) );
  AOI21X1 U19316 ( .A(n32055), .B(n32056), .C(n25493), .Y(rd1data1033_82_) );
  NOR2X1 U19317 ( .A(n32057), .B(n32058), .Y(n32056) );
  NAND3X1 U19318 ( .A(n32059), .B(n32060), .C(n32061), .Y(n32058) );
  NOR2X1 U19319 ( .A(n32062), .B(n32063), .Y(n32061) );
  OAI22X1 U19320 ( .A(n26935), .B(n25504), .C(n26936), .D(n25514), .Y(n32063)
         );
  OAI22X1 U19321 ( .A(n26937), .B(n25525), .C(n26938), .D(n25535), .Y(n32062)
         );
  AOI22X1 U19322 ( .A(n25546), .B(reg_file[1490]), .C(n25557), .D(
        reg_file[1362]), .Y(n32060) );
  AOI22X1 U19323 ( .A(n25568), .B(reg_file[1234]), .C(n25579), .D(
        reg_file[1106]), .Y(n32059) );
  NAND3X1 U19324 ( .A(n32064), .B(n32065), .C(n32066), .Y(n32057) );
  NOR2X1 U19325 ( .A(n32067), .B(n32068), .Y(n32066) );
  OAI22X1 U19326 ( .A(n26944), .B(n25590), .C(n26945), .D(n25600), .Y(n32068)
         );
  OAI22X1 U19327 ( .A(n26946), .B(n25611), .C(n26947), .D(n25621), .Y(n32067)
         );
  AOI22X1 U19328 ( .A(n25632), .B(reg_file[594]), .C(n25643), .D(reg_file[722]), .Y(n32065) );
  AOI22X1 U19329 ( .A(n25654), .B(reg_file[850]), .C(n25665), .D(reg_file[978]), .Y(n32064) );
  NOR2X1 U19330 ( .A(n32069), .B(n32070), .Y(n32055) );
  NAND3X1 U19331 ( .A(n32071), .B(n32072), .C(n32073), .Y(n32070) );
  NOR2X1 U19332 ( .A(n32074), .B(n32075), .Y(n32073) );
  OAI22X1 U19333 ( .A(n26955), .B(n25676), .C(n26956), .D(n25686), .Y(n32075)
         );
  OAI22X1 U19334 ( .A(n26957), .B(n25697), .C(n26958), .D(n25707), .Y(n32074)
         );
  AOI22X1 U19335 ( .A(n25718), .B(reg_file[3538]), .C(n25729), .D(
        reg_file[3410]), .Y(n32072) );
  AOI22X1 U19336 ( .A(n25740), .B(reg_file[3282]), .C(n25751), .D(
        reg_file[3154]), .Y(n32071) );
  NAND3X1 U19337 ( .A(n32076), .B(n32077), .C(n32078), .Y(n32069) );
  NOR2X1 U19338 ( .A(n32079), .B(n32080), .Y(n32078) );
  OAI22X1 U19339 ( .A(n26964), .B(n25762), .C(n26965), .D(n25772), .Y(n32080)
         );
  OAI22X1 U19340 ( .A(n26966), .B(n25783), .C(n26967), .D(n25793), .Y(n32079)
         );
  AOI22X1 U19341 ( .A(n25804), .B(reg_file[2514]), .C(n25815), .D(
        reg_file[2386]), .Y(n32077) );
  AOI22X1 U19342 ( .A(n25826), .B(reg_file[2258]), .C(n25837), .D(
        reg_file[2130]), .Y(n32076) );
  AOI21X1 U19343 ( .A(n32081), .B(n32082), .C(n25492), .Y(rd1data1033_81_) );
  NOR2X1 U19344 ( .A(n32083), .B(n32084), .Y(n32082) );
  NAND3X1 U19345 ( .A(n32085), .B(n32086), .C(n32087), .Y(n32084) );
  NOR2X1 U19346 ( .A(n32088), .B(n32089), .Y(n32087) );
  OAI22X1 U19347 ( .A(n26977), .B(n25503), .C(n26978), .D(n25514), .Y(n32089)
         );
  OAI22X1 U19348 ( .A(n26979), .B(n25524), .C(n26980), .D(n25535), .Y(n32088)
         );
  AOI22X1 U19349 ( .A(n25545), .B(reg_file[1489]), .C(n25556), .D(
        reg_file[1361]), .Y(n32086) );
  AOI22X1 U19350 ( .A(n25567), .B(reg_file[1233]), .C(n25578), .D(
        reg_file[1105]), .Y(n32085) );
  NAND3X1 U19351 ( .A(n32090), .B(n32091), .C(n32092), .Y(n32083) );
  NOR2X1 U19352 ( .A(n32093), .B(n32094), .Y(n32092) );
  OAI22X1 U19353 ( .A(n26986), .B(n25589), .C(n26987), .D(n25600), .Y(n32094)
         );
  OAI22X1 U19354 ( .A(n26988), .B(n25610), .C(n26989), .D(n25621), .Y(n32093)
         );
  AOI22X1 U19355 ( .A(n25631), .B(reg_file[593]), .C(n25642), .D(reg_file[721]), .Y(n32091) );
  AOI22X1 U19356 ( .A(n25653), .B(reg_file[849]), .C(n25664), .D(reg_file[977]), .Y(n32090) );
  NOR2X1 U19357 ( .A(n32095), .B(n32096), .Y(n32081) );
  NAND3X1 U19358 ( .A(n32097), .B(n32098), .C(n32099), .Y(n32096) );
  NOR2X1 U19359 ( .A(n32100), .B(n32101), .Y(n32099) );
  OAI22X1 U19360 ( .A(n26997), .B(n25675), .C(n26998), .D(n25686), .Y(n32101)
         );
  OAI22X1 U19361 ( .A(n26999), .B(n25696), .C(n27000), .D(n25707), .Y(n32100)
         );
  AOI22X1 U19362 ( .A(n25717), .B(reg_file[3537]), .C(n25728), .D(
        reg_file[3409]), .Y(n32098) );
  AOI22X1 U19363 ( .A(n25739), .B(reg_file[3281]), .C(n25750), .D(
        reg_file[3153]), .Y(n32097) );
  NAND3X1 U19364 ( .A(n32102), .B(n32103), .C(n32104), .Y(n32095) );
  NOR2X1 U19365 ( .A(n32105), .B(n32106), .Y(n32104) );
  OAI22X1 U19366 ( .A(n27006), .B(n25761), .C(n27007), .D(n25772), .Y(n32106)
         );
  OAI22X1 U19367 ( .A(n27008), .B(n25782), .C(n27009), .D(n25793), .Y(n32105)
         );
  AOI22X1 U19368 ( .A(n25803), .B(reg_file[2513]), .C(n25814), .D(
        reg_file[2385]), .Y(n32103) );
  AOI22X1 U19369 ( .A(n25825), .B(reg_file[2257]), .C(n25836), .D(
        reg_file[2129]), .Y(n32102) );
  AOI21X1 U19370 ( .A(n32107), .B(n32108), .C(n25492), .Y(rd1data1033_80_) );
  NOR2X1 U19371 ( .A(n32109), .B(n32110), .Y(n32108) );
  NAND3X1 U19372 ( .A(n32111), .B(n32112), .C(n32113), .Y(n32110) );
  NOR2X1 U19373 ( .A(n32114), .B(n32115), .Y(n32113) );
  OAI22X1 U19374 ( .A(n27019), .B(n25503), .C(n27020), .D(n25514), .Y(n32115)
         );
  OAI22X1 U19375 ( .A(n27021), .B(n25524), .C(n27022), .D(n25535), .Y(n32114)
         );
  AOI22X1 U19376 ( .A(n25545), .B(reg_file[1488]), .C(n25556), .D(
        reg_file[1360]), .Y(n32112) );
  AOI22X1 U19377 ( .A(n25567), .B(reg_file[1232]), .C(n25578), .D(
        reg_file[1104]), .Y(n32111) );
  NAND3X1 U19378 ( .A(n32116), .B(n32117), .C(n32118), .Y(n32109) );
  NOR2X1 U19379 ( .A(n32119), .B(n32120), .Y(n32118) );
  OAI22X1 U19380 ( .A(n27028), .B(n25589), .C(n27029), .D(n25600), .Y(n32120)
         );
  OAI22X1 U19381 ( .A(n27030), .B(n25610), .C(n27031), .D(n25621), .Y(n32119)
         );
  AOI22X1 U19382 ( .A(n25631), .B(reg_file[592]), .C(n25642), .D(reg_file[720]), .Y(n32117) );
  AOI22X1 U19383 ( .A(n25653), .B(reg_file[848]), .C(n25664), .D(reg_file[976]), .Y(n32116) );
  NOR2X1 U19384 ( .A(n32121), .B(n32122), .Y(n32107) );
  NAND3X1 U19385 ( .A(n32123), .B(n32124), .C(n32125), .Y(n32122) );
  NOR2X1 U19386 ( .A(n32126), .B(n32127), .Y(n32125) );
  OAI22X1 U19387 ( .A(n27039), .B(n25675), .C(n27040), .D(n25686), .Y(n32127)
         );
  OAI22X1 U19388 ( .A(n27041), .B(n25696), .C(n27042), .D(n25707), .Y(n32126)
         );
  AOI22X1 U19389 ( .A(n25717), .B(reg_file[3536]), .C(n25728), .D(
        reg_file[3408]), .Y(n32124) );
  AOI22X1 U19390 ( .A(n25739), .B(reg_file[3280]), .C(n25750), .D(
        reg_file[3152]), .Y(n32123) );
  NAND3X1 U19391 ( .A(n32128), .B(n32129), .C(n32130), .Y(n32121) );
  NOR2X1 U19392 ( .A(n32131), .B(n32132), .Y(n32130) );
  OAI22X1 U19393 ( .A(n27048), .B(n25761), .C(n27049), .D(n25772), .Y(n32132)
         );
  OAI22X1 U19394 ( .A(n27050), .B(n25782), .C(n27051), .D(n25793), .Y(n32131)
         );
  AOI22X1 U19395 ( .A(n25803), .B(reg_file[2512]), .C(n25814), .D(
        reg_file[2384]), .Y(n32129) );
  AOI22X1 U19396 ( .A(n25825), .B(reg_file[2256]), .C(n25836), .D(
        reg_file[2128]), .Y(n32128) );
  AOI21X1 U19397 ( .A(n32133), .B(n32134), .C(n25492), .Y(rd1data1033_7_) );
  NOR2X1 U19398 ( .A(n32135), .B(n32136), .Y(n32134) );
  NAND3X1 U19399 ( .A(n32137), .B(n32138), .C(n32139), .Y(n32136) );
  NOR2X1 U19400 ( .A(n32140), .B(n32141), .Y(n32139) );
  OAI22X1 U19401 ( .A(n27061), .B(n25503), .C(n27062), .D(n25514), .Y(n32141)
         );
  OAI22X1 U19402 ( .A(n27063), .B(n25524), .C(n27064), .D(n25535), .Y(n32140)
         );
  AOI22X1 U19403 ( .A(n25545), .B(reg_file[1415]), .C(n25556), .D(
        reg_file[1287]), .Y(n32138) );
  AOI22X1 U19404 ( .A(n25567), .B(reg_file[1159]), .C(n25578), .D(
        reg_file[1031]), .Y(n32137) );
  NAND3X1 U19405 ( .A(n32142), .B(n32143), .C(n32144), .Y(n32135) );
  NOR2X1 U19406 ( .A(n32145), .B(n32146), .Y(n32144) );
  OAI22X1 U19407 ( .A(n27070), .B(n25589), .C(n27071), .D(n25600), .Y(n32146)
         );
  OAI22X1 U19408 ( .A(n27072), .B(n25610), .C(n27073), .D(n25621), .Y(n32145)
         );
  AOI22X1 U19409 ( .A(n25631), .B(reg_file[519]), .C(n25642), .D(reg_file[647]), .Y(n32143) );
  AOI22X1 U19410 ( .A(n25653), .B(reg_file[775]), .C(n25664), .D(reg_file[903]), .Y(n32142) );
  NOR2X1 U19411 ( .A(n32147), .B(n32148), .Y(n32133) );
  NAND3X1 U19412 ( .A(n32149), .B(n32150), .C(n32151), .Y(n32148) );
  NOR2X1 U19413 ( .A(n32152), .B(n32153), .Y(n32151) );
  OAI22X1 U19414 ( .A(n27081), .B(n25675), .C(n27082), .D(n25686), .Y(n32153)
         );
  OAI22X1 U19415 ( .A(n27083), .B(n25696), .C(n27084), .D(n25707), .Y(n32152)
         );
  AOI22X1 U19416 ( .A(n25717), .B(reg_file[3463]), .C(n25728), .D(
        reg_file[3335]), .Y(n32150) );
  AOI22X1 U19417 ( .A(n25739), .B(reg_file[3207]), .C(n25750), .D(
        reg_file[3079]), .Y(n32149) );
  NAND3X1 U19418 ( .A(n32154), .B(n32155), .C(n32156), .Y(n32147) );
  NOR2X1 U19419 ( .A(n32157), .B(n32158), .Y(n32156) );
  OAI22X1 U19420 ( .A(n27090), .B(n25761), .C(n27091), .D(n25772), .Y(n32158)
         );
  OAI22X1 U19421 ( .A(n27092), .B(n25782), .C(n27093), .D(n25793), .Y(n32157)
         );
  AOI22X1 U19422 ( .A(n25803), .B(reg_file[2439]), .C(n25814), .D(
        reg_file[2311]), .Y(n32155) );
  AOI22X1 U19423 ( .A(n25825), .B(reg_file[2183]), .C(n25836), .D(
        reg_file[2055]), .Y(n32154) );
  AOI21X1 U19424 ( .A(n32159), .B(n32160), .C(n25492), .Y(rd1data1033_79_) );
  NOR2X1 U19425 ( .A(n32161), .B(n32162), .Y(n32160) );
  NAND3X1 U19426 ( .A(n32163), .B(n32164), .C(n32165), .Y(n32162) );
  NOR2X1 U19427 ( .A(n32166), .B(n32167), .Y(n32165) );
  OAI22X1 U19428 ( .A(n27103), .B(n25503), .C(n27104), .D(n25514), .Y(n32167)
         );
  OAI22X1 U19429 ( .A(n27105), .B(n25524), .C(n27106), .D(n25535), .Y(n32166)
         );
  AOI22X1 U19430 ( .A(n25545), .B(reg_file[1487]), .C(n25556), .D(
        reg_file[1359]), .Y(n32164) );
  AOI22X1 U19431 ( .A(n25567), .B(reg_file[1231]), .C(n25578), .D(
        reg_file[1103]), .Y(n32163) );
  NAND3X1 U19432 ( .A(n32168), .B(n32169), .C(n32170), .Y(n32161) );
  NOR2X1 U19433 ( .A(n32171), .B(n32172), .Y(n32170) );
  OAI22X1 U19434 ( .A(n27112), .B(n25589), .C(n27113), .D(n25600), .Y(n32172)
         );
  OAI22X1 U19435 ( .A(n27114), .B(n25610), .C(n27115), .D(n25621), .Y(n32171)
         );
  AOI22X1 U19436 ( .A(n25631), .B(reg_file[591]), .C(n25642), .D(reg_file[719]), .Y(n32169) );
  AOI22X1 U19437 ( .A(n25653), .B(reg_file[847]), .C(n25664), .D(reg_file[975]), .Y(n32168) );
  NOR2X1 U19438 ( .A(n32173), .B(n32174), .Y(n32159) );
  NAND3X1 U19439 ( .A(n32175), .B(n32176), .C(n32177), .Y(n32174) );
  NOR2X1 U19440 ( .A(n32178), .B(n32179), .Y(n32177) );
  OAI22X1 U19441 ( .A(n27123), .B(n25675), .C(n27124), .D(n25686), .Y(n32179)
         );
  OAI22X1 U19442 ( .A(n27125), .B(n25696), .C(n27126), .D(n25707), .Y(n32178)
         );
  AOI22X1 U19443 ( .A(n25717), .B(reg_file[3535]), .C(n25728), .D(
        reg_file[3407]), .Y(n32176) );
  AOI22X1 U19444 ( .A(n25739), .B(reg_file[3279]), .C(n25750), .D(
        reg_file[3151]), .Y(n32175) );
  NAND3X1 U19445 ( .A(n32180), .B(n32181), .C(n32182), .Y(n32173) );
  NOR2X1 U19446 ( .A(n32183), .B(n32184), .Y(n32182) );
  OAI22X1 U19447 ( .A(n27132), .B(n25761), .C(n27133), .D(n25772), .Y(n32184)
         );
  OAI22X1 U19448 ( .A(n27134), .B(n25782), .C(n27135), .D(n25793), .Y(n32183)
         );
  AOI22X1 U19449 ( .A(n25803), .B(reg_file[2511]), .C(n25814), .D(
        reg_file[2383]), .Y(n32181) );
  AOI22X1 U19450 ( .A(n25825), .B(reg_file[2255]), .C(n25836), .D(
        reg_file[2127]), .Y(n32180) );
  AOI21X1 U19451 ( .A(n32185), .B(n32186), .C(n25492), .Y(rd1data1033_78_) );
  NOR2X1 U19452 ( .A(n32187), .B(n32188), .Y(n32186) );
  NAND3X1 U19453 ( .A(n32189), .B(n32190), .C(n32191), .Y(n32188) );
  NOR2X1 U19454 ( .A(n32192), .B(n32193), .Y(n32191) );
  OAI22X1 U19455 ( .A(n27145), .B(n25503), .C(n27146), .D(n25513), .Y(n32193)
         );
  OAI22X1 U19456 ( .A(n27147), .B(n25524), .C(n27148), .D(n25534), .Y(n32192)
         );
  AOI22X1 U19457 ( .A(n25545), .B(reg_file[1486]), .C(n25556), .D(
        reg_file[1358]), .Y(n32190) );
  AOI22X1 U19458 ( .A(n25567), .B(reg_file[1230]), .C(n25578), .D(
        reg_file[1102]), .Y(n32189) );
  NAND3X1 U19459 ( .A(n32194), .B(n32195), .C(n32196), .Y(n32187) );
  NOR2X1 U19460 ( .A(n32197), .B(n32198), .Y(n32196) );
  OAI22X1 U19461 ( .A(n27154), .B(n25589), .C(n27155), .D(n25599), .Y(n32198)
         );
  OAI22X1 U19462 ( .A(n27156), .B(n25610), .C(n27157), .D(n25620), .Y(n32197)
         );
  AOI22X1 U19463 ( .A(n25631), .B(reg_file[590]), .C(n25642), .D(reg_file[718]), .Y(n32195) );
  AOI22X1 U19464 ( .A(n25653), .B(reg_file[846]), .C(n25664), .D(reg_file[974]), .Y(n32194) );
  NOR2X1 U19465 ( .A(n32199), .B(n32200), .Y(n32185) );
  NAND3X1 U19466 ( .A(n32201), .B(n32202), .C(n32203), .Y(n32200) );
  NOR2X1 U19467 ( .A(n32204), .B(n32205), .Y(n32203) );
  OAI22X1 U19468 ( .A(n27165), .B(n25675), .C(n27166), .D(n25685), .Y(n32205)
         );
  OAI22X1 U19469 ( .A(n27167), .B(n25696), .C(n27168), .D(n25706), .Y(n32204)
         );
  AOI22X1 U19470 ( .A(n25717), .B(reg_file[3534]), .C(n25728), .D(
        reg_file[3406]), .Y(n32202) );
  AOI22X1 U19471 ( .A(n25739), .B(reg_file[3278]), .C(n25750), .D(
        reg_file[3150]), .Y(n32201) );
  NAND3X1 U19472 ( .A(n32206), .B(n32207), .C(n32208), .Y(n32199) );
  NOR2X1 U19473 ( .A(n32209), .B(n32210), .Y(n32208) );
  OAI22X1 U19474 ( .A(n27174), .B(n25761), .C(n27175), .D(n25771), .Y(n32210)
         );
  OAI22X1 U19475 ( .A(n27176), .B(n25782), .C(n27177), .D(n25792), .Y(n32209)
         );
  AOI22X1 U19476 ( .A(n25803), .B(reg_file[2510]), .C(n25814), .D(
        reg_file[2382]), .Y(n32207) );
  AOI22X1 U19477 ( .A(n25825), .B(reg_file[2254]), .C(n25836), .D(
        reg_file[2126]), .Y(n32206) );
  AOI21X1 U19478 ( .A(n32211), .B(n32212), .C(n25492), .Y(rd1data1033_77_) );
  NOR2X1 U19479 ( .A(n32213), .B(n32214), .Y(n32212) );
  NAND3X1 U19480 ( .A(n32215), .B(n32216), .C(n32217), .Y(n32214) );
  NOR2X1 U19481 ( .A(n32218), .B(n32219), .Y(n32217) );
  OAI22X1 U19482 ( .A(n27187), .B(n25503), .C(n27188), .D(n25513), .Y(n32219)
         );
  OAI22X1 U19483 ( .A(n27189), .B(n25524), .C(n27190), .D(n25534), .Y(n32218)
         );
  AOI22X1 U19484 ( .A(n25545), .B(reg_file[1485]), .C(n25556), .D(
        reg_file[1357]), .Y(n32216) );
  AOI22X1 U19485 ( .A(n25567), .B(reg_file[1229]), .C(n25578), .D(
        reg_file[1101]), .Y(n32215) );
  NAND3X1 U19486 ( .A(n32220), .B(n32221), .C(n32222), .Y(n32213) );
  NOR2X1 U19487 ( .A(n32223), .B(n32224), .Y(n32222) );
  OAI22X1 U19488 ( .A(n27196), .B(n25589), .C(n27197), .D(n25599), .Y(n32224)
         );
  OAI22X1 U19489 ( .A(n27198), .B(n25610), .C(n27199), .D(n25620), .Y(n32223)
         );
  AOI22X1 U19490 ( .A(n25631), .B(reg_file[589]), .C(n25642), .D(reg_file[717]), .Y(n32221) );
  AOI22X1 U19491 ( .A(n25653), .B(reg_file[845]), .C(n25664), .D(reg_file[973]), .Y(n32220) );
  NOR2X1 U19492 ( .A(n32225), .B(n32226), .Y(n32211) );
  NAND3X1 U19493 ( .A(n32227), .B(n32228), .C(n32229), .Y(n32226) );
  NOR2X1 U19494 ( .A(n32230), .B(n32231), .Y(n32229) );
  OAI22X1 U19495 ( .A(n27207), .B(n25675), .C(n27208), .D(n25685), .Y(n32231)
         );
  OAI22X1 U19496 ( .A(n27209), .B(n25696), .C(n27210), .D(n25706), .Y(n32230)
         );
  AOI22X1 U19497 ( .A(n25717), .B(reg_file[3533]), .C(n25728), .D(
        reg_file[3405]), .Y(n32228) );
  AOI22X1 U19498 ( .A(n25739), .B(reg_file[3277]), .C(n25750), .D(
        reg_file[3149]), .Y(n32227) );
  NAND3X1 U19499 ( .A(n32232), .B(n32233), .C(n32234), .Y(n32225) );
  NOR2X1 U19500 ( .A(n32235), .B(n32236), .Y(n32234) );
  OAI22X1 U19501 ( .A(n27216), .B(n25761), .C(n27217), .D(n25771), .Y(n32236)
         );
  OAI22X1 U19502 ( .A(n27218), .B(n25782), .C(n27219), .D(n25792), .Y(n32235)
         );
  AOI22X1 U19503 ( .A(n25803), .B(reg_file[2509]), .C(n25814), .D(
        reg_file[2381]), .Y(n32233) );
  AOI22X1 U19504 ( .A(n25825), .B(reg_file[2253]), .C(n25836), .D(
        reg_file[2125]), .Y(n32232) );
  AOI21X1 U19505 ( .A(n32237), .B(n32238), .C(n25492), .Y(rd1data1033_76_) );
  NOR2X1 U19506 ( .A(n32239), .B(n32240), .Y(n32238) );
  NAND3X1 U19507 ( .A(n32241), .B(n32242), .C(n32243), .Y(n32240) );
  NOR2X1 U19508 ( .A(n32244), .B(n32245), .Y(n32243) );
  OAI22X1 U19509 ( .A(n27229), .B(n25503), .C(n27230), .D(n25513), .Y(n32245)
         );
  OAI22X1 U19510 ( .A(n27231), .B(n25524), .C(n27232), .D(n25534), .Y(n32244)
         );
  AOI22X1 U19511 ( .A(n25545), .B(reg_file[1484]), .C(n25556), .D(
        reg_file[1356]), .Y(n32242) );
  AOI22X1 U19512 ( .A(n25567), .B(reg_file[1228]), .C(n25578), .D(
        reg_file[1100]), .Y(n32241) );
  NAND3X1 U19513 ( .A(n32246), .B(n32247), .C(n32248), .Y(n32239) );
  NOR2X1 U19514 ( .A(n32249), .B(n32250), .Y(n32248) );
  OAI22X1 U19515 ( .A(n27238), .B(n25589), .C(n27239), .D(n25599), .Y(n32250)
         );
  OAI22X1 U19516 ( .A(n27240), .B(n25610), .C(n27241), .D(n25620), .Y(n32249)
         );
  AOI22X1 U19517 ( .A(n25631), .B(reg_file[588]), .C(n25642), .D(reg_file[716]), .Y(n32247) );
  AOI22X1 U19518 ( .A(n25653), .B(reg_file[844]), .C(n25664), .D(reg_file[972]), .Y(n32246) );
  NOR2X1 U19519 ( .A(n32251), .B(n32252), .Y(n32237) );
  NAND3X1 U19520 ( .A(n32253), .B(n32254), .C(n32255), .Y(n32252) );
  NOR2X1 U19521 ( .A(n32256), .B(n32257), .Y(n32255) );
  OAI22X1 U19522 ( .A(n27249), .B(n25675), .C(n27250), .D(n25685), .Y(n32257)
         );
  OAI22X1 U19523 ( .A(n27251), .B(n25696), .C(n27252), .D(n25706), .Y(n32256)
         );
  AOI22X1 U19524 ( .A(n25717), .B(reg_file[3532]), .C(n25728), .D(
        reg_file[3404]), .Y(n32254) );
  AOI22X1 U19525 ( .A(n25739), .B(reg_file[3276]), .C(n25750), .D(
        reg_file[3148]), .Y(n32253) );
  NAND3X1 U19526 ( .A(n32258), .B(n32259), .C(n32260), .Y(n32251) );
  NOR2X1 U19527 ( .A(n32261), .B(n32262), .Y(n32260) );
  OAI22X1 U19528 ( .A(n27258), .B(n25761), .C(n27259), .D(n25771), .Y(n32262)
         );
  OAI22X1 U19529 ( .A(n27260), .B(n25782), .C(n27261), .D(n25792), .Y(n32261)
         );
  AOI22X1 U19530 ( .A(n25803), .B(reg_file[2508]), .C(n25814), .D(
        reg_file[2380]), .Y(n32259) );
  AOI22X1 U19531 ( .A(n25825), .B(reg_file[2252]), .C(n25836), .D(
        reg_file[2124]), .Y(n32258) );
  AOI21X1 U19532 ( .A(n32263), .B(n32264), .C(n25492), .Y(rd1data1033_75_) );
  NOR2X1 U19533 ( .A(n32265), .B(n32266), .Y(n32264) );
  NAND3X1 U19534 ( .A(n32267), .B(n32268), .C(n32269), .Y(n32266) );
  NOR2X1 U19535 ( .A(n32270), .B(n32271), .Y(n32269) );
  OAI22X1 U19536 ( .A(n27271), .B(n25503), .C(n27272), .D(n25513), .Y(n32271)
         );
  OAI22X1 U19537 ( .A(n27273), .B(n25524), .C(n27274), .D(n25534), .Y(n32270)
         );
  AOI22X1 U19538 ( .A(n25545), .B(reg_file[1483]), .C(n25556), .D(
        reg_file[1355]), .Y(n32268) );
  AOI22X1 U19539 ( .A(n25567), .B(reg_file[1227]), .C(n25578), .D(
        reg_file[1099]), .Y(n32267) );
  NAND3X1 U19540 ( .A(n32272), .B(n32273), .C(n32274), .Y(n32265) );
  NOR2X1 U19541 ( .A(n32275), .B(n32276), .Y(n32274) );
  OAI22X1 U19542 ( .A(n27280), .B(n25589), .C(n27281), .D(n25599), .Y(n32276)
         );
  OAI22X1 U19543 ( .A(n27282), .B(n25610), .C(n27283), .D(n25620), .Y(n32275)
         );
  AOI22X1 U19544 ( .A(n25631), .B(reg_file[587]), .C(n25642), .D(reg_file[715]), .Y(n32273) );
  AOI22X1 U19545 ( .A(n25653), .B(reg_file[843]), .C(n25664), .D(reg_file[971]), .Y(n32272) );
  NOR2X1 U19546 ( .A(n32277), .B(n32278), .Y(n32263) );
  NAND3X1 U19547 ( .A(n32279), .B(n32280), .C(n32281), .Y(n32278) );
  NOR2X1 U19548 ( .A(n32282), .B(n32283), .Y(n32281) );
  OAI22X1 U19549 ( .A(n27291), .B(n25675), .C(n27292), .D(n25685), .Y(n32283)
         );
  OAI22X1 U19550 ( .A(n27293), .B(n25696), .C(n27294), .D(n25706), .Y(n32282)
         );
  AOI22X1 U19551 ( .A(n25717), .B(reg_file[3531]), .C(n25728), .D(
        reg_file[3403]), .Y(n32280) );
  AOI22X1 U19552 ( .A(n25739), .B(reg_file[3275]), .C(n25750), .D(
        reg_file[3147]), .Y(n32279) );
  NAND3X1 U19553 ( .A(n32284), .B(n32285), .C(n32286), .Y(n32277) );
  NOR2X1 U19554 ( .A(n32287), .B(n32288), .Y(n32286) );
  OAI22X1 U19555 ( .A(n27300), .B(n25761), .C(n27301), .D(n25771), .Y(n32288)
         );
  OAI22X1 U19556 ( .A(n27302), .B(n25782), .C(n27303), .D(n25792), .Y(n32287)
         );
  AOI22X1 U19557 ( .A(n25803), .B(reg_file[2507]), .C(n25814), .D(
        reg_file[2379]), .Y(n32285) );
  AOI22X1 U19558 ( .A(n25825), .B(reg_file[2251]), .C(n25836), .D(
        reg_file[2123]), .Y(n32284) );
  AOI21X1 U19559 ( .A(n32289), .B(n32290), .C(n25492), .Y(rd1data1033_74_) );
  NOR2X1 U19560 ( .A(n32291), .B(n32292), .Y(n32290) );
  NAND3X1 U19561 ( .A(n32293), .B(n32294), .C(n32295), .Y(n32292) );
  NOR2X1 U19562 ( .A(n32296), .B(n32297), .Y(n32295) );
  OAI22X1 U19563 ( .A(n27313), .B(n25503), .C(n27314), .D(n25513), .Y(n32297)
         );
  OAI22X1 U19564 ( .A(n27315), .B(n25524), .C(n27316), .D(n25534), .Y(n32296)
         );
  AOI22X1 U19565 ( .A(n25545), .B(reg_file[1482]), .C(n25556), .D(
        reg_file[1354]), .Y(n32294) );
  AOI22X1 U19566 ( .A(n25567), .B(reg_file[1226]), .C(n25578), .D(
        reg_file[1098]), .Y(n32293) );
  NAND3X1 U19567 ( .A(n32298), .B(n32299), .C(n32300), .Y(n32291) );
  NOR2X1 U19568 ( .A(n32301), .B(n32302), .Y(n32300) );
  OAI22X1 U19569 ( .A(n27322), .B(n25589), .C(n27323), .D(n25599), .Y(n32302)
         );
  OAI22X1 U19570 ( .A(n27324), .B(n25610), .C(n27325), .D(n25620), .Y(n32301)
         );
  AOI22X1 U19571 ( .A(n25631), .B(reg_file[586]), .C(n25642), .D(reg_file[714]), .Y(n32299) );
  AOI22X1 U19572 ( .A(n25653), .B(reg_file[842]), .C(n25664), .D(reg_file[970]), .Y(n32298) );
  NOR2X1 U19573 ( .A(n32303), .B(n32304), .Y(n32289) );
  NAND3X1 U19574 ( .A(n32305), .B(n32306), .C(n32307), .Y(n32304) );
  NOR2X1 U19575 ( .A(n32308), .B(n32309), .Y(n32307) );
  OAI22X1 U19576 ( .A(n27333), .B(n25675), .C(n27334), .D(n25685), .Y(n32309)
         );
  OAI22X1 U19577 ( .A(n27335), .B(n25696), .C(n27336), .D(n25706), .Y(n32308)
         );
  AOI22X1 U19578 ( .A(n25717), .B(reg_file[3530]), .C(n25728), .D(
        reg_file[3402]), .Y(n32306) );
  AOI22X1 U19579 ( .A(n25739), .B(reg_file[3274]), .C(n25750), .D(
        reg_file[3146]), .Y(n32305) );
  NAND3X1 U19580 ( .A(n32310), .B(n32311), .C(n32312), .Y(n32303) );
  NOR2X1 U19581 ( .A(n32313), .B(n32314), .Y(n32312) );
  OAI22X1 U19582 ( .A(n27342), .B(n25761), .C(n27343), .D(n25771), .Y(n32314)
         );
  OAI22X1 U19583 ( .A(n27344), .B(n25782), .C(n27345), .D(n25792), .Y(n32313)
         );
  AOI22X1 U19584 ( .A(n25803), .B(reg_file[2506]), .C(n25814), .D(
        reg_file[2378]), .Y(n32311) );
  AOI22X1 U19585 ( .A(n25825), .B(reg_file[2250]), .C(n25836), .D(
        reg_file[2122]), .Y(n32310) );
  AOI21X1 U19586 ( .A(n32315), .B(n32316), .C(n25492), .Y(rd1data1033_73_) );
  NOR2X1 U19587 ( .A(n32317), .B(n32318), .Y(n32316) );
  NAND3X1 U19588 ( .A(n32319), .B(n32320), .C(n32321), .Y(n32318) );
  NOR2X1 U19589 ( .A(n32322), .B(n32323), .Y(n32321) );
  OAI22X1 U19590 ( .A(n27355), .B(n25503), .C(n27356), .D(n25513), .Y(n32323)
         );
  OAI22X1 U19591 ( .A(n27357), .B(n25524), .C(n27358), .D(n25534), .Y(n32322)
         );
  AOI22X1 U19592 ( .A(n25545), .B(reg_file[1481]), .C(n25556), .D(
        reg_file[1353]), .Y(n32320) );
  AOI22X1 U19593 ( .A(n25567), .B(reg_file[1225]), .C(n25578), .D(
        reg_file[1097]), .Y(n32319) );
  NAND3X1 U19594 ( .A(n32324), .B(n32325), .C(n32326), .Y(n32317) );
  NOR2X1 U19595 ( .A(n32327), .B(n32328), .Y(n32326) );
  OAI22X1 U19596 ( .A(n27364), .B(n25589), .C(n27365), .D(n25599), .Y(n32328)
         );
  OAI22X1 U19597 ( .A(n27366), .B(n25610), .C(n27367), .D(n25620), .Y(n32327)
         );
  AOI22X1 U19598 ( .A(n25631), .B(reg_file[585]), .C(n25642), .D(reg_file[713]), .Y(n32325) );
  AOI22X1 U19599 ( .A(n25653), .B(reg_file[841]), .C(n25664), .D(reg_file[969]), .Y(n32324) );
  NOR2X1 U19600 ( .A(n32329), .B(n32330), .Y(n32315) );
  NAND3X1 U19601 ( .A(n32331), .B(n32332), .C(n32333), .Y(n32330) );
  NOR2X1 U19602 ( .A(n32334), .B(n32335), .Y(n32333) );
  OAI22X1 U19603 ( .A(n27375), .B(n25675), .C(n27376), .D(n25685), .Y(n32335)
         );
  OAI22X1 U19604 ( .A(n27377), .B(n25696), .C(n27378), .D(n25706), .Y(n32334)
         );
  AOI22X1 U19605 ( .A(n25717), .B(reg_file[3529]), .C(n25728), .D(
        reg_file[3401]), .Y(n32332) );
  AOI22X1 U19606 ( .A(n25739), .B(reg_file[3273]), .C(n25750), .D(
        reg_file[3145]), .Y(n32331) );
  NAND3X1 U19607 ( .A(n32336), .B(n32337), .C(n32338), .Y(n32329) );
  NOR2X1 U19608 ( .A(n32339), .B(n32340), .Y(n32338) );
  OAI22X1 U19609 ( .A(n27384), .B(n25761), .C(n27385), .D(n25771), .Y(n32340)
         );
  OAI22X1 U19610 ( .A(n27386), .B(n25782), .C(n27387), .D(n25792), .Y(n32339)
         );
  AOI22X1 U19611 ( .A(n25803), .B(reg_file[2505]), .C(n25814), .D(
        reg_file[2377]), .Y(n32337) );
  AOI22X1 U19612 ( .A(n25825), .B(reg_file[2249]), .C(n25836), .D(
        reg_file[2121]), .Y(n32336) );
  AOI21X1 U19613 ( .A(n32341), .B(n32342), .C(n25492), .Y(rd1data1033_72_) );
  NOR2X1 U19614 ( .A(n32343), .B(n32344), .Y(n32342) );
  NAND3X1 U19615 ( .A(n32345), .B(n32346), .C(n32347), .Y(n32344) );
  NOR2X1 U19616 ( .A(n32348), .B(n32349), .Y(n32347) );
  OAI22X1 U19617 ( .A(n27397), .B(n25503), .C(n27398), .D(n25513), .Y(n32349)
         );
  OAI22X1 U19618 ( .A(n27399), .B(n25524), .C(n27400), .D(n25534), .Y(n32348)
         );
  AOI22X1 U19619 ( .A(n25545), .B(reg_file[1480]), .C(n25556), .D(
        reg_file[1352]), .Y(n32346) );
  AOI22X1 U19620 ( .A(n25567), .B(reg_file[1224]), .C(n25578), .D(
        reg_file[1096]), .Y(n32345) );
  NAND3X1 U19621 ( .A(n32350), .B(n32351), .C(n32352), .Y(n32343) );
  NOR2X1 U19622 ( .A(n32353), .B(n32354), .Y(n32352) );
  OAI22X1 U19623 ( .A(n27406), .B(n25589), .C(n27407), .D(n25599), .Y(n32354)
         );
  OAI22X1 U19624 ( .A(n27408), .B(n25610), .C(n27409), .D(n25620), .Y(n32353)
         );
  AOI22X1 U19625 ( .A(n25631), .B(reg_file[584]), .C(n25642), .D(reg_file[712]), .Y(n32351) );
  AOI22X1 U19626 ( .A(n25653), .B(reg_file[840]), .C(n25664), .D(reg_file[968]), .Y(n32350) );
  NOR2X1 U19627 ( .A(n32355), .B(n32356), .Y(n32341) );
  NAND3X1 U19628 ( .A(n32357), .B(n32358), .C(n32359), .Y(n32356) );
  NOR2X1 U19629 ( .A(n32360), .B(n32361), .Y(n32359) );
  OAI22X1 U19630 ( .A(n27417), .B(n25675), .C(n27418), .D(n25685), .Y(n32361)
         );
  OAI22X1 U19631 ( .A(n27419), .B(n25696), .C(n27420), .D(n25706), .Y(n32360)
         );
  AOI22X1 U19632 ( .A(n25717), .B(reg_file[3528]), .C(n25728), .D(
        reg_file[3400]), .Y(n32358) );
  AOI22X1 U19633 ( .A(n25739), .B(reg_file[3272]), .C(n25750), .D(
        reg_file[3144]), .Y(n32357) );
  NAND3X1 U19634 ( .A(n32362), .B(n32363), .C(n32364), .Y(n32355) );
  NOR2X1 U19635 ( .A(n32365), .B(n32366), .Y(n32364) );
  OAI22X1 U19636 ( .A(n27426), .B(n25761), .C(n27427), .D(n25771), .Y(n32366)
         );
  OAI22X1 U19637 ( .A(n27428), .B(n25782), .C(n27429), .D(n25792), .Y(n32365)
         );
  AOI22X1 U19638 ( .A(n25803), .B(reg_file[2504]), .C(n25814), .D(
        reg_file[2376]), .Y(n32363) );
  AOI22X1 U19639 ( .A(n25825), .B(reg_file[2248]), .C(n25836), .D(
        reg_file[2120]), .Y(n32362) );
  AOI21X1 U19640 ( .A(n32367), .B(n32368), .C(n25492), .Y(rd1data1033_71_) );
  NOR2X1 U19641 ( .A(n32369), .B(n32370), .Y(n32368) );
  NAND3X1 U19642 ( .A(n32371), .B(n32372), .C(n32373), .Y(n32370) );
  NOR2X1 U19643 ( .A(n32374), .B(n32375), .Y(n32373) );
  OAI22X1 U19644 ( .A(n27439), .B(n25503), .C(n27440), .D(n25513), .Y(n32375)
         );
  OAI22X1 U19645 ( .A(n27441), .B(n25524), .C(n27442), .D(n25534), .Y(n32374)
         );
  AOI22X1 U19646 ( .A(n25545), .B(reg_file[1479]), .C(n25556), .D(
        reg_file[1351]), .Y(n32372) );
  AOI22X1 U19647 ( .A(n25567), .B(reg_file[1223]), .C(n25578), .D(
        reg_file[1095]), .Y(n32371) );
  NAND3X1 U19648 ( .A(n32376), .B(n32377), .C(n32378), .Y(n32369) );
  NOR2X1 U19649 ( .A(n32379), .B(n32380), .Y(n32378) );
  OAI22X1 U19650 ( .A(n27448), .B(n25589), .C(n27449), .D(n25599), .Y(n32380)
         );
  OAI22X1 U19651 ( .A(n27450), .B(n25610), .C(n27451), .D(n25620), .Y(n32379)
         );
  AOI22X1 U19652 ( .A(n25631), .B(reg_file[583]), .C(n25642), .D(reg_file[711]), .Y(n32377) );
  AOI22X1 U19653 ( .A(n25653), .B(reg_file[839]), .C(n25664), .D(reg_file[967]), .Y(n32376) );
  NOR2X1 U19654 ( .A(n32381), .B(n32382), .Y(n32367) );
  NAND3X1 U19655 ( .A(n32383), .B(n32384), .C(n32385), .Y(n32382) );
  NOR2X1 U19656 ( .A(n32386), .B(n32387), .Y(n32385) );
  OAI22X1 U19657 ( .A(n27459), .B(n25675), .C(n27460), .D(n25685), .Y(n32387)
         );
  OAI22X1 U19658 ( .A(n27461), .B(n25696), .C(n27462), .D(n25706), .Y(n32386)
         );
  AOI22X1 U19659 ( .A(n25717), .B(reg_file[3527]), .C(n25728), .D(
        reg_file[3399]), .Y(n32384) );
  AOI22X1 U19660 ( .A(n25739), .B(reg_file[3271]), .C(n25750), .D(
        reg_file[3143]), .Y(n32383) );
  NAND3X1 U19661 ( .A(n32388), .B(n32389), .C(n32390), .Y(n32381) );
  NOR2X1 U19662 ( .A(n32391), .B(n32392), .Y(n32390) );
  OAI22X1 U19663 ( .A(n27468), .B(n25761), .C(n27469), .D(n25771), .Y(n32392)
         );
  OAI22X1 U19664 ( .A(n27470), .B(n25782), .C(n27471), .D(n25792), .Y(n32391)
         );
  AOI22X1 U19665 ( .A(n25803), .B(reg_file[2503]), .C(n25814), .D(
        reg_file[2375]), .Y(n32389) );
  AOI22X1 U19666 ( .A(n25825), .B(reg_file[2247]), .C(n25836), .D(
        reg_file[2119]), .Y(n32388) );
  AOI21X1 U19667 ( .A(n32393), .B(n32394), .C(n25491), .Y(rd1data1033_70_) );
  NOR2X1 U19668 ( .A(n32395), .B(n32396), .Y(n32394) );
  NAND3X1 U19669 ( .A(n32397), .B(n32398), .C(n32399), .Y(n32396) );
  NOR2X1 U19670 ( .A(n32400), .B(n32401), .Y(n32399) );
  OAI22X1 U19671 ( .A(n27481), .B(n25502), .C(n27482), .D(n25513), .Y(n32401)
         );
  OAI22X1 U19672 ( .A(n27483), .B(n25523), .C(n27484), .D(n25534), .Y(n32400)
         );
  AOI22X1 U19673 ( .A(n25544), .B(reg_file[1478]), .C(n25555), .D(
        reg_file[1350]), .Y(n32398) );
  AOI22X1 U19674 ( .A(n25566), .B(reg_file[1222]), .C(n25577), .D(
        reg_file[1094]), .Y(n32397) );
  NAND3X1 U19675 ( .A(n32402), .B(n32403), .C(n32404), .Y(n32395) );
  NOR2X1 U19676 ( .A(n32405), .B(n32406), .Y(n32404) );
  OAI22X1 U19677 ( .A(n27490), .B(n25588), .C(n27491), .D(n25599), .Y(n32406)
         );
  OAI22X1 U19678 ( .A(n27492), .B(n25609), .C(n27493), .D(n25620), .Y(n32405)
         );
  AOI22X1 U19679 ( .A(n25630), .B(reg_file[582]), .C(n25641), .D(reg_file[710]), .Y(n32403) );
  AOI22X1 U19680 ( .A(n25652), .B(reg_file[838]), .C(n25663), .D(reg_file[966]), .Y(n32402) );
  NOR2X1 U19681 ( .A(n32407), .B(n32408), .Y(n32393) );
  NAND3X1 U19682 ( .A(n32409), .B(n32410), .C(n32411), .Y(n32408) );
  NOR2X1 U19683 ( .A(n32412), .B(n32413), .Y(n32411) );
  OAI22X1 U19684 ( .A(n27501), .B(n25674), .C(n27502), .D(n25685), .Y(n32413)
         );
  OAI22X1 U19685 ( .A(n27503), .B(n25695), .C(n27504), .D(n25706), .Y(n32412)
         );
  AOI22X1 U19686 ( .A(n25716), .B(reg_file[3526]), .C(n25727), .D(
        reg_file[3398]), .Y(n32410) );
  AOI22X1 U19687 ( .A(n25738), .B(reg_file[3270]), .C(n25749), .D(
        reg_file[3142]), .Y(n32409) );
  NAND3X1 U19688 ( .A(n32414), .B(n32415), .C(n32416), .Y(n32407) );
  NOR2X1 U19689 ( .A(n32417), .B(n32418), .Y(n32416) );
  OAI22X1 U19690 ( .A(n27510), .B(n25760), .C(n27511), .D(n25771), .Y(n32418)
         );
  OAI22X1 U19691 ( .A(n27512), .B(n25781), .C(n27513), .D(n25792), .Y(n32417)
         );
  AOI22X1 U19692 ( .A(n25802), .B(reg_file[2502]), .C(n25813), .D(
        reg_file[2374]), .Y(n32415) );
  AOI22X1 U19693 ( .A(n25824), .B(reg_file[2246]), .C(n25835), .D(
        reg_file[2118]), .Y(n32414) );
  AOI21X1 U19694 ( .A(n32419), .B(n32420), .C(n25491), .Y(rd1data1033_6_) );
  NOR2X1 U19695 ( .A(n32421), .B(n32422), .Y(n32420) );
  NAND3X1 U19696 ( .A(n32423), .B(n32424), .C(n32425), .Y(n32422) );
  NOR2X1 U19697 ( .A(n32426), .B(n32427), .Y(n32425) );
  OAI22X1 U19698 ( .A(n27523), .B(n25502), .C(n27524), .D(n25513), .Y(n32427)
         );
  OAI22X1 U19699 ( .A(n27525), .B(n25523), .C(n27526), .D(n25534), .Y(n32426)
         );
  AOI22X1 U19700 ( .A(n25544), .B(reg_file[1414]), .C(n25555), .D(
        reg_file[1286]), .Y(n32424) );
  AOI22X1 U19701 ( .A(n25566), .B(reg_file[1158]), .C(n25577), .D(
        reg_file[1030]), .Y(n32423) );
  NAND3X1 U19702 ( .A(n32428), .B(n32429), .C(n32430), .Y(n32421) );
  NOR2X1 U19703 ( .A(n32431), .B(n32432), .Y(n32430) );
  OAI22X1 U19704 ( .A(n27532), .B(n25588), .C(n27533), .D(n25599), .Y(n32432)
         );
  OAI22X1 U19705 ( .A(n27534), .B(n25609), .C(n27535), .D(n25620), .Y(n32431)
         );
  AOI22X1 U19706 ( .A(n25630), .B(reg_file[518]), .C(n25641), .D(reg_file[646]), .Y(n32429) );
  AOI22X1 U19707 ( .A(n25652), .B(reg_file[774]), .C(n25663), .D(reg_file[902]), .Y(n32428) );
  NOR2X1 U19708 ( .A(n32433), .B(n32434), .Y(n32419) );
  NAND3X1 U19709 ( .A(n32435), .B(n32436), .C(n32437), .Y(n32434) );
  NOR2X1 U19710 ( .A(n32438), .B(n32439), .Y(n32437) );
  OAI22X1 U19711 ( .A(n27543), .B(n25674), .C(n27544), .D(n25685), .Y(n32439)
         );
  OAI22X1 U19712 ( .A(n27545), .B(n25695), .C(n27546), .D(n25706), .Y(n32438)
         );
  AOI22X1 U19713 ( .A(n25716), .B(reg_file[3462]), .C(n25727), .D(
        reg_file[3334]), .Y(n32436) );
  AOI22X1 U19714 ( .A(n25738), .B(reg_file[3206]), .C(n25749), .D(
        reg_file[3078]), .Y(n32435) );
  NAND3X1 U19715 ( .A(n32440), .B(n32441), .C(n32442), .Y(n32433) );
  NOR2X1 U19716 ( .A(n32443), .B(n32444), .Y(n32442) );
  OAI22X1 U19717 ( .A(n27552), .B(n25760), .C(n27553), .D(n25771), .Y(n32444)
         );
  OAI22X1 U19718 ( .A(n27554), .B(n25781), .C(n27555), .D(n25792), .Y(n32443)
         );
  AOI22X1 U19719 ( .A(n25802), .B(reg_file[2438]), .C(n25813), .D(
        reg_file[2310]), .Y(n32441) );
  AOI22X1 U19720 ( .A(n25824), .B(reg_file[2182]), .C(n25835), .D(
        reg_file[2054]), .Y(n32440) );
  AOI21X1 U19721 ( .A(n32445), .B(n32446), .C(n25491), .Y(rd1data1033_69_) );
  NOR2X1 U19722 ( .A(n32447), .B(n32448), .Y(n32446) );
  NAND3X1 U19723 ( .A(n32449), .B(n32450), .C(n32451), .Y(n32448) );
  NOR2X1 U19724 ( .A(n32452), .B(n32453), .Y(n32451) );
  OAI22X1 U19725 ( .A(n27565), .B(n25502), .C(n27566), .D(n25513), .Y(n32453)
         );
  OAI22X1 U19726 ( .A(n27567), .B(n25523), .C(n27568), .D(n25534), .Y(n32452)
         );
  AOI22X1 U19727 ( .A(n25544), .B(reg_file[1477]), .C(n25555), .D(
        reg_file[1349]), .Y(n32450) );
  AOI22X1 U19728 ( .A(n25566), .B(reg_file[1221]), .C(n25577), .D(
        reg_file[1093]), .Y(n32449) );
  NAND3X1 U19729 ( .A(n32454), .B(n32455), .C(n32456), .Y(n32447) );
  NOR2X1 U19730 ( .A(n32457), .B(n32458), .Y(n32456) );
  OAI22X1 U19731 ( .A(n27574), .B(n25588), .C(n27575), .D(n25599), .Y(n32458)
         );
  OAI22X1 U19732 ( .A(n27576), .B(n25609), .C(n27577), .D(n25620), .Y(n32457)
         );
  AOI22X1 U19733 ( .A(n25630), .B(reg_file[581]), .C(n25641), .D(reg_file[709]), .Y(n32455) );
  AOI22X1 U19734 ( .A(n25652), .B(reg_file[837]), .C(n25663), .D(reg_file[965]), .Y(n32454) );
  NOR2X1 U19735 ( .A(n32459), .B(n32460), .Y(n32445) );
  NAND3X1 U19736 ( .A(n32461), .B(n32462), .C(n32463), .Y(n32460) );
  NOR2X1 U19737 ( .A(n32464), .B(n32465), .Y(n32463) );
  OAI22X1 U19738 ( .A(n27585), .B(n25674), .C(n27586), .D(n25685), .Y(n32465)
         );
  OAI22X1 U19739 ( .A(n27587), .B(n25695), .C(n27588), .D(n25706), .Y(n32464)
         );
  AOI22X1 U19740 ( .A(n25716), .B(reg_file[3525]), .C(n25727), .D(
        reg_file[3397]), .Y(n32462) );
  AOI22X1 U19741 ( .A(n25738), .B(reg_file[3269]), .C(n25749), .D(
        reg_file[3141]), .Y(n32461) );
  NAND3X1 U19742 ( .A(n32466), .B(n32467), .C(n32468), .Y(n32459) );
  NOR2X1 U19743 ( .A(n32469), .B(n32470), .Y(n32468) );
  OAI22X1 U19744 ( .A(n27594), .B(n25760), .C(n27595), .D(n25771), .Y(n32470)
         );
  OAI22X1 U19745 ( .A(n27596), .B(n25781), .C(n27597), .D(n25792), .Y(n32469)
         );
  AOI22X1 U19746 ( .A(n25802), .B(reg_file[2501]), .C(n25813), .D(
        reg_file[2373]), .Y(n32467) );
  AOI22X1 U19747 ( .A(n25824), .B(reg_file[2245]), .C(n25835), .D(
        reg_file[2117]), .Y(n32466) );
  AOI21X1 U19748 ( .A(n32471), .B(n32472), .C(n25491), .Y(rd1data1033_68_) );
  NOR2X1 U19749 ( .A(n32473), .B(n32474), .Y(n32472) );
  NAND3X1 U19750 ( .A(n32475), .B(n32476), .C(n32477), .Y(n32474) );
  NOR2X1 U19751 ( .A(n32478), .B(n32479), .Y(n32477) );
  OAI22X1 U19752 ( .A(n27607), .B(n25502), .C(n27608), .D(n25513), .Y(n32479)
         );
  OAI22X1 U19753 ( .A(n27609), .B(n25523), .C(n27610), .D(n25534), .Y(n32478)
         );
  AOI22X1 U19754 ( .A(n25544), .B(reg_file[1476]), .C(n25555), .D(
        reg_file[1348]), .Y(n32476) );
  AOI22X1 U19755 ( .A(n25566), .B(reg_file[1220]), .C(n25577), .D(
        reg_file[1092]), .Y(n32475) );
  NAND3X1 U19756 ( .A(n32480), .B(n32481), .C(n32482), .Y(n32473) );
  NOR2X1 U19757 ( .A(n32483), .B(n32484), .Y(n32482) );
  OAI22X1 U19758 ( .A(n27616), .B(n25588), .C(n27617), .D(n25599), .Y(n32484)
         );
  OAI22X1 U19759 ( .A(n27618), .B(n25609), .C(n27619), .D(n25620), .Y(n32483)
         );
  AOI22X1 U19760 ( .A(n25630), .B(reg_file[580]), .C(n25641), .D(reg_file[708]), .Y(n32481) );
  AOI22X1 U19761 ( .A(n25652), .B(reg_file[836]), .C(n25663), .D(reg_file[964]), .Y(n32480) );
  NOR2X1 U19762 ( .A(n32485), .B(n32486), .Y(n32471) );
  NAND3X1 U19763 ( .A(n32487), .B(n32488), .C(n32489), .Y(n32486) );
  NOR2X1 U19764 ( .A(n32490), .B(n32491), .Y(n32489) );
  OAI22X1 U19765 ( .A(n27627), .B(n25674), .C(n27628), .D(n25685), .Y(n32491)
         );
  OAI22X1 U19766 ( .A(n27629), .B(n25695), .C(n27630), .D(n25706), .Y(n32490)
         );
  AOI22X1 U19767 ( .A(n25716), .B(reg_file[3524]), .C(n25727), .D(
        reg_file[3396]), .Y(n32488) );
  AOI22X1 U19768 ( .A(n25738), .B(reg_file[3268]), .C(n25749), .D(
        reg_file[3140]), .Y(n32487) );
  NAND3X1 U19769 ( .A(n32492), .B(n32493), .C(n32494), .Y(n32485) );
  NOR2X1 U19770 ( .A(n32495), .B(n32496), .Y(n32494) );
  OAI22X1 U19771 ( .A(n27636), .B(n25760), .C(n27637), .D(n25771), .Y(n32496)
         );
  OAI22X1 U19772 ( .A(n27638), .B(n25781), .C(n27639), .D(n25792), .Y(n32495)
         );
  AOI22X1 U19773 ( .A(n25802), .B(reg_file[2500]), .C(n25813), .D(
        reg_file[2372]), .Y(n32493) );
  AOI22X1 U19774 ( .A(n25824), .B(reg_file[2244]), .C(n25835), .D(
        reg_file[2116]), .Y(n32492) );
  AOI21X1 U19775 ( .A(n32497), .B(n32498), .C(n25491), .Y(rd1data1033_67_) );
  NOR2X1 U19776 ( .A(n32499), .B(n32500), .Y(n32498) );
  NAND3X1 U19777 ( .A(n32501), .B(n32502), .C(n32503), .Y(n32500) );
  NOR2X1 U19778 ( .A(n32504), .B(n32505), .Y(n32503) );
  OAI22X1 U19779 ( .A(n27649), .B(n25502), .C(n27650), .D(n25513), .Y(n32505)
         );
  OAI22X1 U19780 ( .A(n27651), .B(n25523), .C(n27652), .D(n25534), .Y(n32504)
         );
  AOI22X1 U19781 ( .A(n25544), .B(reg_file[1475]), .C(n25555), .D(
        reg_file[1347]), .Y(n32502) );
  AOI22X1 U19782 ( .A(n25566), .B(reg_file[1219]), .C(n25577), .D(
        reg_file[1091]), .Y(n32501) );
  NAND3X1 U19783 ( .A(n32506), .B(n32507), .C(n32508), .Y(n32499) );
  NOR2X1 U19784 ( .A(n32509), .B(n32510), .Y(n32508) );
  OAI22X1 U19785 ( .A(n27658), .B(n25588), .C(n27659), .D(n25599), .Y(n32510)
         );
  OAI22X1 U19786 ( .A(n27660), .B(n25609), .C(n27661), .D(n25620), .Y(n32509)
         );
  AOI22X1 U19787 ( .A(n25630), .B(reg_file[579]), .C(n25641), .D(reg_file[707]), .Y(n32507) );
  AOI22X1 U19788 ( .A(n25652), .B(reg_file[835]), .C(n25663), .D(reg_file[963]), .Y(n32506) );
  NOR2X1 U19789 ( .A(n32511), .B(n32512), .Y(n32497) );
  NAND3X1 U19790 ( .A(n32513), .B(n32514), .C(n32515), .Y(n32512) );
  NOR2X1 U19791 ( .A(n32516), .B(n32517), .Y(n32515) );
  OAI22X1 U19792 ( .A(n27669), .B(n25674), .C(n27670), .D(n25685), .Y(n32517)
         );
  OAI22X1 U19793 ( .A(n27671), .B(n25695), .C(n27672), .D(n25706), .Y(n32516)
         );
  AOI22X1 U19794 ( .A(n25716), .B(reg_file[3523]), .C(n25727), .D(
        reg_file[3395]), .Y(n32514) );
  AOI22X1 U19795 ( .A(n25738), .B(reg_file[3267]), .C(n25749), .D(
        reg_file[3139]), .Y(n32513) );
  NAND3X1 U19796 ( .A(n32518), .B(n32519), .C(n32520), .Y(n32511) );
  NOR2X1 U19797 ( .A(n32521), .B(n32522), .Y(n32520) );
  OAI22X1 U19798 ( .A(n27678), .B(n25760), .C(n27679), .D(n25771), .Y(n32522)
         );
  OAI22X1 U19799 ( .A(n27680), .B(n25781), .C(n27681), .D(n25792), .Y(n32521)
         );
  AOI22X1 U19800 ( .A(n25802), .B(reg_file[2499]), .C(n25813), .D(
        reg_file[2371]), .Y(n32519) );
  AOI22X1 U19801 ( .A(n25824), .B(reg_file[2243]), .C(n25835), .D(
        reg_file[2115]), .Y(n32518) );
  AOI21X1 U19802 ( .A(n32523), .B(n32524), .C(n25491), .Y(rd1data1033_66_) );
  NOR2X1 U19803 ( .A(n32525), .B(n32526), .Y(n32524) );
  NAND3X1 U19804 ( .A(n32527), .B(n32528), .C(n32529), .Y(n32526) );
  NOR2X1 U19805 ( .A(n32530), .B(n32531), .Y(n32529) );
  OAI22X1 U19806 ( .A(n27691), .B(n25502), .C(n27692), .D(n25512), .Y(n32531)
         );
  OAI22X1 U19807 ( .A(n27693), .B(n25523), .C(n27694), .D(n25533), .Y(n32530)
         );
  AOI22X1 U19808 ( .A(n25544), .B(reg_file[1474]), .C(n25555), .D(
        reg_file[1346]), .Y(n32528) );
  AOI22X1 U19809 ( .A(n25566), .B(reg_file[1218]), .C(n25577), .D(
        reg_file[1090]), .Y(n32527) );
  NAND3X1 U19810 ( .A(n32532), .B(n32533), .C(n32534), .Y(n32525) );
  NOR2X1 U19811 ( .A(n32535), .B(n32536), .Y(n32534) );
  OAI22X1 U19812 ( .A(n27700), .B(n25588), .C(n27701), .D(n25598), .Y(n32536)
         );
  OAI22X1 U19813 ( .A(n27702), .B(n25609), .C(n27703), .D(n25619), .Y(n32535)
         );
  AOI22X1 U19814 ( .A(n25630), .B(reg_file[578]), .C(n25641), .D(reg_file[706]), .Y(n32533) );
  AOI22X1 U19815 ( .A(n25652), .B(reg_file[834]), .C(n25663), .D(reg_file[962]), .Y(n32532) );
  NOR2X1 U19816 ( .A(n32537), .B(n32538), .Y(n32523) );
  NAND3X1 U19817 ( .A(n32539), .B(n32540), .C(n32541), .Y(n32538) );
  NOR2X1 U19818 ( .A(n32542), .B(n32543), .Y(n32541) );
  OAI22X1 U19819 ( .A(n27711), .B(n25674), .C(n27712), .D(n25684), .Y(n32543)
         );
  OAI22X1 U19820 ( .A(n27713), .B(n25695), .C(n27714), .D(n25705), .Y(n32542)
         );
  AOI22X1 U19821 ( .A(n25716), .B(reg_file[3522]), .C(n25727), .D(
        reg_file[3394]), .Y(n32540) );
  AOI22X1 U19822 ( .A(n25738), .B(reg_file[3266]), .C(n25749), .D(
        reg_file[3138]), .Y(n32539) );
  NAND3X1 U19823 ( .A(n32544), .B(n32545), .C(n32546), .Y(n32537) );
  NOR2X1 U19824 ( .A(n32547), .B(n32548), .Y(n32546) );
  OAI22X1 U19825 ( .A(n27720), .B(n25760), .C(n27721), .D(n25770), .Y(n32548)
         );
  OAI22X1 U19826 ( .A(n27722), .B(n25781), .C(n27723), .D(n25791), .Y(n32547)
         );
  AOI22X1 U19827 ( .A(n25802), .B(reg_file[2498]), .C(n25813), .D(
        reg_file[2370]), .Y(n32545) );
  AOI22X1 U19828 ( .A(n25824), .B(reg_file[2242]), .C(n25835), .D(
        reg_file[2114]), .Y(n32544) );
  AOI21X1 U19829 ( .A(n32549), .B(n32550), .C(n25491), .Y(rd1data1033_65_) );
  NOR2X1 U19830 ( .A(n32551), .B(n32552), .Y(n32550) );
  NAND3X1 U19831 ( .A(n32553), .B(n32554), .C(n32555), .Y(n32552) );
  NOR2X1 U19832 ( .A(n32556), .B(n32557), .Y(n32555) );
  OAI22X1 U19833 ( .A(n27733), .B(n25502), .C(n27734), .D(n25512), .Y(n32557)
         );
  OAI22X1 U19834 ( .A(n27735), .B(n25523), .C(n27736), .D(n25533), .Y(n32556)
         );
  AOI22X1 U19835 ( .A(n25544), .B(reg_file[1473]), .C(n25555), .D(
        reg_file[1345]), .Y(n32554) );
  AOI22X1 U19836 ( .A(n25566), .B(reg_file[1217]), .C(n25577), .D(
        reg_file[1089]), .Y(n32553) );
  NAND3X1 U19837 ( .A(n32558), .B(n32559), .C(n32560), .Y(n32551) );
  NOR2X1 U19838 ( .A(n32561), .B(n32562), .Y(n32560) );
  OAI22X1 U19839 ( .A(n27742), .B(n25588), .C(n27743), .D(n25598), .Y(n32562)
         );
  OAI22X1 U19840 ( .A(n27744), .B(n25609), .C(n27745), .D(n25619), .Y(n32561)
         );
  AOI22X1 U19841 ( .A(n25630), .B(reg_file[577]), .C(n25641), .D(reg_file[705]), .Y(n32559) );
  AOI22X1 U19842 ( .A(n25652), .B(reg_file[833]), .C(n25663), .D(reg_file[961]), .Y(n32558) );
  NOR2X1 U19843 ( .A(n32563), .B(n32564), .Y(n32549) );
  NAND3X1 U19844 ( .A(n32565), .B(n32566), .C(n32567), .Y(n32564) );
  NOR2X1 U19845 ( .A(n32568), .B(n32569), .Y(n32567) );
  OAI22X1 U19846 ( .A(n27753), .B(n25674), .C(n27754), .D(n25684), .Y(n32569)
         );
  OAI22X1 U19847 ( .A(n27755), .B(n25695), .C(n27756), .D(n25705), .Y(n32568)
         );
  AOI22X1 U19848 ( .A(n25716), .B(reg_file[3521]), .C(n25727), .D(
        reg_file[3393]), .Y(n32566) );
  AOI22X1 U19849 ( .A(n25738), .B(reg_file[3265]), .C(n25749), .D(
        reg_file[3137]), .Y(n32565) );
  NAND3X1 U19850 ( .A(n32570), .B(n32571), .C(n32572), .Y(n32563) );
  NOR2X1 U19851 ( .A(n32573), .B(n32574), .Y(n32572) );
  OAI22X1 U19852 ( .A(n27762), .B(n25760), .C(n27763), .D(n25770), .Y(n32574)
         );
  OAI22X1 U19853 ( .A(n27764), .B(n25781), .C(n27765), .D(n25791), .Y(n32573)
         );
  AOI22X1 U19854 ( .A(n25802), .B(reg_file[2497]), .C(n25813), .D(
        reg_file[2369]), .Y(n32571) );
  AOI22X1 U19855 ( .A(n25824), .B(reg_file[2241]), .C(n25835), .D(
        reg_file[2113]), .Y(n32570) );
  AOI21X1 U19856 ( .A(n32575), .B(n32576), .C(n25491), .Y(rd1data1033_64_) );
  NOR2X1 U19857 ( .A(n32577), .B(n32578), .Y(n32576) );
  NAND3X1 U19858 ( .A(n32579), .B(n32580), .C(n32581), .Y(n32578) );
  NOR2X1 U19859 ( .A(n32582), .B(n32583), .Y(n32581) );
  OAI22X1 U19860 ( .A(n27775), .B(n25502), .C(n27776), .D(n25512), .Y(n32583)
         );
  OAI22X1 U19861 ( .A(n27777), .B(n25523), .C(n27778), .D(n25533), .Y(n32582)
         );
  AOI22X1 U19862 ( .A(n25544), .B(reg_file[1472]), .C(n25555), .D(
        reg_file[1344]), .Y(n32580) );
  AOI22X1 U19863 ( .A(n25566), .B(reg_file[1216]), .C(n25577), .D(
        reg_file[1088]), .Y(n32579) );
  NAND3X1 U19864 ( .A(n32584), .B(n32585), .C(n32586), .Y(n32577) );
  NOR2X1 U19865 ( .A(n32587), .B(n32588), .Y(n32586) );
  OAI22X1 U19866 ( .A(n27784), .B(n25588), .C(n27785), .D(n25598), .Y(n32588)
         );
  OAI22X1 U19867 ( .A(n27786), .B(n25609), .C(n27787), .D(n25619), .Y(n32587)
         );
  AOI22X1 U19868 ( .A(n25630), .B(reg_file[576]), .C(n25641), .D(reg_file[704]), .Y(n32585) );
  AOI22X1 U19869 ( .A(n25652), .B(reg_file[832]), .C(n25663), .D(reg_file[960]), .Y(n32584) );
  NOR2X1 U19870 ( .A(n32589), .B(n32590), .Y(n32575) );
  NAND3X1 U19871 ( .A(n32591), .B(n32592), .C(n32593), .Y(n32590) );
  NOR2X1 U19872 ( .A(n32594), .B(n32595), .Y(n32593) );
  OAI22X1 U19873 ( .A(n27795), .B(n25674), .C(n27796), .D(n25684), .Y(n32595)
         );
  OAI22X1 U19874 ( .A(n27797), .B(n25695), .C(n27798), .D(n25705), .Y(n32594)
         );
  AOI22X1 U19875 ( .A(n25716), .B(reg_file[3520]), .C(n25727), .D(
        reg_file[3392]), .Y(n32592) );
  AOI22X1 U19876 ( .A(n25738), .B(reg_file[3264]), .C(n25749), .D(
        reg_file[3136]), .Y(n32591) );
  NAND3X1 U19877 ( .A(n32596), .B(n32597), .C(n32598), .Y(n32589) );
  NOR2X1 U19878 ( .A(n32599), .B(n32600), .Y(n32598) );
  OAI22X1 U19879 ( .A(n27804), .B(n25760), .C(n27805), .D(n25770), .Y(n32600)
         );
  OAI22X1 U19880 ( .A(n27806), .B(n25781), .C(n27807), .D(n25791), .Y(n32599)
         );
  AOI22X1 U19881 ( .A(n25802), .B(reg_file[2496]), .C(n25813), .D(
        reg_file[2368]), .Y(n32597) );
  AOI22X1 U19882 ( .A(n25824), .B(reg_file[2240]), .C(n25835), .D(
        reg_file[2112]), .Y(n32596) );
  AOI21X1 U19883 ( .A(n32601), .B(n32602), .C(n25491), .Y(rd1data1033_63_) );
  NOR2X1 U19884 ( .A(n32603), .B(n32604), .Y(n32602) );
  NAND3X1 U19885 ( .A(n32605), .B(n32606), .C(n32607), .Y(n32604) );
  NOR2X1 U19886 ( .A(n32608), .B(n32609), .Y(n32607) );
  OAI22X1 U19887 ( .A(n27817), .B(n25502), .C(n27818), .D(n25512), .Y(n32609)
         );
  OAI22X1 U19888 ( .A(n27819), .B(n25523), .C(n27820), .D(n25533), .Y(n32608)
         );
  AOI22X1 U19889 ( .A(n25544), .B(reg_file[1471]), .C(n25555), .D(
        reg_file[1343]), .Y(n32606) );
  AOI22X1 U19890 ( .A(n25566), .B(reg_file[1215]), .C(n25577), .D(
        reg_file[1087]), .Y(n32605) );
  NAND3X1 U19891 ( .A(n32610), .B(n32611), .C(n32612), .Y(n32603) );
  NOR2X1 U19892 ( .A(n32613), .B(n32614), .Y(n32612) );
  OAI22X1 U19893 ( .A(n27826), .B(n25588), .C(n27827), .D(n25598), .Y(n32614)
         );
  OAI22X1 U19894 ( .A(n27828), .B(n25609), .C(n27829), .D(n25619), .Y(n32613)
         );
  AOI22X1 U19895 ( .A(n25630), .B(reg_file[575]), .C(n25641), .D(reg_file[703]), .Y(n32611) );
  AOI22X1 U19896 ( .A(n25652), .B(reg_file[831]), .C(n25663), .D(reg_file[959]), .Y(n32610) );
  NOR2X1 U19897 ( .A(n32615), .B(n32616), .Y(n32601) );
  NAND3X1 U19898 ( .A(n32617), .B(n32618), .C(n32619), .Y(n32616) );
  NOR2X1 U19899 ( .A(n32620), .B(n32621), .Y(n32619) );
  OAI22X1 U19900 ( .A(n27837), .B(n25674), .C(n27838), .D(n25684), .Y(n32621)
         );
  OAI22X1 U19901 ( .A(n27839), .B(n25695), .C(n27840), .D(n25705), .Y(n32620)
         );
  AOI22X1 U19902 ( .A(n25716), .B(reg_file[3519]), .C(n25727), .D(
        reg_file[3391]), .Y(n32618) );
  AOI22X1 U19903 ( .A(n25738), .B(reg_file[3263]), .C(n25749), .D(
        reg_file[3135]), .Y(n32617) );
  NAND3X1 U19904 ( .A(n32622), .B(n32623), .C(n32624), .Y(n32615) );
  NOR2X1 U19905 ( .A(n32625), .B(n32626), .Y(n32624) );
  OAI22X1 U19906 ( .A(n27846), .B(n25760), .C(n27847), .D(n25770), .Y(n32626)
         );
  OAI22X1 U19907 ( .A(n27848), .B(n25781), .C(n27849), .D(n25791), .Y(n32625)
         );
  AOI22X1 U19908 ( .A(n25802), .B(reg_file[2495]), .C(n25813), .D(
        reg_file[2367]), .Y(n32623) );
  AOI22X1 U19909 ( .A(n25824), .B(reg_file[2239]), .C(n25835), .D(
        reg_file[2111]), .Y(n32622) );
  AOI21X1 U19910 ( .A(n32627), .B(n32628), .C(n25491), .Y(rd1data1033_62_) );
  NOR2X1 U19911 ( .A(n32629), .B(n32630), .Y(n32628) );
  NAND3X1 U19912 ( .A(n32631), .B(n32632), .C(n32633), .Y(n32630) );
  NOR2X1 U19913 ( .A(n32634), .B(n32635), .Y(n32633) );
  OAI22X1 U19914 ( .A(n27859), .B(n25502), .C(n27860), .D(n25512), .Y(n32635)
         );
  OAI22X1 U19915 ( .A(n27861), .B(n25523), .C(n27862), .D(n25533), .Y(n32634)
         );
  AOI22X1 U19916 ( .A(n25544), .B(reg_file[1470]), .C(n25555), .D(
        reg_file[1342]), .Y(n32632) );
  AOI22X1 U19917 ( .A(n25566), .B(reg_file[1214]), .C(n25577), .D(
        reg_file[1086]), .Y(n32631) );
  NAND3X1 U19918 ( .A(n32636), .B(n32637), .C(n32638), .Y(n32629) );
  NOR2X1 U19919 ( .A(n32639), .B(n32640), .Y(n32638) );
  OAI22X1 U19920 ( .A(n27868), .B(n25588), .C(n27869), .D(n25598), .Y(n32640)
         );
  OAI22X1 U19921 ( .A(n27870), .B(n25609), .C(n27871), .D(n25619), .Y(n32639)
         );
  AOI22X1 U19922 ( .A(n25630), .B(reg_file[574]), .C(n25641), .D(reg_file[702]), .Y(n32637) );
  AOI22X1 U19923 ( .A(n25652), .B(reg_file[830]), .C(n25663), .D(reg_file[958]), .Y(n32636) );
  NOR2X1 U19924 ( .A(n32641), .B(n32642), .Y(n32627) );
  NAND3X1 U19925 ( .A(n32643), .B(n32644), .C(n32645), .Y(n32642) );
  NOR2X1 U19926 ( .A(n32646), .B(n32647), .Y(n32645) );
  OAI22X1 U19927 ( .A(n27879), .B(n25674), .C(n27880), .D(n25684), .Y(n32647)
         );
  OAI22X1 U19928 ( .A(n27881), .B(n25695), .C(n27882), .D(n25705), .Y(n32646)
         );
  AOI22X1 U19929 ( .A(n25716), .B(reg_file[3518]), .C(n25727), .D(
        reg_file[3390]), .Y(n32644) );
  AOI22X1 U19930 ( .A(n25738), .B(reg_file[3262]), .C(n25749), .D(
        reg_file[3134]), .Y(n32643) );
  NAND3X1 U19931 ( .A(n32648), .B(n32649), .C(n32650), .Y(n32641) );
  NOR2X1 U19932 ( .A(n32651), .B(n32652), .Y(n32650) );
  OAI22X1 U19933 ( .A(n27888), .B(n25760), .C(n27889), .D(n25770), .Y(n32652)
         );
  OAI22X1 U19934 ( .A(n27890), .B(n25781), .C(n27891), .D(n25791), .Y(n32651)
         );
  AOI22X1 U19935 ( .A(n25802), .B(reg_file[2494]), .C(n25813), .D(
        reg_file[2366]), .Y(n32649) );
  AOI22X1 U19936 ( .A(n25824), .B(reg_file[2238]), .C(n25835), .D(
        reg_file[2110]), .Y(n32648) );
  AOI21X1 U19937 ( .A(n32653), .B(n32654), .C(n25491), .Y(rd1data1033_61_) );
  NOR2X1 U19938 ( .A(n32655), .B(n32656), .Y(n32654) );
  NAND3X1 U19939 ( .A(n32657), .B(n32658), .C(n32659), .Y(n32656) );
  NOR2X1 U19940 ( .A(n32660), .B(n32661), .Y(n32659) );
  OAI22X1 U19941 ( .A(n27901), .B(n25502), .C(n27902), .D(n25512), .Y(n32661)
         );
  OAI22X1 U19942 ( .A(n27903), .B(n25523), .C(n27904), .D(n25533), .Y(n32660)
         );
  AOI22X1 U19943 ( .A(n25544), .B(reg_file[1469]), .C(n25555), .D(
        reg_file[1341]), .Y(n32658) );
  AOI22X1 U19944 ( .A(n25566), .B(reg_file[1213]), .C(n25577), .D(
        reg_file[1085]), .Y(n32657) );
  NAND3X1 U19945 ( .A(n32662), .B(n32663), .C(n32664), .Y(n32655) );
  NOR2X1 U19946 ( .A(n32665), .B(n32666), .Y(n32664) );
  OAI22X1 U19947 ( .A(n27910), .B(n25588), .C(n27911), .D(n25598), .Y(n32666)
         );
  OAI22X1 U19948 ( .A(n27912), .B(n25609), .C(n27913), .D(n25619), .Y(n32665)
         );
  AOI22X1 U19949 ( .A(n25630), .B(reg_file[573]), .C(n25641), .D(reg_file[701]), .Y(n32663) );
  AOI22X1 U19950 ( .A(n25652), .B(reg_file[829]), .C(n25663), .D(reg_file[957]), .Y(n32662) );
  NOR2X1 U19951 ( .A(n32667), .B(n32668), .Y(n32653) );
  NAND3X1 U19952 ( .A(n32669), .B(n32670), .C(n32671), .Y(n32668) );
  NOR2X1 U19953 ( .A(n32672), .B(n32673), .Y(n32671) );
  OAI22X1 U19954 ( .A(n27921), .B(n25674), .C(n27922), .D(n25684), .Y(n32673)
         );
  OAI22X1 U19955 ( .A(n27923), .B(n25695), .C(n27924), .D(n25705), .Y(n32672)
         );
  AOI22X1 U19956 ( .A(n25716), .B(reg_file[3517]), .C(n25727), .D(
        reg_file[3389]), .Y(n32670) );
  AOI22X1 U19957 ( .A(n25738), .B(reg_file[3261]), .C(n25749), .D(
        reg_file[3133]), .Y(n32669) );
  NAND3X1 U19958 ( .A(n32674), .B(n32675), .C(n32676), .Y(n32667) );
  NOR2X1 U19959 ( .A(n32677), .B(n32678), .Y(n32676) );
  OAI22X1 U19960 ( .A(n27930), .B(n25760), .C(n27931), .D(n25770), .Y(n32678)
         );
  OAI22X1 U19961 ( .A(n27932), .B(n25781), .C(n27933), .D(n25791), .Y(n32677)
         );
  AOI22X1 U19962 ( .A(n25802), .B(reg_file[2493]), .C(n25813), .D(
        reg_file[2365]), .Y(n32675) );
  AOI22X1 U19963 ( .A(n25824), .B(reg_file[2237]), .C(n25835), .D(
        reg_file[2109]), .Y(n32674) );
  AOI21X1 U19964 ( .A(n32679), .B(n32680), .C(n25491), .Y(rd1data1033_60_) );
  NOR2X1 U19965 ( .A(n32681), .B(n32682), .Y(n32680) );
  NAND3X1 U19966 ( .A(n32683), .B(n32684), .C(n32685), .Y(n32682) );
  NOR2X1 U19967 ( .A(n32686), .B(n32687), .Y(n32685) );
  OAI22X1 U19968 ( .A(n27943), .B(n25502), .C(n27944), .D(n25512), .Y(n32687)
         );
  OAI22X1 U19969 ( .A(n27945), .B(n25523), .C(n27946), .D(n25533), .Y(n32686)
         );
  AOI22X1 U19970 ( .A(n25544), .B(reg_file[1468]), .C(n25555), .D(
        reg_file[1340]), .Y(n32684) );
  AOI22X1 U19971 ( .A(n25566), .B(reg_file[1212]), .C(n25577), .D(
        reg_file[1084]), .Y(n32683) );
  NAND3X1 U19972 ( .A(n32688), .B(n32689), .C(n32690), .Y(n32681) );
  NOR2X1 U19973 ( .A(n32691), .B(n32692), .Y(n32690) );
  OAI22X1 U19974 ( .A(n27952), .B(n25588), .C(n27953), .D(n25598), .Y(n32692)
         );
  OAI22X1 U19975 ( .A(n27954), .B(n25609), .C(n27955), .D(n25619), .Y(n32691)
         );
  AOI22X1 U19976 ( .A(n25630), .B(reg_file[572]), .C(n25641), .D(reg_file[700]), .Y(n32689) );
  AOI22X1 U19977 ( .A(n25652), .B(reg_file[828]), .C(n25663), .D(reg_file[956]), .Y(n32688) );
  NOR2X1 U19978 ( .A(n32693), .B(n32694), .Y(n32679) );
  NAND3X1 U19979 ( .A(n32695), .B(n32696), .C(n32697), .Y(n32694) );
  NOR2X1 U19980 ( .A(n32698), .B(n32699), .Y(n32697) );
  OAI22X1 U19981 ( .A(n27963), .B(n25674), .C(n27964), .D(n25684), .Y(n32699)
         );
  OAI22X1 U19982 ( .A(n27965), .B(n25695), .C(n27966), .D(n25705), .Y(n32698)
         );
  AOI22X1 U19983 ( .A(n25716), .B(reg_file[3516]), .C(n25727), .D(
        reg_file[3388]), .Y(n32696) );
  AOI22X1 U19984 ( .A(n25738), .B(reg_file[3260]), .C(n25749), .D(
        reg_file[3132]), .Y(n32695) );
  NAND3X1 U19985 ( .A(n32700), .B(n32701), .C(n32702), .Y(n32693) );
  NOR2X1 U19986 ( .A(n32703), .B(n32704), .Y(n32702) );
  OAI22X1 U19987 ( .A(n27972), .B(n25760), .C(n27973), .D(n25770), .Y(n32704)
         );
  OAI22X1 U19988 ( .A(n27974), .B(n25781), .C(n27975), .D(n25791), .Y(n32703)
         );
  AOI22X1 U19989 ( .A(n25802), .B(reg_file[2492]), .C(n25813), .D(
        reg_file[2364]), .Y(n32701) );
  AOI22X1 U19990 ( .A(n25824), .B(reg_file[2236]), .C(n25835), .D(
        reg_file[2108]), .Y(n32700) );
  AOI21X1 U19991 ( .A(n32705), .B(n32706), .C(n25490), .Y(rd1data1033_5_) );
  NOR2X1 U19992 ( .A(n32707), .B(n32708), .Y(n32706) );
  NAND3X1 U19993 ( .A(n32709), .B(n32710), .C(n32711), .Y(n32708) );
  NOR2X1 U19994 ( .A(n32712), .B(n32713), .Y(n32711) );
  OAI22X1 U19995 ( .A(n27985), .B(n25501), .C(n27986), .D(n25512), .Y(n32713)
         );
  OAI22X1 U19996 ( .A(n27987), .B(n25522), .C(n27988), .D(n25533), .Y(n32712)
         );
  AOI22X1 U19997 ( .A(n25543), .B(reg_file[1413]), .C(n25554), .D(
        reg_file[1285]), .Y(n32710) );
  AOI22X1 U19998 ( .A(n25565), .B(reg_file[1157]), .C(n25576), .D(
        reg_file[1029]), .Y(n32709) );
  NAND3X1 U19999 ( .A(n32714), .B(n32715), .C(n32716), .Y(n32707) );
  NOR2X1 U20000 ( .A(n32717), .B(n32718), .Y(n32716) );
  OAI22X1 U20001 ( .A(n27994), .B(n25587), .C(n27995), .D(n25598), .Y(n32718)
         );
  OAI22X1 U20002 ( .A(n27996), .B(n25608), .C(n27997), .D(n25619), .Y(n32717)
         );
  AOI22X1 U20003 ( .A(n25629), .B(reg_file[517]), .C(n25640), .D(reg_file[645]), .Y(n32715) );
  AOI22X1 U20004 ( .A(n25651), .B(reg_file[773]), .C(n25662), .D(reg_file[901]), .Y(n32714) );
  NOR2X1 U20005 ( .A(n32719), .B(n32720), .Y(n32705) );
  NAND3X1 U20006 ( .A(n32721), .B(n32722), .C(n32723), .Y(n32720) );
  NOR2X1 U20007 ( .A(n32724), .B(n32725), .Y(n32723) );
  OAI22X1 U20008 ( .A(n28005), .B(n25673), .C(n28006), .D(n25684), .Y(n32725)
         );
  OAI22X1 U20009 ( .A(n28007), .B(n25694), .C(n28008), .D(n25705), .Y(n32724)
         );
  AOI22X1 U20010 ( .A(n25715), .B(reg_file[3461]), .C(n25726), .D(
        reg_file[3333]), .Y(n32722) );
  AOI22X1 U20011 ( .A(n25737), .B(reg_file[3205]), .C(n25748), .D(
        reg_file[3077]), .Y(n32721) );
  NAND3X1 U20012 ( .A(n32726), .B(n32727), .C(n32728), .Y(n32719) );
  NOR2X1 U20013 ( .A(n32729), .B(n32730), .Y(n32728) );
  OAI22X1 U20014 ( .A(n28014), .B(n25759), .C(n28015), .D(n25770), .Y(n32730)
         );
  OAI22X1 U20015 ( .A(n28016), .B(n25780), .C(n28017), .D(n25791), .Y(n32729)
         );
  AOI22X1 U20016 ( .A(n25801), .B(reg_file[2437]), .C(n25812), .D(
        reg_file[2309]), .Y(n32727) );
  AOI22X1 U20017 ( .A(n25823), .B(reg_file[2181]), .C(n25834), .D(
        reg_file[2053]), .Y(n32726) );
  AOI21X1 U20018 ( .A(n32731), .B(n32732), .C(n25490), .Y(rd1data1033_59_) );
  NOR2X1 U20019 ( .A(n32733), .B(n32734), .Y(n32732) );
  NAND3X1 U20020 ( .A(n32735), .B(n32736), .C(n32737), .Y(n32734) );
  NOR2X1 U20021 ( .A(n32738), .B(n32739), .Y(n32737) );
  OAI22X1 U20022 ( .A(n28027), .B(n25501), .C(n28028), .D(n25512), .Y(n32739)
         );
  OAI22X1 U20023 ( .A(n28029), .B(n25522), .C(n28030), .D(n25533), .Y(n32738)
         );
  AOI22X1 U20024 ( .A(n25543), .B(reg_file[1467]), .C(n25554), .D(
        reg_file[1339]), .Y(n32736) );
  AOI22X1 U20025 ( .A(n25565), .B(reg_file[1211]), .C(n25576), .D(
        reg_file[1083]), .Y(n32735) );
  NAND3X1 U20026 ( .A(n32740), .B(n32741), .C(n32742), .Y(n32733) );
  NOR2X1 U20027 ( .A(n32743), .B(n32744), .Y(n32742) );
  OAI22X1 U20028 ( .A(n28036), .B(n25587), .C(n28037), .D(n25598), .Y(n32744)
         );
  OAI22X1 U20029 ( .A(n28038), .B(n25608), .C(n28039), .D(n25619), .Y(n32743)
         );
  AOI22X1 U20030 ( .A(n25629), .B(reg_file[571]), .C(n25640), .D(reg_file[699]), .Y(n32741) );
  AOI22X1 U20031 ( .A(n25651), .B(reg_file[827]), .C(n25662), .D(reg_file[955]), .Y(n32740) );
  NOR2X1 U20032 ( .A(n32745), .B(n32746), .Y(n32731) );
  NAND3X1 U20033 ( .A(n32747), .B(n32748), .C(n32749), .Y(n32746) );
  NOR2X1 U20034 ( .A(n32750), .B(n32751), .Y(n32749) );
  OAI22X1 U20035 ( .A(n28047), .B(n25673), .C(n28048), .D(n25684), .Y(n32751)
         );
  OAI22X1 U20036 ( .A(n28049), .B(n25694), .C(n28050), .D(n25705), .Y(n32750)
         );
  AOI22X1 U20037 ( .A(n25715), .B(reg_file[3515]), .C(n25726), .D(
        reg_file[3387]), .Y(n32748) );
  AOI22X1 U20038 ( .A(n25737), .B(reg_file[3259]), .C(n25748), .D(
        reg_file[3131]), .Y(n32747) );
  NAND3X1 U20039 ( .A(n32752), .B(n32753), .C(n32754), .Y(n32745) );
  NOR2X1 U20040 ( .A(n32755), .B(n32756), .Y(n32754) );
  OAI22X1 U20041 ( .A(n28056), .B(n25759), .C(n28057), .D(n25770), .Y(n32756)
         );
  OAI22X1 U20042 ( .A(n28058), .B(n25780), .C(n28059), .D(n25791), .Y(n32755)
         );
  AOI22X1 U20043 ( .A(n25801), .B(reg_file[2491]), .C(n25812), .D(
        reg_file[2363]), .Y(n32753) );
  AOI22X1 U20044 ( .A(n25823), .B(reg_file[2235]), .C(n25834), .D(
        reg_file[2107]), .Y(n32752) );
  AOI21X1 U20045 ( .A(n32757), .B(n32758), .C(n25490), .Y(rd1data1033_58_) );
  NOR2X1 U20046 ( .A(n32759), .B(n32760), .Y(n32758) );
  NAND3X1 U20047 ( .A(n32761), .B(n32762), .C(n32763), .Y(n32760) );
  NOR2X1 U20048 ( .A(n32764), .B(n32765), .Y(n32763) );
  OAI22X1 U20049 ( .A(n28069), .B(n25501), .C(n28070), .D(n25512), .Y(n32765)
         );
  OAI22X1 U20050 ( .A(n28071), .B(n25522), .C(n28072), .D(n25533), .Y(n32764)
         );
  AOI22X1 U20051 ( .A(n25543), .B(reg_file[1466]), .C(n25554), .D(
        reg_file[1338]), .Y(n32762) );
  AOI22X1 U20052 ( .A(n25565), .B(reg_file[1210]), .C(n25576), .D(
        reg_file[1082]), .Y(n32761) );
  NAND3X1 U20053 ( .A(n32766), .B(n32767), .C(n32768), .Y(n32759) );
  NOR2X1 U20054 ( .A(n32769), .B(n32770), .Y(n32768) );
  OAI22X1 U20055 ( .A(n28078), .B(n25587), .C(n28079), .D(n25598), .Y(n32770)
         );
  OAI22X1 U20056 ( .A(n28080), .B(n25608), .C(n28081), .D(n25619), .Y(n32769)
         );
  AOI22X1 U20057 ( .A(n25629), .B(reg_file[570]), .C(n25640), .D(reg_file[698]), .Y(n32767) );
  AOI22X1 U20058 ( .A(n25651), .B(reg_file[826]), .C(n25662), .D(reg_file[954]), .Y(n32766) );
  NOR2X1 U20059 ( .A(n32771), .B(n32772), .Y(n32757) );
  NAND3X1 U20060 ( .A(n32773), .B(n32774), .C(n32775), .Y(n32772) );
  NOR2X1 U20061 ( .A(n32776), .B(n32777), .Y(n32775) );
  OAI22X1 U20062 ( .A(n28089), .B(n25673), .C(n28090), .D(n25684), .Y(n32777)
         );
  OAI22X1 U20063 ( .A(n28091), .B(n25694), .C(n28092), .D(n25705), .Y(n32776)
         );
  AOI22X1 U20064 ( .A(n25715), .B(reg_file[3514]), .C(n25726), .D(
        reg_file[3386]), .Y(n32774) );
  AOI22X1 U20065 ( .A(n25737), .B(reg_file[3258]), .C(n25748), .D(
        reg_file[3130]), .Y(n32773) );
  NAND3X1 U20066 ( .A(n32778), .B(n32779), .C(n32780), .Y(n32771) );
  NOR2X1 U20067 ( .A(n32781), .B(n32782), .Y(n32780) );
  OAI22X1 U20068 ( .A(n28098), .B(n25759), .C(n28099), .D(n25770), .Y(n32782)
         );
  OAI22X1 U20069 ( .A(n28100), .B(n25780), .C(n28101), .D(n25791), .Y(n32781)
         );
  AOI22X1 U20070 ( .A(n25801), .B(reg_file[2490]), .C(n25812), .D(
        reg_file[2362]), .Y(n32779) );
  AOI22X1 U20071 ( .A(n25823), .B(reg_file[2234]), .C(n25834), .D(
        reg_file[2106]), .Y(n32778) );
  AOI21X1 U20072 ( .A(n32783), .B(n32784), .C(n25490), .Y(rd1data1033_57_) );
  NOR2X1 U20073 ( .A(n32785), .B(n32786), .Y(n32784) );
  NAND3X1 U20074 ( .A(n32787), .B(n32788), .C(n32789), .Y(n32786) );
  NOR2X1 U20075 ( .A(n32790), .B(n32791), .Y(n32789) );
  OAI22X1 U20076 ( .A(n28111), .B(n25501), .C(n28112), .D(n25512), .Y(n32791)
         );
  OAI22X1 U20077 ( .A(n28113), .B(n25522), .C(n28114), .D(n25533), .Y(n32790)
         );
  AOI22X1 U20078 ( .A(n25543), .B(reg_file[1465]), .C(n25554), .D(
        reg_file[1337]), .Y(n32788) );
  AOI22X1 U20079 ( .A(n25565), .B(reg_file[1209]), .C(n25576), .D(
        reg_file[1081]), .Y(n32787) );
  NAND3X1 U20080 ( .A(n32792), .B(n32793), .C(n32794), .Y(n32785) );
  NOR2X1 U20081 ( .A(n32795), .B(n32796), .Y(n32794) );
  OAI22X1 U20082 ( .A(n28120), .B(n25587), .C(n28121), .D(n25598), .Y(n32796)
         );
  OAI22X1 U20083 ( .A(n28122), .B(n25608), .C(n28123), .D(n25619), .Y(n32795)
         );
  AOI22X1 U20084 ( .A(n25629), .B(reg_file[569]), .C(n25640), .D(reg_file[697]), .Y(n32793) );
  AOI22X1 U20085 ( .A(n25651), .B(reg_file[825]), .C(n25662), .D(reg_file[953]), .Y(n32792) );
  NOR2X1 U20086 ( .A(n32797), .B(n32798), .Y(n32783) );
  NAND3X1 U20087 ( .A(n32799), .B(n32800), .C(n32801), .Y(n32798) );
  NOR2X1 U20088 ( .A(n32802), .B(n32803), .Y(n32801) );
  OAI22X1 U20089 ( .A(n28131), .B(n25673), .C(n28132), .D(n25684), .Y(n32803)
         );
  OAI22X1 U20090 ( .A(n28133), .B(n25694), .C(n28134), .D(n25705), .Y(n32802)
         );
  AOI22X1 U20091 ( .A(n25715), .B(reg_file[3513]), .C(n25726), .D(
        reg_file[3385]), .Y(n32800) );
  AOI22X1 U20092 ( .A(n25737), .B(reg_file[3257]), .C(n25748), .D(
        reg_file[3129]), .Y(n32799) );
  NAND3X1 U20093 ( .A(n32804), .B(n32805), .C(n32806), .Y(n32797) );
  NOR2X1 U20094 ( .A(n32807), .B(n32808), .Y(n32806) );
  OAI22X1 U20095 ( .A(n28140), .B(n25759), .C(n28141), .D(n25770), .Y(n32808)
         );
  OAI22X1 U20096 ( .A(n28142), .B(n25780), .C(n28143), .D(n25791), .Y(n32807)
         );
  AOI22X1 U20097 ( .A(n25801), .B(reg_file[2489]), .C(n25812), .D(
        reg_file[2361]), .Y(n32805) );
  AOI22X1 U20098 ( .A(n25823), .B(reg_file[2233]), .C(n25834), .D(
        reg_file[2105]), .Y(n32804) );
  AOI21X1 U20099 ( .A(n32809), .B(n32810), .C(n25490), .Y(rd1data1033_56_) );
  NOR2X1 U20100 ( .A(n32811), .B(n32812), .Y(n32810) );
  NAND3X1 U20101 ( .A(n32813), .B(n32814), .C(n32815), .Y(n32812) );
  NOR2X1 U20102 ( .A(n32816), .B(n32817), .Y(n32815) );
  OAI22X1 U20103 ( .A(n28153), .B(n25501), .C(n28154), .D(n25512), .Y(n32817)
         );
  OAI22X1 U20104 ( .A(n28155), .B(n25522), .C(n28156), .D(n25533), .Y(n32816)
         );
  AOI22X1 U20105 ( .A(n25543), .B(reg_file[1464]), .C(n25554), .D(
        reg_file[1336]), .Y(n32814) );
  AOI22X1 U20106 ( .A(n25565), .B(reg_file[1208]), .C(n25576), .D(
        reg_file[1080]), .Y(n32813) );
  NAND3X1 U20107 ( .A(n32818), .B(n32819), .C(n32820), .Y(n32811) );
  NOR2X1 U20108 ( .A(n32821), .B(n32822), .Y(n32820) );
  OAI22X1 U20109 ( .A(n28162), .B(n25587), .C(n28163), .D(n25598), .Y(n32822)
         );
  OAI22X1 U20110 ( .A(n28164), .B(n25608), .C(n28165), .D(n25619), .Y(n32821)
         );
  AOI22X1 U20111 ( .A(n25629), .B(reg_file[568]), .C(n25640), .D(reg_file[696]), .Y(n32819) );
  AOI22X1 U20112 ( .A(n25651), .B(reg_file[824]), .C(n25662), .D(reg_file[952]), .Y(n32818) );
  NOR2X1 U20113 ( .A(n32823), .B(n32824), .Y(n32809) );
  NAND3X1 U20114 ( .A(n32825), .B(n32826), .C(n32827), .Y(n32824) );
  NOR2X1 U20115 ( .A(n32828), .B(n32829), .Y(n32827) );
  OAI22X1 U20116 ( .A(n28173), .B(n25673), .C(n28174), .D(n25684), .Y(n32829)
         );
  OAI22X1 U20117 ( .A(n28175), .B(n25694), .C(n28176), .D(n25705), .Y(n32828)
         );
  AOI22X1 U20118 ( .A(n25715), .B(reg_file[3512]), .C(n25726), .D(
        reg_file[3384]), .Y(n32826) );
  AOI22X1 U20119 ( .A(n25737), .B(reg_file[3256]), .C(n25748), .D(
        reg_file[3128]), .Y(n32825) );
  NAND3X1 U20120 ( .A(n32830), .B(n32831), .C(n32832), .Y(n32823) );
  NOR2X1 U20121 ( .A(n32833), .B(n32834), .Y(n32832) );
  OAI22X1 U20122 ( .A(n28182), .B(n25759), .C(n28183), .D(n25770), .Y(n32834)
         );
  OAI22X1 U20123 ( .A(n28184), .B(n25780), .C(n28185), .D(n25791), .Y(n32833)
         );
  AOI22X1 U20124 ( .A(n25801), .B(reg_file[2488]), .C(n25812), .D(
        reg_file[2360]), .Y(n32831) );
  AOI22X1 U20125 ( .A(n25823), .B(reg_file[2232]), .C(n25834), .D(
        reg_file[2104]), .Y(n32830) );
  AOI21X1 U20126 ( .A(n32835), .B(n32836), .C(n25490), .Y(rd1data1033_55_) );
  NOR2X1 U20127 ( .A(n32837), .B(n32838), .Y(n32836) );
  NAND3X1 U20128 ( .A(n32839), .B(n32840), .C(n32841), .Y(n32838) );
  NOR2X1 U20129 ( .A(n32842), .B(n32843), .Y(n32841) );
  OAI22X1 U20130 ( .A(n28195), .B(n25501), .C(n28196), .D(n25512), .Y(n32843)
         );
  OAI22X1 U20131 ( .A(n28197), .B(n25522), .C(n28198), .D(n25533), .Y(n32842)
         );
  AOI22X1 U20132 ( .A(n25543), .B(reg_file[1463]), .C(n25554), .D(
        reg_file[1335]), .Y(n32840) );
  AOI22X1 U20133 ( .A(n25565), .B(reg_file[1207]), .C(n25576), .D(
        reg_file[1079]), .Y(n32839) );
  NAND3X1 U20134 ( .A(n32844), .B(n32845), .C(n32846), .Y(n32837) );
  NOR2X1 U20135 ( .A(n32847), .B(n32848), .Y(n32846) );
  OAI22X1 U20136 ( .A(n28204), .B(n25587), .C(n28205), .D(n25598), .Y(n32848)
         );
  OAI22X1 U20137 ( .A(n28206), .B(n25608), .C(n28207), .D(n25619), .Y(n32847)
         );
  AOI22X1 U20138 ( .A(n25629), .B(reg_file[567]), .C(n25640), .D(reg_file[695]), .Y(n32845) );
  AOI22X1 U20139 ( .A(n25651), .B(reg_file[823]), .C(n25662), .D(reg_file[951]), .Y(n32844) );
  NOR2X1 U20140 ( .A(n32849), .B(n32850), .Y(n32835) );
  NAND3X1 U20141 ( .A(n32851), .B(n32852), .C(n32853), .Y(n32850) );
  NOR2X1 U20142 ( .A(n32854), .B(n32855), .Y(n32853) );
  OAI22X1 U20143 ( .A(n28215), .B(n25673), .C(n28216), .D(n25684), .Y(n32855)
         );
  OAI22X1 U20144 ( .A(n28217), .B(n25694), .C(n28218), .D(n25705), .Y(n32854)
         );
  AOI22X1 U20145 ( .A(n25715), .B(reg_file[3511]), .C(n25726), .D(
        reg_file[3383]), .Y(n32852) );
  AOI22X1 U20146 ( .A(n25737), .B(reg_file[3255]), .C(n25748), .D(
        reg_file[3127]), .Y(n32851) );
  NAND3X1 U20147 ( .A(n32856), .B(n32857), .C(n32858), .Y(n32849) );
  NOR2X1 U20148 ( .A(n32859), .B(n32860), .Y(n32858) );
  OAI22X1 U20149 ( .A(n28224), .B(n25759), .C(n28225), .D(n25770), .Y(n32860)
         );
  OAI22X1 U20150 ( .A(n28226), .B(n25780), .C(n28227), .D(n25791), .Y(n32859)
         );
  AOI22X1 U20151 ( .A(n25801), .B(reg_file[2487]), .C(n25812), .D(
        reg_file[2359]), .Y(n32857) );
  AOI22X1 U20152 ( .A(n25823), .B(reg_file[2231]), .C(n25834), .D(
        reg_file[2103]), .Y(n32856) );
  AOI21X1 U20153 ( .A(n32861), .B(n32862), .C(n25490), .Y(rd1data1033_54_) );
  NOR2X1 U20154 ( .A(n32863), .B(n32864), .Y(n32862) );
  NAND3X1 U20155 ( .A(n32865), .B(n32866), .C(n32867), .Y(n32864) );
  NOR2X1 U20156 ( .A(n32868), .B(n32869), .Y(n32867) );
  OAI22X1 U20157 ( .A(n28237), .B(n25501), .C(n28238), .D(n25511), .Y(n32869)
         );
  OAI22X1 U20158 ( .A(n28239), .B(n25522), .C(n28240), .D(n25532), .Y(n32868)
         );
  AOI22X1 U20159 ( .A(n25543), .B(reg_file[1462]), .C(n25554), .D(
        reg_file[1334]), .Y(n32866) );
  AOI22X1 U20160 ( .A(n25565), .B(reg_file[1206]), .C(n25576), .D(
        reg_file[1078]), .Y(n32865) );
  NAND3X1 U20161 ( .A(n32870), .B(n32871), .C(n32872), .Y(n32863) );
  NOR2X1 U20162 ( .A(n32873), .B(n32874), .Y(n32872) );
  OAI22X1 U20163 ( .A(n28246), .B(n25587), .C(n28247), .D(n25597), .Y(n32874)
         );
  OAI22X1 U20164 ( .A(n28248), .B(n25608), .C(n28249), .D(n25618), .Y(n32873)
         );
  AOI22X1 U20165 ( .A(n25629), .B(reg_file[566]), .C(n25640), .D(reg_file[694]), .Y(n32871) );
  AOI22X1 U20166 ( .A(n25651), .B(reg_file[822]), .C(n25662), .D(reg_file[950]), .Y(n32870) );
  NOR2X1 U20167 ( .A(n32875), .B(n32876), .Y(n32861) );
  NAND3X1 U20168 ( .A(n32877), .B(n32878), .C(n32879), .Y(n32876) );
  NOR2X1 U20169 ( .A(n32880), .B(n32881), .Y(n32879) );
  OAI22X1 U20170 ( .A(n28257), .B(n25673), .C(n28258), .D(n25683), .Y(n32881)
         );
  OAI22X1 U20171 ( .A(n28259), .B(n25694), .C(n28260), .D(n25704), .Y(n32880)
         );
  AOI22X1 U20172 ( .A(n25715), .B(reg_file[3510]), .C(n25726), .D(
        reg_file[3382]), .Y(n32878) );
  AOI22X1 U20173 ( .A(n25737), .B(reg_file[3254]), .C(n25748), .D(
        reg_file[3126]), .Y(n32877) );
  NAND3X1 U20174 ( .A(n32882), .B(n32883), .C(n32884), .Y(n32875) );
  NOR2X1 U20175 ( .A(n32885), .B(n32886), .Y(n32884) );
  OAI22X1 U20176 ( .A(n28266), .B(n25759), .C(n28267), .D(n25769), .Y(n32886)
         );
  OAI22X1 U20177 ( .A(n28268), .B(n25780), .C(n28269), .D(n25790), .Y(n32885)
         );
  AOI22X1 U20178 ( .A(n25801), .B(reg_file[2486]), .C(n25812), .D(
        reg_file[2358]), .Y(n32883) );
  AOI22X1 U20179 ( .A(n25823), .B(reg_file[2230]), .C(n25834), .D(
        reg_file[2102]), .Y(n32882) );
  AOI21X1 U20180 ( .A(n32887), .B(n32888), .C(n25490), .Y(rd1data1033_53_) );
  NOR2X1 U20181 ( .A(n32889), .B(n32890), .Y(n32888) );
  NAND3X1 U20182 ( .A(n32891), .B(n32892), .C(n32893), .Y(n32890) );
  NOR2X1 U20183 ( .A(n32894), .B(n32895), .Y(n32893) );
  OAI22X1 U20184 ( .A(n28279), .B(n25501), .C(n28280), .D(n25511), .Y(n32895)
         );
  OAI22X1 U20185 ( .A(n28281), .B(n25522), .C(n28282), .D(n25532), .Y(n32894)
         );
  AOI22X1 U20186 ( .A(n25543), .B(reg_file[1461]), .C(n25554), .D(
        reg_file[1333]), .Y(n32892) );
  AOI22X1 U20187 ( .A(n25565), .B(reg_file[1205]), .C(n25576), .D(
        reg_file[1077]), .Y(n32891) );
  NAND3X1 U20188 ( .A(n32896), .B(n32897), .C(n32898), .Y(n32889) );
  NOR2X1 U20189 ( .A(n32899), .B(n32900), .Y(n32898) );
  OAI22X1 U20190 ( .A(n28288), .B(n25587), .C(n28289), .D(n25597), .Y(n32900)
         );
  OAI22X1 U20191 ( .A(n28290), .B(n25608), .C(n28291), .D(n25618), .Y(n32899)
         );
  AOI22X1 U20192 ( .A(n25629), .B(reg_file[565]), .C(n25640), .D(reg_file[693]), .Y(n32897) );
  AOI22X1 U20193 ( .A(n25651), .B(reg_file[821]), .C(n25662), .D(reg_file[949]), .Y(n32896) );
  NOR2X1 U20194 ( .A(n32901), .B(n32902), .Y(n32887) );
  NAND3X1 U20195 ( .A(n32903), .B(n32904), .C(n32905), .Y(n32902) );
  NOR2X1 U20196 ( .A(n32906), .B(n32907), .Y(n32905) );
  OAI22X1 U20197 ( .A(n28299), .B(n25673), .C(n28300), .D(n25683), .Y(n32907)
         );
  OAI22X1 U20198 ( .A(n28301), .B(n25694), .C(n28302), .D(n25704), .Y(n32906)
         );
  AOI22X1 U20199 ( .A(n25715), .B(reg_file[3509]), .C(n25726), .D(
        reg_file[3381]), .Y(n32904) );
  AOI22X1 U20200 ( .A(n25737), .B(reg_file[3253]), .C(n25748), .D(
        reg_file[3125]), .Y(n32903) );
  NAND3X1 U20201 ( .A(n32908), .B(n32909), .C(n32910), .Y(n32901) );
  NOR2X1 U20202 ( .A(n32911), .B(n32912), .Y(n32910) );
  OAI22X1 U20203 ( .A(n28308), .B(n25759), .C(n28309), .D(n25769), .Y(n32912)
         );
  OAI22X1 U20204 ( .A(n28310), .B(n25780), .C(n28311), .D(n25790), .Y(n32911)
         );
  AOI22X1 U20205 ( .A(n25801), .B(reg_file[2485]), .C(n25812), .D(
        reg_file[2357]), .Y(n32909) );
  AOI22X1 U20206 ( .A(n25823), .B(reg_file[2229]), .C(n25834), .D(
        reg_file[2101]), .Y(n32908) );
  AOI21X1 U20207 ( .A(n32913), .B(n32914), .C(n25490), .Y(rd1data1033_52_) );
  NOR2X1 U20208 ( .A(n32915), .B(n32916), .Y(n32914) );
  NAND3X1 U20209 ( .A(n32917), .B(n32918), .C(n32919), .Y(n32916) );
  NOR2X1 U20210 ( .A(n32920), .B(n32921), .Y(n32919) );
  OAI22X1 U20211 ( .A(n28321), .B(n25501), .C(n28322), .D(n25511), .Y(n32921)
         );
  OAI22X1 U20212 ( .A(n28323), .B(n25522), .C(n28324), .D(n25532), .Y(n32920)
         );
  AOI22X1 U20213 ( .A(n25543), .B(reg_file[1460]), .C(n25554), .D(
        reg_file[1332]), .Y(n32918) );
  AOI22X1 U20214 ( .A(n25565), .B(reg_file[1204]), .C(n25576), .D(
        reg_file[1076]), .Y(n32917) );
  NAND3X1 U20215 ( .A(n32922), .B(n32923), .C(n32924), .Y(n32915) );
  NOR2X1 U20216 ( .A(n32925), .B(n32926), .Y(n32924) );
  OAI22X1 U20217 ( .A(n28330), .B(n25587), .C(n28331), .D(n25597), .Y(n32926)
         );
  OAI22X1 U20218 ( .A(n28332), .B(n25608), .C(n28333), .D(n25618), .Y(n32925)
         );
  AOI22X1 U20219 ( .A(n25629), .B(reg_file[564]), .C(n25640), .D(reg_file[692]), .Y(n32923) );
  AOI22X1 U20220 ( .A(n25651), .B(reg_file[820]), .C(n25662), .D(reg_file[948]), .Y(n32922) );
  NOR2X1 U20221 ( .A(n32927), .B(n32928), .Y(n32913) );
  NAND3X1 U20222 ( .A(n32929), .B(n32930), .C(n32931), .Y(n32928) );
  NOR2X1 U20223 ( .A(n32932), .B(n32933), .Y(n32931) );
  OAI22X1 U20224 ( .A(n28341), .B(n25673), .C(n28342), .D(n25683), .Y(n32933)
         );
  OAI22X1 U20225 ( .A(n28343), .B(n25694), .C(n28344), .D(n25704), .Y(n32932)
         );
  AOI22X1 U20226 ( .A(n25715), .B(reg_file[3508]), .C(n25726), .D(
        reg_file[3380]), .Y(n32930) );
  AOI22X1 U20227 ( .A(n25737), .B(reg_file[3252]), .C(n25748), .D(
        reg_file[3124]), .Y(n32929) );
  NAND3X1 U20228 ( .A(n32934), .B(n32935), .C(n32936), .Y(n32927) );
  NOR2X1 U20229 ( .A(n32937), .B(n32938), .Y(n32936) );
  OAI22X1 U20230 ( .A(n28350), .B(n25759), .C(n28351), .D(n25769), .Y(n32938)
         );
  OAI22X1 U20231 ( .A(n28352), .B(n25780), .C(n28353), .D(n25790), .Y(n32937)
         );
  AOI22X1 U20232 ( .A(n25801), .B(reg_file[2484]), .C(n25812), .D(
        reg_file[2356]), .Y(n32935) );
  AOI22X1 U20233 ( .A(n25823), .B(reg_file[2228]), .C(n25834), .D(
        reg_file[2100]), .Y(n32934) );
  AOI21X1 U20234 ( .A(n32939), .B(n32940), .C(n25490), .Y(rd1data1033_51_) );
  NOR2X1 U20235 ( .A(n32941), .B(n32942), .Y(n32940) );
  NAND3X1 U20236 ( .A(n32943), .B(n32944), .C(n32945), .Y(n32942) );
  NOR2X1 U20237 ( .A(n32946), .B(n32947), .Y(n32945) );
  OAI22X1 U20238 ( .A(n28363), .B(n25501), .C(n28364), .D(n25511), .Y(n32947)
         );
  OAI22X1 U20239 ( .A(n28365), .B(n25522), .C(n28366), .D(n25532), .Y(n32946)
         );
  AOI22X1 U20240 ( .A(n25543), .B(reg_file[1459]), .C(n25554), .D(
        reg_file[1331]), .Y(n32944) );
  AOI22X1 U20241 ( .A(n25565), .B(reg_file[1203]), .C(n25576), .D(
        reg_file[1075]), .Y(n32943) );
  NAND3X1 U20242 ( .A(n32948), .B(n32949), .C(n32950), .Y(n32941) );
  NOR2X1 U20243 ( .A(n32951), .B(n32952), .Y(n32950) );
  OAI22X1 U20244 ( .A(n28372), .B(n25587), .C(n28373), .D(n25597), .Y(n32952)
         );
  OAI22X1 U20245 ( .A(n28374), .B(n25608), .C(n28375), .D(n25618), .Y(n32951)
         );
  AOI22X1 U20246 ( .A(n25629), .B(reg_file[563]), .C(n25640), .D(reg_file[691]), .Y(n32949) );
  AOI22X1 U20247 ( .A(n25651), .B(reg_file[819]), .C(n25662), .D(reg_file[947]), .Y(n32948) );
  NOR2X1 U20248 ( .A(n32953), .B(n32954), .Y(n32939) );
  NAND3X1 U20249 ( .A(n32955), .B(n32956), .C(n32957), .Y(n32954) );
  NOR2X1 U20250 ( .A(n32958), .B(n32959), .Y(n32957) );
  OAI22X1 U20251 ( .A(n28383), .B(n25673), .C(n28384), .D(n25683), .Y(n32959)
         );
  OAI22X1 U20252 ( .A(n28385), .B(n25694), .C(n28386), .D(n25704), .Y(n32958)
         );
  AOI22X1 U20253 ( .A(n25715), .B(reg_file[3507]), .C(n25726), .D(
        reg_file[3379]), .Y(n32956) );
  AOI22X1 U20254 ( .A(n25737), .B(reg_file[3251]), .C(n25748), .D(
        reg_file[3123]), .Y(n32955) );
  NAND3X1 U20255 ( .A(n32960), .B(n32961), .C(n32962), .Y(n32953) );
  NOR2X1 U20256 ( .A(n32963), .B(n32964), .Y(n32962) );
  OAI22X1 U20257 ( .A(n28392), .B(n25759), .C(n28393), .D(n25769), .Y(n32964)
         );
  OAI22X1 U20258 ( .A(n28394), .B(n25780), .C(n28395), .D(n25790), .Y(n32963)
         );
  AOI22X1 U20259 ( .A(n25801), .B(reg_file[2483]), .C(n25812), .D(
        reg_file[2355]), .Y(n32961) );
  AOI22X1 U20260 ( .A(n25823), .B(reg_file[2227]), .C(n25834), .D(
        reg_file[2099]), .Y(n32960) );
  AOI21X1 U20261 ( .A(n32965), .B(n32966), .C(n25490), .Y(rd1data1033_50_) );
  NOR2X1 U20262 ( .A(n32967), .B(n32968), .Y(n32966) );
  NAND3X1 U20263 ( .A(n32969), .B(n32970), .C(n32971), .Y(n32968) );
  NOR2X1 U20264 ( .A(n32972), .B(n32973), .Y(n32971) );
  OAI22X1 U20265 ( .A(n28405), .B(n25501), .C(n28406), .D(n25511), .Y(n32973)
         );
  OAI22X1 U20266 ( .A(n28407), .B(n25522), .C(n28408), .D(n25532), .Y(n32972)
         );
  AOI22X1 U20267 ( .A(n25543), .B(reg_file[1458]), .C(n25554), .D(
        reg_file[1330]), .Y(n32970) );
  AOI22X1 U20268 ( .A(n25565), .B(reg_file[1202]), .C(n25576), .D(
        reg_file[1074]), .Y(n32969) );
  NAND3X1 U20269 ( .A(n32974), .B(n32975), .C(n32976), .Y(n32967) );
  NOR2X1 U20270 ( .A(n32977), .B(n32978), .Y(n32976) );
  OAI22X1 U20271 ( .A(n28414), .B(n25587), .C(n28415), .D(n25597), .Y(n32978)
         );
  OAI22X1 U20272 ( .A(n28416), .B(n25608), .C(n28417), .D(n25618), .Y(n32977)
         );
  AOI22X1 U20273 ( .A(n25629), .B(reg_file[562]), .C(n25640), .D(reg_file[690]), .Y(n32975) );
  AOI22X1 U20274 ( .A(n25651), .B(reg_file[818]), .C(n25662), .D(reg_file[946]), .Y(n32974) );
  NOR2X1 U20275 ( .A(n32979), .B(n32980), .Y(n32965) );
  NAND3X1 U20276 ( .A(n32981), .B(n32982), .C(n32983), .Y(n32980) );
  NOR2X1 U20277 ( .A(n32984), .B(n32985), .Y(n32983) );
  OAI22X1 U20278 ( .A(n28425), .B(n25673), .C(n28426), .D(n25683), .Y(n32985)
         );
  OAI22X1 U20279 ( .A(n28427), .B(n25694), .C(n28428), .D(n25704), .Y(n32984)
         );
  AOI22X1 U20280 ( .A(n25715), .B(reg_file[3506]), .C(n25726), .D(
        reg_file[3378]), .Y(n32982) );
  AOI22X1 U20281 ( .A(n25737), .B(reg_file[3250]), .C(n25748), .D(
        reg_file[3122]), .Y(n32981) );
  NAND3X1 U20282 ( .A(n32986), .B(n32987), .C(n32988), .Y(n32979) );
  NOR2X1 U20283 ( .A(n32989), .B(n32990), .Y(n32988) );
  OAI22X1 U20284 ( .A(n28434), .B(n25759), .C(n28435), .D(n25769), .Y(n32990)
         );
  OAI22X1 U20285 ( .A(n28436), .B(n25780), .C(n28437), .D(n25790), .Y(n32989)
         );
  AOI22X1 U20286 ( .A(n25801), .B(reg_file[2482]), .C(n25812), .D(
        reg_file[2354]), .Y(n32987) );
  AOI22X1 U20287 ( .A(n25823), .B(reg_file[2226]), .C(n25834), .D(
        reg_file[2098]), .Y(n32986) );
  AOI21X1 U20288 ( .A(n32991), .B(n32992), .C(n25490), .Y(rd1data1033_4_) );
  NOR2X1 U20289 ( .A(n32993), .B(n32994), .Y(n32992) );
  NAND3X1 U20290 ( .A(n32995), .B(n32996), .C(n32997), .Y(n32994) );
  NOR2X1 U20291 ( .A(n32998), .B(n32999), .Y(n32997) );
  OAI22X1 U20292 ( .A(n28447), .B(n25501), .C(n28448), .D(n25511), .Y(n32999)
         );
  OAI22X1 U20293 ( .A(n28449), .B(n25522), .C(n28450), .D(n25532), .Y(n32998)
         );
  AOI22X1 U20294 ( .A(n25543), .B(reg_file[1412]), .C(n25554), .D(
        reg_file[1284]), .Y(n32996) );
  AOI22X1 U20295 ( .A(n25565), .B(reg_file[1156]), .C(n25576), .D(
        reg_file[1028]), .Y(n32995) );
  NAND3X1 U20296 ( .A(n33000), .B(n33001), .C(n33002), .Y(n32993) );
  NOR2X1 U20297 ( .A(n33003), .B(n33004), .Y(n33002) );
  OAI22X1 U20298 ( .A(n28456), .B(n25587), .C(n28457), .D(n25597), .Y(n33004)
         );
  OAI22X1 U20299 ( .A(n28458), .B(n25608), .C(n28459), .D(n25618), .Y(n33003)
         );
  AOI22X1 U20300 ( .A(n25629), .B(reg_file[516]), .C(n25640), .D(reg_file[644]), .Y(n33001) );
  AOI22X1 U20301 ( .A(n25651), .B(reg_file[772]), .C(n25662), .D(reg_file[900]), .Y(n33000) );
  NOR2X1 U20302 ( .A(n33005), .B(n33006), .Y(n32991) );
  NAND3X1 U20303 ( .A(n33007), .B(n33008), .C(n33009), .Y(n33006) );
  NOR2X1 U20304 ( .A(n33010), .B(n33011), .Y(n33009) );
  OAI22X1 U20305 ( .A(n28467), .B(n25673), .C(n28468), .D(n25683), .Y(n33011)
         );
  OAI22X1 U20306 ( .A(n28469), .B(n25694), .C(n28470), .D(n25704), .Y(n33010)
         );
  AOI22X1 U20307 ( .A(n25715), .B(reg_file[3460]), .C(n25726), .D(
        reg_file[3332]), .Y(n33008) );
  AOI22X1 U20308 ( .A(n25737), .B(reg_file[3204]), .C(n25748), .D(
        reg_file[3076]), .Y(n33007) );
  NAND3X1 U20309 ( .A(n33012), .B(n33013), .C(n33014), .Y(n33005) );
  NOR2X1 U20310 ( .A(n33015), .B(n33016), .Y(n33014) );
  OAI22X1 U20311 ( .A(n28476), .B(n25759), .C(n28477), .D(n25769), .Y(n33016)
         );
  OAI22X1 U20312 ( .A(n28478), .B(n25780), .C(n28479), .D(n25790), .Y(n33015)
         );
  AOI22X1 U20313 ( .A(n25801), .B(reg_file[2436]), .C(n25812), .D(
        reg_file[2308]), .Y(n33013) );
  AOI22X1 U20314 ( .A(n25823), .B(reg_file[2180]), .C(n25834), .D(
        reg_file[2052]), .Y(n33012) );
  AOI21X1 U20315 ( .A(n33017), .B(n33018), .C(n25489), .Y(rd1data1033_49_) );
  NOR2X1 U20316 ( .A(n33019), .B(n33020), .Y(n33018) );
  NAND3X1 U20317 ( .A(n33021), .B(n33022), .C(n33023), .Y(n33020) );
  NOR2X1 U20318 ( .A(n33024), .B(n33025), .Y(n33023) );
  OAI22X1 U20319 ( .A(n28489), .B(n25500), .C(n28490), .D(n25511), .Y(n33025)
         );
  OAI22X1 U20320 ( .A(n28491), .B(n25521), .C(n28492), .D(n25532), .Y(n33024)
         );
  AOI22X1 U20321 ( .A(n25542), .B(reg_file[1457]), .C(n25553), .D(
        reg_file[1329]), .Y(n33022) );
  AOI22X1 U20322 ( .A(n25564), .B(reg_file[1201]), .C(n25575), .D(
        reg_file[1073]), .Y(n33021) );
  NAND3X1 U20323 ( .A(n33026), .B(n33027), .C(n33028), .Y(n33019) );
  NOR2X1 U20324 ( .A(n33029), .B(n33030), .Y(n33028) );
  OAI22X1 U20325 ( .A(n28498), .B(n25586), .C(n28499), .D(n25597), .Y(n33030)
         );
  OAI22X1 U20326 ( .A(n28500), .B(n25607), .C(n28501), .D(n25618), .Y(n33029)
         );
  AOI22X1 U20327 ( .A(n25628), .B(reg_file[561]), .C(n25639), .D(reg_file[689]), .Y(n33027) );
  AOI22X1 U20328 ( .A(n25650), .B(reg_file[817]), .C(n25661), .D(reg_file[945]), .Y(n33026) );
  NOR2X1 U20329 ( .A(n33031), .B(n33032), .Y(n33017) );
  NAND3X1 U20330 ( .A(n33033), .B(n33034), .C(n33035), .Y(n33032) );
  NOR2X1 U20331 ( .A(n33036), .B(n33037), .Y(n33035) );
  OAI22X1 U20332 ( .A(n28509), .B(n25672), .C(n28510), .D(n25683), .Y(n33037)
         );
  OAI22X1 U20333 ( .A(n28511), .B(n25693), .C(n28512), .D(n25704), .Y(n33036)
         );
  AOI22X1 U20334 ( .A(n25714), .B(reg_file[3505]), .C(n25725), .D(
        reg_file[3377]), .Y(n33034) );
  AOI22X1 U20335 ( .A(n25736), .B(reg_file[3249]), .C(n25747), .D(
        reg_file[3121]), .Y(n33033) );
  NAND3X1 U20336 ( .A(n33038), .B(n33039), .C(n33040), .Y(n33031) );
  NOR2X1 U20337 ( .A(n33041), .B(n33042), .Y(n33040) );
  OAI22X1 U20338 ( .A(n28518), .B(n25758), .C(n28519), .D(n25769), .Y(n33042)
         );
  OAI22X1 U20339 ( .A(n28520), .B(n25779), .C(n28521), .D(n25790), .Y(n33041)
         );
  AOI22X1 U20340 ( .A(n25800), .B(reg_file[2481]), .C(n25811), .D(
        reg_file[2353]), .Y(n33039) );
  AOI22X1 U20341 ( .A(n25822), .B(reg_file[2225]), .C(n25833), .D(
        reg_file[2097]), .Y(n33038) );
  AOI21X1 U20342 ( .A(n33043), .B(n33044), .C(n25489), .Y(rd1data1033_48_) );
  NOR2X1 U20343 ( .A(n33045), .B(n33046), .Y(n33044) );
  NAND3X1 U20344 ( .A(n33047), .B(n33048), .C(n33049), .Y(n33046) );
  NOR2X1 U20345 ( .A(n33050), .B(n33051), .Y(n33049) );
  OAI22X1 U20346 ( .A(n28531), .B(n25500), .C(n28532), .D(n25511), .Y(n33051)
         );
  OAI22X1 U20347 ( .A(n28533), .B(n25521), .C(n28534), .D(n25532), .Y(n33050)
         );
  AOI22X1 U20348 ( .A(n25542), .B(reg_file[1456]), .C(n25553), .D(
        reg_file[1328]), .Y(n33048) );
  AOI22X1 U20349 ( .A(n25564), .B(reg_file[1200]), .C(n25575), .D(
        reg_file[1072]), .Y(n33047) );
  NAND3X1 U20350 ( .A(n33052), .B(n33053), .C(n33054), .Y(n33045) );
  NOR2X1 U20351 ( .A(n33055), .B(n33056), .Y(n33054) );
  OAI22X1 U20352 ( .A(n28540), .B(n25586), .C(n28541), .D(n25597), .Y(n33056)
         );
  OAI22X1 U20353 ( .A(n28542), .B(n25607), .C(n28543), .D(n25618), .Y(n33055)
         );
  AOI22X1 U20354 ( .A(n25628), .B(reg_file[560]), .C(n25639), .D(reg_file[688]), .Y(n33053) );
  AOI22X1 U20355 ( .A(n25650), .B(reg_file[816]), .C(n25661), .D(reg_file[944]), .Y(n33052) );
  NOR2X1 U20356 ( .A(n33057), .B(n33058), .Y(n33043) );
  NAND3X1 U20357 ( .A(n33059), .B(n33060), .C(n33061), .Y(n33058) );
  NOR2X1 U20358 ( .A(n33062), .B(n33063), .Y(n33061) );
  OAI22X1 U20359 ( .A(n28551), .B(n25672), .C(n28552), .D(n25683), .Y(n33063)
         );
  OAI22X1 U20360 ( .A(n28553), .B(n25693), .C(n28554), .D(n25704), .Y(n33062)
         );
  AOI22X1 U20361 ( .A(n25714), .B(reg_file[3504]), .C(n25725), .D(
        reg_file[3376]), .Y(n33060) );
  AOI22X1 U20362 ( .A(n25736), .B(reg_file[3248]), .C(n25747), .D(
        reg_file[3120]), .Y(n33059) );
  NAND3X1 U20363 ( .A(n33064), .B(n33065), .C(n33066), .Y(n33057) );
  NOR2X1 U20364 ( .A(n33067), .B(n33068), .Y(n33066) );
  OAI22X1 U20365 ( .A(n28560), .B(n25758), .C(n28561), .D(n25769), .Y(n33068)
         );
  OAI22X1 U20366 ( .A(n28562), .B(n25779), .C(n28563), .D(n25790), .Y(n33067)
         );
  AOI22X1 U20367 ( .A(n25800), .B(reg_file[2480]), .C(n25811), .D(
        reg_file[2352]), .Y(n33065) );
  AOI22X1 U20368 ( .A(n25822), .B(reg_file[2224]), .C(n25833), .D(
        reg_file[2096]), .Y(n33064) );
  AOI21X1 U20369 ( .A(n33069), .B(n33070), .C(n25489), .Y(rd1data1033_47_) );
  NOR2X1 U20370 ( .A(n33071), .B(n33072), .Y(n33070) );
  NAND3X1 U20371 ( .A(n33073), .B(n33074), .C(n33075), .Y(n33072) );
  NOR2X1 U20372 ( .A(n33076), .B(n33077), .Y(n33075) );
  OAI22X1 U20373 ( .A(n28573), .B(n25500), .C(n28574), .D(n25511), .Y(n33077)
         );
  OAI22X1 U20374 ( .A(n28575), .B(n25521), .C(n28576), .D(n25532), .Y(n33076)
         );
  AOI22X1 U20375 ( .A(n25542), .B(reg_file[1455]), .C(n25553), .D(
        reg_file[1327]), .Y(n33074) );
  AOI22X1 U20376 ( .A(n25564), .B(reg_file[1199]), .C(n25575), .D(
        reg_file[1071]), .Y(n33073) );
  NAND3X1 U20377 ( .A(n33078), .B(n33079), .C(n33080), .Y(n33071) );
  NOR2X1 U20378 ( .A(n33081), .B(n33082), .Y(n33080) );
  OAI22X1 U20379 ( .A(n28582), .B(n25586), .C(n28583), .D(n25597), .Y(n33082)
         );
  OAI22X1 U20380 ( .A(n28584), .B(n25607), .C(n28585), .D(n25618), .Y(n33081)
         );
  AOI22X1 U20381 ( .A(n25628), .B(reg_file[559]), .C(n25639), .D(reg_file[687]), .Y(n33079) );
  AOI22X1 U20382 ( .A(n25650), .B(reg_file[815]), .C(n25661), .D(reg_file[943]), .Y(n33078) );
  NOR2X1 U20383 ( .A(n33083), .B(n33084), .Y(n33069) );
  NAND3X1 U20384 ( .A(n33085), .B(n33086), .C(n33087), .Y(n33084) );
  NOR2X1 U20385 ( .A(n33088), .B(n33089), .Y(n33087) );
  OAI22X1 U20386 ( .A(n28593), .B(n25672), .C(n28594), .D(n25683), .Y(n33089)
         );
  OAI22X1 U20387 ( .A(n28595), .B(n25693), .C(n28596), .D(n25704), .Y(n33088)
         );
  AOI22X1 U20388 ( .A(n25714), .B(reg_file[3503]), .C(n25725), .D(
        reg_file[3375]), .Y(n33086) );
  AOI22X1 U20389 ( .A(n25736), .B(reg_file[3247]), .C(n25747), .D(
        reg_file[3119]), .Y(n33085) );
  NAND3X1 U20390 ( .A(n33090), .B(n33091), .C(n33092), .Y(n33083) );
  NOR2X1 U20391 ( .A(n33093), .B(n33094), .Y(n33092) );
  OAI22X1 U20392 ( .A(n28602), .B(n25758), .C(n28603), .D(n25769), .Y(n33094)
         );
  OAI22X1 U20393 ( .A(n28604), .B(n25779), .C(n28605), .D(n25790), .Y(n33093)
         );
  AOI22X1 U20394 ( .A(n25800), .B(reg_file[2479]), .C(n25811), .D(
        reg_file[2351]), .Y(n33091) );
  AOI22X1 U20395 ( .A(n25822), .B(reg_file[2223]), .C(n25833), .D(
        reg_file[2095]), .Y(n33090) );
  AOI21X1 U20396 ( .A(n33095), .B(n33096), .C(n25489), .Y(rd1data1033_46_) );
  NOR2X1 U20397 ( .A(n33097), .B(n33098), .Y(n33096) );
  NAND3X1 U20398 ( .A(n33099), .B(n33100), .C(n33101), .Y(n33098) );
  NOR2X1 U20399 ( .A(n33102), .B(n33103), .Y(n33101) );
  OAI22X1 U20400 ( .A(n28615), .B(n25500), .C(n28616), .D(n25511), .Y(n33103)
         );
  OAI22X1 U20401 ( .A(n28617), .B(n25521), .C(n28618), .D(n25532), .Y(n33102)
         );
  AOI22X1 U20402 ( .A(n25542), .B(reg_file[1454]), .C(n25553), .D(
        reg_file[1326]), .Y(n33100) );
  AOI22X1 U20403 ( .A(n25564), .B(reg_file[1198]), .C(n25575), .D(
        reg_file[1070]), .Y(n33099) );
  NAND3X1 U20404 ( .A(n33104), .B(n33105), .C(n33106), .Y(n33097) );
  NOR2X1 U20405 ( .A(n33107), .B(n33108), .Y(n33106) );
  OAI22X1 U20406 ( .A(n28624), .B(n25586), .C(n28625), .D(n25597), .Y(n33108)
         );
  OAI22X1 U20407 ( .A(n28626), .B(n25607), .C(n28627), .D(n25618), .Y(n33107)
         );
  AOI22X1 U20408 ( .A(n25628), .B(reg_file[558]), .C(n25639), .D(reg_file[686]), .Y(n33105) );
  AOI22X1 U20409 ( .A(n25650), .B(reg_file[814]), .C(n25661), .D(reg_file[942]), .Y(n33104) );
  NOR2X1 U20410 ( .A(n33109), .B(n33110), .Y(n33095) );
  NAND3X1 U20411 ( .A(n33111), .B(n33112), .C(n33113), .Y(n33110) );
  NOR2X1 U20412 ( .A(n33114), .B(n33115), .Y(n33113) );
  OAI22X1 U20413 ( .A(n28635), .B(n25672), .C(n28636), .D(n25683), .Y(n33115)
         );
  OAI22X1 U20414 ( .A(n28637), .B(n25693), .C(n28638), .D(n25704), .Y(n33114)
         );
  AOI22X1 U20415 ( .A(n25714), .B(reg_file[3502]), .C(n25725), .D(
        reg_file[3374]), .Y(n33112) );
  AOI22X1 U20416 ( .A(n25736), .B(reg_file[3246]), .C(n25747), .D(
        reg_file[3118]), .Y(n33111) );
  NAND3X1 U20417 ( .A(n33116), .B(n33117), .C(n33118), .Y(n33109) );
  NOR2X1 U20418 ( .A(n33119), .B(n33120), .Y(n33118) );
  OAI22X1 U20419 ( .A(n28644), .B(n25758), .C(n28645), .D(n25769), .Y(n33120)
         );
  OAI22X1 U20420 ( .A(n28646), .B(n25779), .C(n28647), .D(n25790), .Y(n33119)
         );
  AOI22X1 U20421 ( .A(n25800), .B(reg_file[2478]), .C(n25811), .D(
        reg_file[2350]), .Y(n33117) );
  AOI22X1 U20422 ( .A(n25822), .B(reg_file[2222]), .C(n25833), .D(
        reg_file[2094]), .Y(n33116) );
  AOI21X1 U20423 ( .A(n33121), .B(n33122), .C(n25489), .Y(rd1data1033_45_) );
  NOR2X1 U20424 ( .A(n33123), .B(n33124), .Y(n33122) );
  NAND3X1 U20425 ( .A(n33125), .B(n33126), .C(n33127), .Y(n33124) );
  NOR2X1 U20426 ( .A(n33128), .B(n33129), .Y(n33127) );
  OAI22X1 U20427 ( .A(n28657), .B(n25500), .C(n28658), .D(n25511), .Y(n33129)
         );
  OAI22X1 U20428 ( .A(n28659), .B(n25521), .C(n28660), .D(n25532), .Y(n33128)
         );
  AOI22X1 U20429 ( .A(n25542), .B(reg_file[1453]), .C(n25553), .D(
        reg_file[1325]), .Y(n33126) );
  AOI22X1 U20430 ( .A(n25564), .B(reg_file[1197]), .C(n25575), .D(
        reg_file[1069]), .Y(n33125) );
  NAND3X1 U20431 ( .A(n33130), .B(n33131), .C(n33132), .Y(n33123) );
  NOR2X1 U20432 ( .A(n33133), .B(n33134), .Y(n33132) );
  OAI22X1 U20433 ( .A(n28666), .B(n25586), .C(n28667), .D(n25597), .Y(n33134)
         );
  OAI22X1 U20434 ( .A(n28668), .B(n25607), .C(n28669), .D(n25618), .Y(n33133)
         );
  AOI22X1 U20435 ( .A(n25628), .B(reg_file[557]), .C(n25639), .D(reg_file[685]), .Y(n33131) );
  AOI22X1 U20436 ( .A(n25650), .B(reg_file[813]), .C(n25661), .D(reg_file[941]), .Y(n33130) );
  NOR2X1 U20437 ( .A(n33135), .B(n33136), .Y(n33121) );
  NAND3X1 U20438 ( .A(n33137), .B(n33138), .C(n33139), .Y(n33136) );
  NOR2X1 U20439 ( .A(n33140), .B(n33141), .Y(n33139) );
  OAI22X1 U20440 ( .A(n28677), .B(n25672), .C(n28678), .D(n25683), .Y(n33141)
         );
  OAI22X1 U20441 ( .A(n28679), .B(n25693), .C(n28680), .D(n25704), .Y(n33140)
         );
  AOI22X1 U20442 ( .A(n25714), .B(reg_file[3501]), .C(n25725), .D(
        reg_file[3373]), .Y(n33138) );
  AOI22X1 U20443 ( .A(n25736), .B(reg_file[3245]), .C(n25747), .D(
        reg_file[3117]), .Y(n33137) );
  NAND3X1 U20444 ( .A(n33142), .B(n33143), .C(n33144), .Y(n33135) );
  NOR2X1 U20445 ( .A(n33145), .B(n33146), .Y(n33144) );
  OAI22X1 U20446 ( .A(n28686), .B(n25758), .C(n28687), .D(n25769), .Y(n33146)
         );
  OAI22X1 U20447 ( .A(n28688), .B(n25779), .C(n28689), .D(n25790), .Y(n33145)
         );
  AOI22X1 U20448 ( .A(n25800), .B(reg_file[2477]), .C(n25811), .D(
        reg_file[2349]), .Y(n33143) );
  AOI22X1 U20449 ( .A(n25822), .B(reg_file[2221]), .C(n25833), .D(
        reg_file[2093]), .Y(n33142) );
  AOI21X1 U20450 ( .A(n33147), .B(n33148), .C(n25489), .Y(rd1data1033_44_) );
  NOR2X1 U20451 ( .A(n33149), .B(n33150), .Y(n33148) );
  NAND3X1 U20452 ( .A(n33151), .B(n33152), .C(n33153), .Y(n33150) );
  NOR2X1 U20453 ( .A(n33154), .B(n33155), .Y(n33153) );
  OAI22X1 U20454 ( .A(n28699), .B(n25500), .C(n28700), .D(n25511), .Y(n33155)
         );
  OAI22X1 U20455 ( .A(n28701), .B(n25521), .C(n28702), .D(n25532), .Y(n33154)
         );
  AOI22X1 U20456 ( .A(n25542), .B(reg_file[1452]), .C(n25553), .D(
        reg_file[1324]), .Y(n33152) );
  AOI22X1 U20457 ( .A(n25564), .B(reg_file[1196]), .C(n25575), .D(
        reg_file[1068]), .Y(n33151) );
  NAND3X1 U20458 ( .A(n33156), .B(n33157), .C(n33158), .Y(n33149) );
  NOR2X1 U20459 ( .A(n33159), .B(n33160), .Y(n33158) );
  OAI22X1 U20460 ( .A(n28708), .B(n25586), .C(n28709), .D(n25597), .Y(n33160)
         );
  OAI22X1 U20461 ( .A(n28710), .B(n25607), .C(n28711), .D(n25618), .Y(n33159)
         );
  AOI22X1 U20462 ( .A(n25628), .B(reg_file[556]), .C(n25639), .D(reg_file[684]), .Y(n33157) );
  AOI22X1 U20463 ( .A(n25650), .B(reg_file[812]), .C(n25661), .D(reg_file[940]), .Y(n33156) );
  NOR2X1 U20464 ( .A(n33161), .B(n33162), .Y(n33147) );
  NAND3X1 U20465 ( .A(n33163), .B(n33164), .C(n33165), .Y(n33162) );
  NOR2X1 U20466 ( .A(n33166), .B(n33167), .Y(n33165) );
  OAI22X1 U20467 ( .A(n28719), .B(n25672), .C(n28720), .D(n25683), .Y(n33167)
         );
  OAI22X1 U20468 ( .A(n28721), .B(n25693), .C(n28722), .D(n25704), .Y(n33166)
         );
  AOI22X1 U20469 ( .A(n25714), .B(reg_file[3500]), .C(n25725), .D(
        reg_file[3372]), .Y(n33164) );
  AOI22X1 U20470 ( .A(n25736), .B(reg_file[3244]), .C(n25747), .D(
        reg_file[3116]), .Y(n33163) );
  NAND3X1 U20471 ( .A(n33168), .B(n33169), .C(n33170), .Y(n33161) );
  NOR2X1 U20472 ( .A(n33171), .B(n33172), .Y(n33170) );
  OAI22X1 U20473 ( .A(n28728), .B(n25758), .C(n28729), .D(n25769), .Y(n33172)
         );
  OAI22X1 U20474 ( .A(n28730), .B(n25779), .C(n28731), .D(n25790), .Y(n33171)
         );
  AOI22X1 U20475 ( .A(n25800), .B(reg_file[2476]), .C(n25811), .D(
        reg_file[2348]), .Y(n33169) );
  AOI22X1 U20476 ( .A(n25822), .B(reg_file[2220]), .C(n25833), .D(
        reg_file[2092]), .Y(n33168) );
  AOI21X1 U20477 ( .A(n33173), .B(n33174), .C(n25489), .Y(rd1data1033_43_) );
  NOR2X1 U20478 ( .A(n33175), .B(n33176), .Y(n33174) );
  NAND3X1 U20479 ( .A(n33177), .B(n33178), .C(n33179), .Y(n33176) );
  NOR2X1 U20480 ( .A(n33180), .B(n33181), .Y(n33179) );
  OAI22X1 U20481 ( .A(n28741), .B(n25500), .C(n28742), .D(n25511), .Y(n33181)
         );
  OAI22X1 U20482 ( .A(n28743), .B(n25521), .C(n28744), .D(n25532), .Y(n33180)
         );
  AOI22X1 U20483 ( .A(n25542), .B(reg_file[1451]), .C(n25553), .D(
        reg_file[1323]), .Y(n33178) );
  AOI22X1 U20484 ( .A(n25564), .B(reg_file[1195]), .C(n25575), .D(
        reg_file[1067]), .Y(n33177) );
  NAND3X1 U20485 ( .A(n33182), .B(n33183), .C(n33184), .Y(n33175) );
  NOR2X1 U20486 ( .A(n33185), .B(n33186), .Y(n33184) );
  OAI22X1 U20487 ( .A(n28750), .B(n25586), .C(n28751), .D(n25597), .Y(n33186)
         );
  OAI22X1 U20488 ( .A(n28752), .B(n25607), .C(n28753), .D(n25618), .Y(n33185)
         );
  AOI22X1 U20489 ( .A(n25628), .B(reg_file[555]), .C(n25639), .D(reg_file[683]), .Y(n33183) );
  AOI22X1 U20490 ( .A(n25650), .B(reg_file[811]), .C(n25661), .D(reg_file[939]), .Y(n33182) );
  NOR2X1 U20491 ( .A(n33187), .B(n33188), .Y(n33173) );
  NAND3X1 U20492 ( .A(n33189), .B(n33190), .C(n33191), .Y(n33188) );
  NOR2X1 U20493 ( .A(n33192), .B(n33193), .Y(n33191) );
  OAI22X1 U20494 ( .A(n28761), .B(n25672), .C(n28762), .D(n25683), .Y(n33193)
         );
  OAI22X1 U20495 ( .A(n28763), .B(n25693), .C(n28764), .D(n25704), .Y(n33192)
         );
  AOI22X1 U20496 ( .A(n25714), .B(reg_file[3499]), .C(n25725), .D(
        reg_file[3371]), .Y(n33190) );
  AOI22X1 U20497 ( .A(n25736), .B(reg_file[3243]), .C(n25747), .D(
        reg_file[3115]), .Y(n33189) );
  NAND3X1 U20498 ( .A(n33194), .B(n33195), .C(n33196), .Y(n33187) );
  NOR2X1 U20499 ( .A(n33197), .B(n33198), .Y(n33196) );
  OAI22X1 U20500 ( .A(n28770), .B(n25758), .C(n28771), .D(n25769), .Y(n33198)
         );
  OAI22X1 U20501 ( .A(n28772), .B(n25779), .C(n28773), .D(n25790), .Y(n33197)
         );
  AOI22X1 U20502 ( .A(n25800), .B(reg_file[2475]), .C(n25811), .D(
        reg_file[2347]), .Y(n33195) );
  AOI22X1 U20503 ( .A(n25822), .B(reg_file[2219]), .C(n25833), .D(
        reg_file[2091]), .Y(n33194) );
  AOI21X1 U20504 ( .A(n33199), .B(n33200), .C(n25489), .Y(rd1data1033_42_) );
  NOR2X1 U20505 ( .A(n33201), .B(n33202), .Y(n33200) );
  NAND3X1 U20506 ( .A(n33203), .B(n33204), .C(n33205), .Y(n33202) );
  NOR2X1 U20507 ( .A(n33206), .B(n33207), .Y(n33205) );
  OAI22X1 U20508 ( .A(n28783), .B(n25500), .C(n28784), .D(n25510), .Y(n33207)
         );
  OAI22X1 U20509 ( .A(n28785), .B(n25521), .C(n28786), .D(n25531), .Y(n33206)
         );
  AOI22X1 U20510 ( .A(n25542), .B(reg_file[1450]), .C(n25553), .D(
        reg_file[1322]), .Y(n33204) );
  AOI22X1 U20511 ( .A(n25564), .B(reg_file[1194]), .C(n25575), .D(
        reg_file[1066]), .Y(n33203) );
  NAND3X1 U20512 ( .A(n33208), .B(n33209), .C(n33210), .Y(n33201) );
  NOR2X1 U20513 ( .A(n33211), .B(n33212), .Y(n33210) );
  OAI22X1 U20514 ( .A(n28792), .B(n25586), .C(n28793), .D(n25596), .Y(n33212)
         );
  OAI22X1 U20515 ( .A(n28794), .B(n25607), .C(n28795), .D(n25617), .Y(n33211)
         );
  AOI22X1 U20516 ( .A(n25628), .B(reg_file[554]), .C(n25639), .D(reg_file[682]), .Y(n33209) );
  AOI22X1 U20517 ( .A(n25650), .B(reg_file[810]), .C(n25661), .D(reg_file[938]), .Y(n33208) );
  NOR2X1 U20518 ( .A(n33213), .B(n33214), .Y(n33199) );
  NAND3X1 U20519 ( .A(n33215), .B(n33216), .C(n33217), .Y(n33214) );
  NOR2X1 U20520 ( .A(n33218), .B(n33219), .Y(n33217) );
  OAI22X1 U20521 ( .A(n28803), .B(n25672), .C(n28804), .D(n25682), .Y(n33219)
         );
  OAI22X1 U20522 ( .A(n28805), .B(n25693), .C(n28806), .D(n25703), .Y(n33218)
         );
  AOI22X1 U20523 ( .A(n25714), .B(reg_file[3498]), .C(n25725), .D(
        reg_file[3370]), .Y(n33216) );
  AOI22X1 U20524 ( .A(n25736), .B(reg_file[3242]), .C(n25747), .D(
        reg_file[3114]), .Y(n33215) );
  NAND3X1 U20525 ( .A(n33220), .B(n33221), .C(n33222), .Y(n33213) );
  NOR2X1 U20526 ( .A(n33223), .B(n33224), .Y(n33222) );
  OAI22X1 U20527 ( .A(n28812), .B(n25758), .C(n28813), .D(n25768), .Y(n33224)
         );
  OAI22X1 U20528 ( .A(n28814), .B(n25779), .C(n28815), .D(n25789), .Y(n33223)
         );
  AOI22X1 U20529 ( .A(n25800), .B(reg_file[2474]), .C(n25811), .D(
        reg_file[2346]), .Y(n33221) );
  AOI22X1 U20530 ( .A(n25822), .B(reg_file[2218]), .C(n25833), .D(
        reg_file[2090]), .Y(n33220) );
  AOI21X1 U20531 ( .A(n33225), .B(n33226), .C(n25489), .Y(rd1data1033_41_) );
  NOR2X1 U20532 ( .A(n33227), .B(n33228), .Y(n33226) );
  NAND3X1 U20533 ( .A(n33229), .B(n33230), .C(n33231), .Y(n33228) );
  NOR2X1 U20534 ( .A(n33232), .B(n33233), .Y(n33231) );
  OAI22X1 U20535 ( .A(n28825), .B(n25500), .C(n28826), .D(n25510), .Y(n33233)
         );
  OAI22X1 U20536 ( .A(n28827), .B(n25521), .C(n28828), .D(n25531), .Y(n33232)
         );
  AOI22X1 U20537 ( .A(n25542), .B(reg_file[1449]), .C(n25553), .D(
        reg_file[1321]), .Y(n33230) );
  AOI22X1 U20538 ( .A(n25564), .B(reg_file[1193]), .C(n25575), .D(
        reg_file[1065]), .Y(n33229) );
  NAND3X1 U20539 ( .A(n33234), .B(n33235), .C(n33236), .Y(n33227) );
  NOR2X1 U20540 ( .A(n33237), .B(n33238), .Y(n33236) );
  OAI22X1 U20541 ( .A(n28834), .B(n25586), .C(n28835), .D(n25596), .Y(n33238)
         );
  OAI22X1 U20542 ( .A(n28836), .B(n25607), .C(n28837), .D(n25617), .Y(n33237)
         );
  AOI22X1 U20543 ( .A(n25628), .B(reg_file[553]), .C(n25639), .D(reg_file[681]), .Y(n33235) );
  AOI22X1 U20544 ( .A(n25650), .B(reg_file[809]), .C(n25661), .D(reg_file[937]), .Y(n33234) );
  NOR2X1 U20545 ( .A(n33239), .B(n33240), .Y(n33225) );
  NAND3X1 U20546 ( .A(n33241), .B(n33242), .C(n33243), .Y(n33240) );
  NOR2X1 U20547 ( .A(n33244), .B(n33245), .Y(n33243) );
  OAI22X1 U20548 ( .A(n28845), .B(n25672), .C(n28846), .D(n25682), .Y(n33245)
         );
  OAI22X1 U20549 ( .A(n28847), .B(n25693), .C(n28848), .D(n25703), .Y(n33244)
         );
  AOI22X1 U20550 ( .A(n25714), .B(reg_file[3497]), .C(n25725), .D(
        reg_file[3369]), .Y(n33242) );
  AOI22X1 U20551 ( .A(n25736), .B(reg_file[3241]), .C(n25747), .D(
        reg_file[3113]), .Y(n33241) );
  NAND3X1 U20552 ( .A(n33246), .B(n33247), .C(n33248), .Y(n33239) );
  NOR2X1 U20553 ( .A(n33249), .B(n33250), .Y(n33248) );
  OAI22X1 U20554 ( .A(n28854), .B(n25758), .C(n28855), .D(n25768), .Y(n33250)
         );
  OAI22X1 U20555 ( .A(n28856), .B(n25779), .C(n28857), .D(n25789), .Y(n33249)
         );
  AOI22X1 U20556 ( .A(n25800), .B(reg_file[2473]), .C(n25811), .D(
        reg_file[2345]), .Y(n33247) );
  AOI22X1 U20557 ( .A(n25822), .B(reg_file[2217]), .C(n25833), .D(
        reg_file[2089]), .Y(n33246) );
  AOI21X1 U20558 ( .A(n33251), .B(n33252), .C(n25489), .Y(rd1data1033_40_) );
  NOR2X1 U20559 ( .A(n33253), .B(n33254), .Y(n33252) );
  NAND3X1 U20560 ( .A(n33255), .B(n33256), .C(n33257), .Y(n33254) );
  NOR2X1 U20561 ( .A(n33258), .B(n33259), .Y(n33257) );
  OAI22X1 U20562 ( .A(n28867), .B(n25500), .C(n28868), .D(n25510), .Y(n33259)
         );
  OAI22X1 U20563 ( .A(n28869), .B(n25521), .C(n28870), .D(n25531), .Y(n33258)
         );
  AOI22X1 U20564 ( .A(n25542), .B(reg_file[1448]), .C(n25553), .D(
        reg_file[1320]), .Y(n33256) );
  AOI22X1 U20565 ( .A(n25564), .B(reg_file[1192]), .C(n25575), .D(
        reg_file[1064]), .Y(n33255) );
  NAND3X1 U20566 ( .A(n33260), .B(n33261), .C(n33262), .Y(n33253) );
  NOR2X1 U20567 ( .A(n33263), .B(n33264), .Y(n33262) );
  OAI22X1 U20568 ( .A(n28876), .B(n25586), .C(n28877), .D(n25596), .Y(n33264)
         );
  OAI22X1 U20569 ( .A(n28878), .B(n25607), .C(n28879), .D(n25617), .Y(n33263)
         );
  AOI22X1 U20570 ( .A(n25628), .B(reg_file[552]), .C(n25639), .D(reg_file[680]), .Y(n33261) );
  AOI22X1 U20571 ( .A(n25650), .B(reg_file[808]), .C(n25661), .D(reg_file[936]), .Y(n33260) );
  NOR2X1 U20572 ( .A(n33265), .B(n33266), .Y(n33251) );
  NAND3X1 U20573 ( .A(n33267), .B(n33268), .C(n33269), .Y(n33266) );
  NOR2X1 U20574 ( .A(n33270), .B(n33271), .Y(n33269) );
  OAI22X1 U20575 ( .A(n28887), .B(n25672), .C(n28888), .D(n25682), .Y(n33271)
         );
  OAI22X1 U20576 ( .A(n28889), .B(n25693), .C(n28890), .D(n25703), .Y(n33270)
         );
  AOI22X1 U20577 ( .A(n25714), .B(reg_file[3496]), .C(n25725), .D(
        reg_file[3368]), .Y(n33268) );
  AOI22X1 U20578 ( .A(n25736), .B(reg_file[3240]), .C(n25747), .D(
        reg_file[3112]), .Y(n33267) );
  NAND3X1 U20579 ( .A(n33272), .B(n33273), .C(n33274), .Y(n33265) );
  NOR2X1 U20580 ( .A(n33275), .B(n33276), .Y(n33274) );
  OAI22X1 U20581 ( .A(n28896), .B(n25758), .C(n28897), .D(n25768), .Y(n33276)
         );
  OAI22X1 U20582 ( .A(n28898), .B(n25779), .C(n28899), .D(n25789), .Y(n33275)
         );
  AOI22X1 U20583 ( .A(n25800), .B(reg_file[2472]), .C(n25811), .D(
        reg_file[2344]), .Y(n33273) );
  AOI22X1 U20584 ( .A(n25822), .B(reg_file[2216]), .C(n25833), .D(
        reg_file[2088]), .Y(n33272) );
  AOI21X1 U20585 ( .A(n33277), .B(n33278), .C(n25489), .Y(rd1data1033_3_) );
  NOR2X1 U20586 ( .A(n33279), .B(n33280), .Y(n33278) );
  NAND3X1 U20587 ( .A(n33281), .B(n33282), .C(n33283), .Y(n33280) );
  NOR2X1 U20588 ( .A(n33284), .B(n33285), .Y(n33283) );
  OAI22X1 U20589 ( .A(n28909), .B(n25500), .C(n28910), .D(n25510), .Y(n33285)
         );
  OAI22X1 U20590 ( .A(n28911), .B(n25521), .C(n28912), .D(n25531), .Y(n33284)
         );
  AOI22X1 U20591 ( .A(n25542), .B(reg_file[1411]), .C(n25553), .D(
        reg_file[1283]), .Y(n33282) );
  AOI22X1 U20592 ( .A(n25564), .B(reg_file[1155]), .C(n25575), .D(
        reg_file[1027]), .Y(n33281) );
  NAND3X1 U20593 ( .A(n33286), .B(n33287), .C(n33288), .Y(n33279) );
  NOR2X1 U20594 ( .A(n33289), .B(n33290), .Y(n33288) );
  OAI22X1 U20595 ( .A(n28918), .B(n25586), .C(n28919), .D(n25596), .Y(n33290)
         );
  OAI22X1 U20596 ( .A(n28920), .B(n25607), .C(n28921), .D(n25617), .Y(n33289)
         );
  AOI22X1 U20597 ( .A(n25628), .B(reg_file[515]), .C(n25639), .D(reg_file[643]), .Y(n33287) );
  AOI22X1 U20598 ( .A(n25650), .B(reg_file[771]), .C(n25661), .D(reg_file[899]), .Y(n33286) );
  NOR2X1 U20599 ( .A(n33291), .B(n33292), .Y(n33277) );
  NAND3X1 U20600 ( .A(n33293), .B(n33294), .C(n33295), .Y(n33292) );
  NOR2X1 U20601 ( .A(n33296), .B(n33297), .Y(n33295) );
  OAI22X1 U20602 ( .A(n28929), .B(n25672), .C(n28930), .D(n25682), .Y(n33297)
         );
  OAI22X1 U20603 ( .A(n28931), .B(n25693), .C(n28932), .D(n25703), .Y(n33296)
         );
  AOI22X1 U20604 ( .A(n25714), .B(reg_file[3459]), .C(n25725), .D(
        reg_file[3331]), .Y(n33294) );
  AOI22X1 U20605 ( .A(n25736), .B(reg_file[3203]), .C(n25747), .D(
        reg_file[3075]), .Y(n33293) );
  NAND3X1 U20606 ( .A(n33298), .B(n33299), .C(n33300), .Y(n33291) );
  NOR2X1 U20607 ( .A(n33301), .B(n33302), .Y(n33300) );
  OAI22X1 U20608 ( .A(n28938), .B(n25758), .C(n28939), .D(n25768), .Y(n33302)
         );
  OAI22X1 U20609 ( .A(n28940), .B(n25779), .C(n28941), .D(n25789), .Y(n33301)
         );
  AOI22X1 U20610 ( .A(n25800), .B(reg_file[2435]), .C(n25811), .D(
        reg_file[2307]), .Y(n33299) );
  AOI22X1 U20611 ( .A(n25822), .B(reg_file[2179]), .C(n25833), .D(
        reg_file[2051]), .Y(n33298) );
  AOI21X1 U20612 ( .A(n33303), .B(n33304), .C(n25489), .Y(rd1data1033_39_) );
  NOR2X1 U20613 ( .A(n33305), .B(n33306), .Y(n33304) );
  NAND3X1 U20614 ( .A(n33307), .B(n33308), .C(n33309), .Y(n33306) );
  NOR2X1 U20615 ( .A(n33310), .B(n33311), .Y(n33309) );
  OAI22X1 U20616 ( .A(n28951), .B(n25500), .C(n28952), .D(n25510), .Y(n33311)
         );
  OAI22X1 U20617 ( .A(n28953), .B(n25521), .C(n28954), .D(n25531), .Y(n33310)
         );
  AOI22X1 U20618 ( .A(n25542), .B(reg_file[1447]), .C(n25553), .D(
        reg_file[1319]), .Y(n33308) );
  AOI22X1 U20619 ( .A(n25564), .B(reg_file[1191]), .C(n25575), .D(
        reg_file[1063]), .Y(n33307) );
  NAND3X1 U20620 ( .A(n33312), .B(n33313), .C(n33314), .Y(n33305) );
  NOR2X1 U20621 ( .A(n33315), .B(n33316), .Y(n33314) );
  OAI22X1 U20622 ( .A(n28960), .B(n25586), .C(n28961), .D(n25596), .Y(n33316)
         );
  OAI22X1 U20623 ( .A(n28962), .B(n25607), .C(n28963), .D(n25617), .Y(n33315)
         );
  AOI22X1 U20624 ( .A(n25628), .B(reg_file[551]), .C(n25639), .D(reg_file[679]), .Y(n33313) );
  AOI22X1 U20625 ( .A(n25650), .B(reg_file[807]), .C(n25661), .D(reg_file[935]), .Y(n33312) );
  NOR2X1 U20626 ( .A(n33317), .B(n33318), .Y(n33303) );
  NAND3X1 U20627 ( .A(n33319), .B(n33320), .C(n33321), .Y(n33318) );
  NOR2X1 U20628 ( .A(n33322), .B(n33323), .Y(n33321) );
  OAI22X1 U20629 ( .A(n28971), .B(n25672), .C(n28972), .D(n25682), .Y(n33323)
         );
  OAI22X1 U20630 ( .A(n28973), .B(n25693), .C(n28974), .D(n25703), .Y(n33322)
         );
  AOI22X1 U20631 ( .A(n25714), .B(reg_file[3495]), .C(n25725), .D(
        reg_file[3367]), .Y(n33320) );
  AOI22X1 U20632 ( .A(n25736), .B(reg_file[3239]), .C(n25747), .D(
        reg_file[3111]), .Y(n33319) );
  NAND3X1 U20633 ( .A(n33324), .B(n33325), .C(n33326), .Y(n33317) );
  NOR2X1 U20634 ( .A(n33327), .B(n33328), .Y(n33326) );
  OAI22X1 U20635 ( .A(n28980), .B(n25758), .C(n28981), .D(n25768), .Y(n33328)
         );
  OAI22X1 U20636 ( .A(n28982), .B(n25779), .C(n28983), .D(n25789), .Y(n33327)
         );
  AOI22X1 U20637 ( .A(n25800), .B(reg_file[2471]), .C(n25811), .D(
        reg_file[2343]), .Y(n33325) );
  AOI22X1 U20638 ( .A(n25822), .B(reg_file[2215]), .C(n25833), .D(
        reg_file[2087]), .Y(n33324) );
  AOI21X1 U20639 ( .A(n33329), .B(n33330), .C(n25488), .Y(rd1data1033_38_) );
  NOR2X1 U20640 ( .A(n33331), .B(n33332), .Y(n33330) );
  NAND3X1 U20641 ( .A(n33333), .B(n33334), .C(n33335), .Y(n33332) );
  NOR2X1 U20642 ( .A(n33336), .B(n33337), .Y(n33335) );
  OAI22X1 U20643 ( .A(n28993), .B(n25499), .C(n28994), .D(n25510), .Y(n33337)
         );
  OAI22X1 U20644 ( .A(n28995), .B(n25520), .C(n28996), .D(n25531), .Y(n33336)
         );
  AOI22X1 U20645 ( .A(n25541), .B(reg_file[1446]), .C(n25552), .D(
        reg_file[1318]), .Y(n33334) );
  AOI22X1 U20646 ( .A(n25563), .B(reg_file[1190]), .C(n25574), .D(
        reg_file[1062]), .Y(n33333) );
  NAND3X1 U20647 ( .A(n33338), .B(n33339), .C(n33340), .Y(n33331) );
  NOR2X1 U20648 ( .A(n33341), .B(n33342), .Y(n33340) );
  OAI22X1 U20649 ( .A(n29002), .B(n25585), .C(n29003), .D(n25596), .Y(n33342)
         );
  OAI22X1 U20650 ( .A(n29004), .B(n25606), .C(n29005), .D(n25617), .Y(n33341)
         );
  AOI22X1 U20651 ( .A(n25627), .B(reg_file[550]), .C(n25638), .D(reg_file[678]), .Y(n33339) );
  AOI22X1 U20652 ( .A(n25649), .B(reg_file[806]), .C(n25660), .D(reg_file[934]), .Y(n33338) );
  NOR2X1 U20653 ( .A(n33343), .B(n33344), .Y(n33329) );
  NAND3X1 U20654 ( .A(n33345), .B(n33346), .C(n33347), .Y(n33344) );
  NOR2X1 U20655 ( .A(n33348), .B(n33349), .Y(n33347) );
  OAI22X1 U20656 ( .A(n29013), .B(n25671), .C(n29014), .D(n25682), .Y(n33349)
         );
  OAI22X1 U20657 ( .A(n29015), .B(n25692), .C(n29016), .D(n25703), .Y(n33348)
         );
  AOI22X1 U20658 ( .A(n25713), .B(reg_file[3494]), .C(n25724), .D(
        reg_file[3366]), .Y(n33346) );
  AOI22X1 U20659 ( .A(n25735), .B(reg_file[3238]), .C(n25746), .D(
        reg_file[3110]), .Y(n33345) );
  NAND3X1 U20660 ( .A(n33350), .B(n33351), .C(n33352), .Y(n33343) );
  NOR2X1 U20661 ( .A(n33353), .B(n33354), .Y(n33352) );
  OAI22X1 U20662 ( .A(n29022), .B(n25757), .C(n29023), .D(n25768), .Y(n33354)
         );
  OAI22X1 U20663 ( .A(n29024), .B(n25778), .C(n29025), .D(n25789), .Y(n33353)
         );
  AOI22X1 U20664 ( .A(n25799), .B(reg_file[2470]), .C(n25810), .D(
        reg_file[2342]), .Y(n33351) );
  AOI22X1 U20665 ( .A(n25821), .B(reg_file[2214]), .C(n25832), .D(
        reg_file[2086]), .Y(n33350) );
  AOI21X1 U20666 ( .A(n33355), .B(n33356), .C(n25488), .Y(rd1data1033_37_) );
  NOR2X1 U20667 ( .A(n33357), .B(n33358), .Y(n33356) );
  NAND3X1 U20668 ( .A(n33359), .B(n33360), .C(n33361), .Y(n33358) );
  NOR2X1 U20669 ( .A(n33362), .B(n33363), .Y(n33361) );
  OAI22X1 U20670 ( .A(n29035), .B(n25499), .C(n29036), .D(n25510), .Y(n33363)
         );
  OAI22X1 U20671 ( .A(n29037), .B(n25520), .C(n29038), .D(n25531), .Y(n33362)
         );
  AOI22X1 U20672 ( .A(n25541), .B(reg_file[1445]), .C(n25552), .D(
        reg_file[1317]), .Y(n33360) );
  AOI22X1 U20673 ( .A(n25563), .B(reg_file[1189]), .C(n25574), .D(
        reg_file[1061]), .Y(n33359) );
  NAND3X1 U20674 ( .A(n33364), .B(n33365), .C(n33366), .Y(n33357) );
  NOR2X1 U20675 ( .A(n33367), .B(n33368), .Y(n33366) );
  OAI22X1 U20676 ( .A(n29044), .B(n25585), .C(n29045), .D(n25596), .Y(n33368)
         );
  OAI22X1 U20677 ( .A(n29046), .B(n25606), .C(n29047), .D(n25617), .Y(n33367)
         );
  AOI22X1 U20678 ( .A(n25627), .B(reg_file[549]), .C(n25638), .D(reg_file[677]), .Y(n33365) );
  AOI22X1 U20679 ( .A(n25649), .B(reg_file[805]), .C(n25660), .D(reg_file[933]), .Y(n33364) );
  NOR2X1 U20680 ( .A(n33369), .B(n33370), .Y(n33355) );
  NAND3X1 U20681 ( .A(n33371), .B(n33372), .C(n33373), .Y(n33370) );
  NOR2X1 U20682 ( .A(n33374), .B(n33375), .Y(n33373) );
  OAI22X1 U20683 ( .A(n29055), .B(n25671), .C(n29056), .D(n25682), .Y(n33375)
         );
  OAI22X1 U20684 ( .A(n29057), .B(n25692), .C(n29058), .D(n25703), .Y(n33374)
         );
  AOI22X1 U20685 ( .A(n25713), .B(reg_file[3493]), .C(n25724), .D(
        reg_file[3365]), .Y(n33372) );
  AOI22X1 U20686 ( .A(n25735), .B(reg_file[3237]), .C(n25746), .D(
        reg_file[3109]), .Y(n33371) );
  NAND3X1 U20687 ( .A(n33376), .B(n33377), .C(n33378), .Y(n33369) );
  NOR2X1 U20688 ( .A(n33379), .B(n33380), .Y(n33378) );
  OAI22X1 U20689 ( .A(n29064), .B(n25757), .C(n29065), .D(n25768), .Y(n33380)
         );
  OAI22X1 U20690 ( .A(n29066), .B(n25778), .C(n29067), .D(n25789), .Y(n33379)
         );
  AOI22X1 U20691 ( .A(n25799), .B(reg_file[2469]), .C(n25810), .D(
        reg_file[2341]), .Y(n33377) );
  AOI22X1 U20692 ( .A(n25821), .B(reg_file[2213]), .C(n25832), .D(
        reg_file[2085]), .Y(n33376) );
  AOI21X1 U20693 ( .A(n33381), .B(n33382), .C(n25488), .Y(rd1data1033_36_) );
  NOR2X1 U20694 ( .A(n33383), .B(n33384), .Y(n33382) );
  NAND3X1 U20695 ( .A(n33385), .B(n33386), .C(n33387), .Y(n33384) );
  NOR2X1 U20696 ( .A(n33388), .B(n33389), .Y(n33387) );
  OAI22X1 U20697 ( .A(n29077), .B(n25499), .C(n29078), .D(n25510), .Y(n33389)
         );
  OAI22X1 U20698 ( .A(n29079), .B(n25520), .C(n29080), .D(n25531), .Y(n33388)
         );
  AOI22X1 U20699 ( .A(n25541), .B(reg_file[1444]), .C(n25552), .D(
        reg_file[1316]), .Y(n33386) );
  AOI22X1 U20700 ( .A(n25563), .B(reg_file[1188]), .C(n25574), .D(
        reg_file[1060]), .Y(n33385) );
  NAND3X1 U20701 ( .A(n33390), .B(n33391), .C(n33392), .Y(n33383) );
  NOR2X1 U20702 ( .A(n33393), .B(n33394), .Y(n33392) );
  OAI22X1 U20703 ( .A(n29086), .B(n25585), .C(n29087), .D(n25596), .Y(n33394)
         );
  OAI22X1 U20704 ( .A(n29088), .B(n25606), .C(n29089), .D(n25617), .Y(n33393)
         );
  AOI22X1 U20705 ( .A(n25627), .B(reg_file[548]), .C(n25638), .D(reg_file[676]), .Y(n33391) );
  AOI22X1 U20706 ( .A(n25649), .B(reg_file[804]), .C(n25660), .D(reg_file[932]), .Y(n33390) );
  NOR2X1 U20707 ( .A(n33395), .B(n33396), .Y(n33381) );
  NAND3X1 U20708 ( .A(n33397), .B(n33398), .C(n33399), .Y(n33396) );
  NOR2X1 U20709 ( .A(n33400), .B(n33401), .Y(n33399) );
  OAI22X1 U20710 ( .A(n29097), .B(n25671), .C(n29098), .D(n25682), .Y(n33401)
         );
  OAI22X1 U20711 ( .A(n29099), .B(n25692), .C(n29100), .D(n25703), .Y(n33400)
         );
  AOI22X1 U20712 ( .A(n25713), .B(reg_file[3492]), .C(n25724), .D(
        reg_file[3364]), .Y(n33398) );
  AOI22X1 U20713 ( .A(n25735), .B(reg_file[3236]), .C(n25746), .D(
        reg_file[3108]), .Y(n33397) );
  NAND3X1 U20714 ( .A(n33402), .B(n33403), .C(n33404), .Y(n33395) );
  NOR2X1 U20715 ( .A(n33405), .B(n33406), .Y(n33404) );
  OAI22X1 U20716 ( .A(n29106), .B(n25757), .C(n29107), .D(n25768), .Y(n33406)
         );
  OAI22X1 U20717 ( .A(n29108), .B(n25778), .C(n29109), .D(n25789), .Y(n33405)
         );
  AOI22X1 U20718 ( .A(n25799), .B(reg_file[2468]), .C(n25810), .D(
        reg_file[2340]), .Y(n33403) );
  AOI22X1 U20719 ( .A(n25821), .B(reg_file[2212]), .C(n25832), .D(
        reg_file[2084]), .Y(n33402) );
  AOI21X1 U20720 ( .A(n33407), .B(n33408), .C(n25488), .Y(rd1data1033_35_) );
  NOR2X1 U20721 ( .A(n33409), .B(n33410), .Y(n33408) );
  NAND3X1 U20722 ( .A(n33411), .B(n33412), .C(n33413), .Y(n33410) );
  NOR2X1 U20723 ( .A(n33414), .B(n33415), .Y(n33413) );
  OAI22X1 U20724 ( .A(n29119), .B(n25499), .C(n29120), .D(n25510), .Y(n33415)
         );
  OAI22X1 U20725 ( .A(n29121), .B(n25520), .C(n29122), .D(n25531), .Y(n33414)
         );
  AOI22X1 U20726 ( .A(n25541), .B(reg_file[1443]), .C(n25552), .D(
        reg_file[1315]), .Y(n33412) );
  AOI22X1 U20727 ( .A(n25563), .B(reg_file[1187]), .C(n25574), .D(
        reg_file[1059]), .Y(n33411) );
  NAND3X1 U20728 ( .A(n33416), .B(n33417), .C(n33418), .Y(n33409) );
  NOR2X1 U20729 ( .A(n33419), .B(n33420), .Y(n33418) );
  OAI22X1 U20730 ( .A(n29128), .B(n25585), .C(n29129), .D(n25596), .Y(n33420)
         );
  OAI22X1 U20731 ( .A(n29130), .B(n25606), .C(n29131), .D(n25617), .Y(n33419)
         );
  AOI22X1 U20732 ( .A(n25627), .B(reg_file[547]), .C(n25638), .D(reg_file[675]), .Y(n33417) );
  AOI22X1 U20733 ( .A(n25649), .B(reg_file[803]), .C(n25660), .D(reg_file[931]), .Y(n33416) );
  NOR2X1 U20734 ( .A(n33421), .B(n33422), .Y(n33407) );
  NAND3X1 U20735 ( .A(n33423), .B(n33424), .C(n33425), .Y(n33422) );
  NOR2X1 U20736 ( .A(n33426), .B(n33427), .Y(n33425) );
  OAI22X1 U20737 ( .A(n29139), .B(n25671), .C(n29140), .D(n25682), .Y(n33427)
         );
  OAI22X1 U20738 ( .A(n29141), .B(n25692), .C(n29142), .D(n25703), .Y(n33426)
         );
  AOI22X1 U20739 ( .A(n25713), .B(reg_file[3491]), .C(n25724), .D(
        reg_file[3363]), .Y(n33424) );
  AOI22X1 U20740 ( .A(n25735), .B(reg_file[3235]), .C(n25746), .D(
        reg_file[3107]), .Y(n33423) );
  NAND3X1 U20741 ( .A(n33428), .B(n33429), .C(n33430), .Y(n33421) );
  NOR2X1 U20742 ( .A(n33431), .B(n33432), .Y(n33430) );
  OAI22X1 U20743 ( .A(n29148), .B(n25757), .C(n29149), .D(n25768), .Y(n33432)
         );
  OAI22X1 U20744 ( .A(n29150), .B(n25778), .C(n29151), .D(n25789), .Y(n33431)
         );
  AOI22X1 U20745 ( .A(n25799), .B(reg_file[2467]), .C(n25810), .D(
        reg_file[2339]), .Y(n33429) );
  AOI22X1 U20746 ( .A(n25821), .B(reg_file[2211]), .C(n25832), .D(
        reg_file[2083]), .Y(n33428) );
  AOI21X1 U20747 ( .A(n33433), .B(n33434), .C(n25488), .Y(rd1data1033_34_) );
  NOR2X1 U20748 ( .A(n33435), .B(n33436), .Y(n33434) );
  NAND3X1 U20749 ( .A(n33437), .B(n33438), .C(n33439), .Y(n33436) );
  NOR2X1 U20750 ( .A(n33440), .B(n33441), .Y(n33439) );
  OAI22X1 U20751 ( .A(n29161), .B(n25499), .C(n29162), .D(n25510), .Y(n33441)
         );
  OAI22X1 U20752 ( .A(n29163), .B(n25520), .C(n29164), .D(n25531), .Y(n33440)
         );
  AOI22X1 U20753 ( .A(n25541), .B(reg_file[1442]), .C(n25552), .D(
        reg_file[1314]), .Y(n33438) );
  AOI22X1 U20754 ( .A(n25563), .B(reg_file[1186]), .C(n25574), .D(
        reg_file[1058]), .Y(n33437) );
  NAND3X1 U20755 ( .A(n33442), .B(n33443), .C(n33444), .Y(n33435) );
  NOR2X1 U20756 ( .A(n33445), .B(n33446), .Y(n33444) );
  OAI22X1 U20757 ( .A(n29170), .B(n25585), .C(n29171), .D(n25596), .Y(n33446)
         );
  OAI22X1 U20758 ( .A(n29172), .B(n25606), .C(n29173), .D(n25617), .Y(n33445)
         );
  AOI22X1 U20759 ( .A(n25627), .B(reg_file[546]), .C(n25638), .D(reg_file[674]), .Y(n33443) );
  AOI22X1 U20760 ( .A(n25649), .B(reg_file[802]), .C(n25660), .D(reg_file[930]), .Y(n33442) );
  NOR2X1 U20761 ( .A(n33447), .B(n33448), .Y(n33433) );
  NAND3X1 U20762 ( .A(n33449), .B(n33450), .C(n33451), .Y(n33448) );
  NOR2X1 U20763 ( .A(n33452), .B(n33453), .Y(n33451) );
  OAI22X1 U20764 ( .A(n29181), .B(n25671), .C(n29182), .D(n25682), .Y(n33453)
         );
  OAI22X1 U20765 ( .A(n29183), .B(n25692), .C(n29184), .D(n25703), .Y(n33452)
         );
  AOI22X1 U20766 ( .A(n25713), .B(reg_file[3490]), .C(n25724), .D(
        reg_file[3362]), .Y(n33450) );
  AOI22X1 U20767 ( .A(n25735), .B(reg_file[3234]), .C(n25746), .D(
        reg_file[3106]), .Y(n33449) );
  NAND3X1 U20768 ( .A(n33454), .B(n33455), .C(n33456), .Y(n33447) );
  NOR2X1 U20769 ( .A(n33457), .B(n33458), .Y(n33456) );
  OAI22X1 U20770 ( .A(n29190), .B(n25757), .C(n29191), .D(n25768), .Y(n33458)
         );
  OAI22X1 U20771 ( .A(n29192), .B(n25778), .C(n29193), .D(n25789), .Y(n33457)
         );
  AOI22X1 U20772 ( .A(n25799), .B(reg_file[2466]), .C(n25810), .D(
        reg_file[2338]), .Y(n33455) );
  AOI22X1 U20773 ( .A(n25821), .B(reg_file[2210]), .C(n25832), .D(
        reg_file[2082]), .Y(n33454) );
  AOI21X1 U20774 ( .A(n33459), .B(n33460), .C(n25488), .Y(rd1data1033_33_) );
  NOR2X1 U20775 ( .A(n33461), .B(n33462), .Y(n33460) );
  NAND3X1 U20776 ( .A(n33463), .B(n33464), .C(n33465), .Y(n33462) );
  NOR2X1 U20777 ( .A(n33466), .B(n33467), .Y(n33465) );
  OAI22X1 U20778 ( .A(n29203), .B(n25499), .C(n29204), .D(n25510), .Y(n33467)
         );
  OAI22X1 U20779 ( .A(n29205), .B(n25520), .C(n29206), .D(n25531), .Y(n33466)
         );
  AOI22X1 U20780 ( .A(n25541), .B(reg_file[1441]), .C(n25552), .D(
        reg_file[1313]), .Y(n33464) );
  AOI22X1 U20781 ( .A(n25563), .B(reg_file[1185]), .C(n25574), .D(
        reg_file[1057]), .Y(n33463) );
  NAND3X1 U20782 ( .A(n33468), .B(n33469), .C(n33470), .Y(n33461) );
  NOR2X1 U20783 ( .A(n33471), .B(n33472), .Y(n33470) );
  OAI22X1 U20784 ( .A(n29212), .B(n25585), .C(n29213), .D(n25596), .Y(n33472)
         );
  OAI22X1 U20785 ( .A(n29214), .B(n25606), .C(n29215), .D(n25617), .Y(n33471)
         );
  AOI22X1 U20786 ( .A(n25627), .B(reg_file[545]), .C(n25638), .D(reg_file[673]), .Y(n33469) );
  AOI22X1 U20787 ( .A(n25649), .B(reg_file[801]), .C(n25660), .D(reg_file[929]), .Y(n33468) );
  NOR2X1 U20788 ( .A(n33473), .B(n33474), .Y(n33459) );
  NAND3X1 U20789 ( .A(n33475), .B(n33476), .C(n33477), .Y(n33474) );
  NOR2X1 U20790 ( .A(n33478), .B(n33479), .Y(n33477) );
  OAI22X1 U20791 ( .A(n29223), .B(n25671), .C(n29224), .D(n25682), .Y(n33479)
         );
  OAI22X1 U20792 ( .A(n29225), .B(n25692), .C(n29226), .D(n25703), .Y(n33478)
         );
  AOI22X1 U20793 ( .A(n25713), .B(reg_file[3489]), .C(n25724), .D(
        reg_file[3361]), .Y(n33476) );
  AOI22X1 U20794 ( .A(n25735), .B(reg_file[3233]), .C(n25746), .D(
        reg_file[3105]), .Y(n33475) );
  NAND3X1 U20795 ( .A(n33480), .B(n33481), .C(n33482), .Y(n33473) );
  NOR2X1 U20796 ( .A(n33483), .B(n33484), .Y(n33482) );
  OAI22X1 U20797 ( .A(n29232), .B(n25757), .C(n29233), .D(n25768), .Y(n33484)
         );
  OAI22X1 U20798 ( .A(n29234), .B(n25778), .C(n29235), .D(n25789), .Y(n33483)
         );
  AOI22X1 U20799 ( .A(n25799), .B(reg_file[2465]), .C(n25810), .D(
        reg_file[2337]), .Y(n33481) );
  AOI22X1 U20800 ( .A(n25821), .B(reg_file[2209]), .C(n25832), .D(
        reg_file[2081]), .Y(n33480) );
  AOI21X1 U20801 ( .A(n33485), .B(n33486), .C(n25488), .Y(rd1data1033_32_) );
  NOR2X1 U20802 ( .A(n33487), .B(n33488), .Y(n33486) );
  NAND3X1 U20803 ( .A(n33489), .B(n33490), .C(n33491), .Y(n33488) );
  NOR2X1 U20804 ( .A(n33492), .B(n33493), .Y(n33491) );
  OAI22X1 U20805 ( .A(n29245), .B(n25499), .C(n29246), .D(n25510), .Y(n33493)
         );
  OAI22X1 U20806 ( .A(n29247), .B(n25520), .C(n29248), .D(n25531), .Y(n33492)
         );
  AOI22X1 U20807 ( .A(n25541), .B(reg_file[1440]), .C(n25552), .D(
        reg_file[1312]), .Y(n33490) );
  AOI22X1 U20808 ( .A(n25563), .B(reg_file[1184]), .C(n25574), .D(
        reg_file[1056]), .Y(n33489) );
  NAND3X1 U20809 ( .A(n33494), .B(n33495), .C(n33496), .Y(n33487) );
  NOR2X1 U20810 ( .A(n33497), .B(n33498), .Y(n33496) );
  OAI22X1 U20811 ( .A(n29254), .B(n25585), .C(n29255), .D(n25596), .Y(n33498)
         );
  OAI22X1 U20812 ( .A(n29256), .B(n25606), .C(n29257), .D(n25617), .Y(n33497)
         );
  AOI22X1 U20813 ( .A(n25627), .B(reg_file[544]), .C(n25638), .D(reg_file[672]), .Y(n33495) );
  AOI22X1 U20814 ( .A(n25649), .B(reg_file[800]), .C(n25660), .D(reg_file[928]), .Y(n33494) );
  NOR2X1 U20815 ( .A(n33499), .B(n33500), .Y(n33485) );
  NAND3X1 U20816 ( .A(n33501), .B(n33502), .C(n33503), .Y(n33500) );
  NOR2X1 U20817 ( .A(n33504), .B(n33505), .Y(n33503) );
  OAI22X1 U20818 ( .A(n29265), .B(n25671), .C(n29266), .D(n25682), .Y(n33505)
         );
  OAI22X1 U20819 ( .A(n29267), .B(n25692), .C(n29268), .D(n25703), .Y(n33504)
         );
  AOI22X1 U20820 ( .A(n25713), .B(reg_file[3488]), .C(n25724), .D(
        reg_file[3360]), .Y(n33502) );
  AOI22X1 U20821 ( .A(n25735), .B(reg_file[3232]), .C(n25746), .D(
        reg_file[3104]), .Y(n33501) );
  NAND3X1 U20822 ( .A(n33506), .B(n33507), .C(n33508), .Y(n33499) );
  NOR2X1 U20823 ( .A(n33509), .B(n33510), .Y(n33508) );
  OAI22X1 U20824 ( .A(n29274), .B(n25757), .C(n29275), .D(n25768), .Y(n33510)
         );
  OAI22X1 U20825 ( .A(n29276), .B(n25778), .C(n29277), .D(n25789), .Y(n33509)
         );
  AOI22X1 U20826 ( .A(n25799), .B(reg_file[2464]), .C(n25810), .D(
        reg_file[2336]), .Y(n33507) );
  AOI22X1 U20827 ( .A(n25821), .B(reg_file[2208]), .C(n25832), .D(
        reg_file[2080]), .Y(n33506) );
  AOI21X1 U20828 ( .A(n33511), .B(n33512), .C(n25488), .Y(rd1data1033_31_) );
  NOR2X1 U20829 ( .A(n33513), .B(n33514), .Y(n33512) );
  NAND3X1 U20830 ( .A(n33515), .B(n33516), .C(n33517), .Y(n33514) );
  NOR2X1 U20831 ( .A(n33518), .B(n33519), .Y(n33517) );
  OAI22X1 U20832 ( .A(n29287), .B(n25499), .C(n29288), .D(n25510), .Y(n33519)
         );
  OAI22X1 U20833 ( .A(n29289), .B(n25520), .C(n29290), .D(n25531), .Y(n33518)
         );
  AOI22X1 U20834 ( .A(n25541), .B(reg_file[1439]), .C(n25552), .D(
        reg_file[1311]), .Y(n33516) );
  AOI22X1 U20835 ( .A(n25563), .B(reg_file[1183]), .C(n25574), .D(
        reg_file[1055]), .Y(n33515) );
  NAND3X1 U20836 ( .A(n33520), .B(n33521), .C(n33522), .Y(n33513) );
  NOR2X1 U20837 ( .A(n33523), .B(n33524), .Y(n33522) );
  OAI22X1 U20838 ( .A(n29296), .B(n25585), .C(n29297), .D(n25596), .Y(n33524)
         );
  OAI22X1 U20839 ( .A(n29298), .B(n25606), .C(n29299), .D(n25617), .Y(n33523)
         );
  AOI22X1 U20840 ( .A(n25627), .B(reg_file[543]), .C(n25638), .D(reg_file[671]), .Y(n33521) );
  AOI22X1 U20841 ( .A(n25649), .B(reg_file[799]), .C(n25660), .D(reg_file[927]), .Y(n33520) );
  NOR2X1 U20842 ( .A(n33525), .B(n33526), .Y(n33511) );
  NAND3X1 U20843 ( .A(n33527), .B(n33528), .C(n33529), .Y(n33526) );
  NOR2X1 U20844 ( .A(n33530), .B(n33531), .Y(n33529) );
  OAI22X1 U20845 ( .A(n29307), .B(n25671), .C(n29308), .D(n25682), .Y(n33531)
         );
  OAI22X1 U20846 ( .A(n29309), .B(n25692), .C(n29310), .D(n25703), .Y(n33530)
         );
  AOI22X1 U20847 ( .A(n25713), .B(reg_file[3487]), .C(n25724), .D(
        reg_file[3359]), .Y(n33528) );
  AOI22X1 U20848 ( .A(n25735), .B(reg_file[3231]), .C(n25746), .D(
        reg_file[3103]), .Y(n33527) );
  NAND3X1 U20849 ( .A(n33532), .B(n33533), .C(n33534), .Y(n33525) );
  NOR2X1 U20850 ( .A(n33535), .B(n33536), .Y(n33534) );
  OAI22X1 U20851 ( .A(n29316), .B(n25757), .C(n29317), .D(n25768), .Y(n33536)
         );
  OAI22X1 U20852 ( .A(n29318), .B(n25778), .C(n29319), .D(n25789), .Y(n33535)
         );
  AOI22X1 U20853 ( .A(n25799), .B(reg_file[2463]), .C(n25810), .D(
        reg_file[2335]), .Y(n33533) );
  AOI22X1 U20854 ( .A(n25821), .B(reg_file[2207]), .C(n25832), .D(
        reg_file[2079]), .Y(n33532) );
  AOI21X1 U20855 ( .A(n33537), .B(n33538), .C(n25488), .Y(rd1data1033_30_) );
  NOR2X1 U20856 ( .A(n33539), .B(n33540), .Y(n33538) );
  NAND3X1 U20857 ( .A(n33541), .B(n33542), .C(n33543), .Y(n33540) );
  NOR2X1 U20858 ( .A(n33544), .B(n33545), .Y(n33543) );
  OAI22X1 U20859 ( .A(n29329), .B(n25499), .C(n29330), .D(n25509), .Y(n33545)
         );
  OAI22X1 U20860 ( .A(n29331), .B(n25520), .C(n29332), .D(n25530), .Y(n33544)
         );
  AOI22X1 U20861 ( .A(n25541), .B(reg_file[1438]), .C(n25552), .D(
        reg_file[1310]), .Y(n33542) );
  AOI22X1 U20862 ( .A(n25563), .B(reg_file[1182]), .C(n25574), .D(
        reg_file[1054]), .Y(n33541) );
  NAND3X1 U20863 ( .A(n33546), .B(n33547), .C(n33548), .Y(n33539) );
  NOR2X1 U20864 ( .A(n33549), .B(n33550), .Y(n33548) );
  OAI22X1 U20865 ( .A(n29338), .B(n25585), .C(n29339), .D(n25595), .Y(n33550)
         );
  OAI22X1 U20866 ( .A(n29340), .B(n25606), .C(n29341), .D(n25616), .Y(n33549)
         );
  AOI22X1 U20867 ( .A(n25627), .B(reg_file[542]), .C(n25638), .D(reg_file[670]), .Y(n33547) );
  AOI22X1 U20868 ( .A(n25649), .B(reg_file[798]), .C(n25660), .D(reg_file[926]), .Y(n33546) );
  NOR2X1 U20869 ( .A(n33551), .B(n33552), .Y(n33537) );
  NAND3X1 U20870 ( .A(n33553), .B(n33554), .C(n33555), .Y(n33552) );
  NOR2X1 U20871 ( .A(n33556), .B(n33557), .Y(n33555) );
  OAI22X1 U20872 ( .A(n29349), .B(n25671), .C(n29350), .D(n25681), .Y(n33557)
         );
  OAI22X1 U20873 ( .A(n29351), .B(n25692), .C(n29352), .D(n25702), .Y(n33556)
         );
  AOI22X1 U20874 ( .A(n25713), .B(reg_file[3486]), .C(n25724), .D(
        reg_file[3358]), .Y(n33554) );
  AOI22X1 U20875 ( .A(n25735), .B(reg_file[3230]), .C(n25746), .D(
        reg_file[3102]), .Y(n33553) );
  NAND3X1 U20876 ( .A(n33558), .B(n33559), .C(n33560), .Y(n33551) );
  NOR2X1 U20877 ( .A(n33561), .B(n33562), .Y(n33560) );
  OAI22X1 U20878 ( .A(n29358), .B(n25757), .C(n29359), .D(n25767), .Y(n33562)
         );
  OAI22X1 U20879 ( .A(n29360), .B(n25778), .C(n29361), .D(n25788), .Y(n33561)
         );
  AOI22X1 U20880 ( .A(n25799), .B(reg_file[2462]), .C(n25810), .D(
        reg_file[2334]), .Y(n33559) );
  AOI22X1 U20881 ( .A(n25821), .B(reg_file[2206]), .C(n25832), .D(
        reg_file[2078]), .Y(n33558) );
  AOI21X1 U20882 ( .A(n33563), .B(n33564), .C(n25488), .Y(rd1data1033_2_) );
  NOR2X1 U20883 ( .A(n33565), .B(n33566), .Y(n33564) );
  NAND3X1 U20884 ( .A(n33567), .B(n33568), .C(n33569), .Y(n33566) );
  NOR2X1 U20885 ( .A(n33570), .B(n33571), .Y(n33569) );
  OAI22X1 U20886 ( .A(n29371), .B(n25499), .C(n29372), .D(n25509), .Y(n33571)
         );
  OAI22X1 U20887 ( .A(n29373), .B(n25520), .C(n29374), .D(n25530), .Y(n33570)
         );
  AOI22X1 U20888 ( .A(n25541), .B(reg_file[1410]), .C(n25552), .D(
        reg_file[1282]), .Y(n33568) );
  AOI22X1 U20889 ( .A(n25563), .B(reg_file[1154]), .C(n25574), .D(
        reg_file[1026]), .Y(n33567) );
  NAND3X1 U20890 ( .A(n33572), .B(n33573), .C(n33574), .Y(n33565) );
  NOR2X1 U20891 ( .A(n33575), .B(n33576), .Y(n33574) );
  OAI22X1 U20892 ( .A(n29380), .B(n25585), .C(n29381), .D(n25595), .Y(n33576)
         );
  OAI22X1 U20893 ( .A(n29382), .B(n25606), .C(n29383), .D(n25616), .Y(n33575)
         );
  AOI22X1 U20894 ( .A(n25627), .B(reg_file[514]), .C(n25638), .D(reg_file[642]), .Y(n33573) );
  AOI22X1 U20895 ( .A(n25649), .B(reg_file[770]), .C(n25660), .D(reg_file[898]), .Y(n33572) );
  NOR2X1 U20896 ( .A(n33577), .B(n33578), .Y(n33563) );
  NAND3X1 U20897 ( .A(n33579), .B(n33580), .C(n33581), .Y(n33578) );
  NOR2X1 U20898 ( .A(n33582), .B(n33583), .Y(n33581) );
  OAI22X1 U20899 ( .A(n29391), .B(n25671), .C(n29392), .D(n25681), .Y(n33583)
         );
  OAI22X1 U20900 ( .A(n29393), .B(n25692), .C(n29394), .D(n25702), .Y(n33582)
         );
  AOI22X1 U20901 ( .A(n25713), .B(reg_file[3458]), .C(n25724), .D(
        reg_file[3330]), .Y(n33580) );
  AOI22X1 U20902 ( .A(n25735), .B(reg_file[3202]), .C(n25746), .D(
        reg_file[3074]), .Y(n33579) );
  NAND3X1 U20903 ( .A(n33584), .B(n33585), .C(n33586), .Y(n33577) );
  NOR2X1 U20904 ( .A(n33587), .B(n33588), .Y(n33586) );
  OAI22X1 U20905 ( .A(n29400), .B(n25757), .C(n29401), .D(n25767), .Y(n33588)
         );
  OAI22X1 U20906 ( .A(n29402), .B(n25778), .C(n29403), .D(n25788), .Y(n33587)
         );
  AOI22X1 U20907 ( .A(n25799), .B(reg_file[2434]), .C(n25810), .D(
        reg_file[2306]), .Y(n33585) );
  AOI22X1 U20908 ( .A(n25821), .B(reg_file[2178]), .C(n25832), .D(
        reg_file[2050]), .Y(n33584) );
  AOI21X1 U20909 ( .A(n33589), .B(n33590), .C(n25488), .Y(rd1data1033_29_) );
  NOR2X1 U20910 ( .A(n33591), .B(n33592), .Y(n33590) );
  NAND3X1 U20911 ( .A(n33593), .B(n33594), .C(n33595), .Y(n33592) );
  NOR2X1 U20912 ( .A(n33596), .B(n33597), .Y(n33595) );
  OAI22X1 U20913 ( .A(n29413), .B(n25499), .C(n29414), .D(n25509), .Y(n33597)
         );
  OAI22X1 U20914 ( .A(n29415), .B(n25520), .C(n29416), .D(n25530), .Y(n33596)
         );
  AOI22X1 U20915 ( .A(n25541), .B(reg_file[1437]), .C(n25552), .D(
        reg_file[1309]), .Y(n33594) );
  AOI22X1 U20916 ( .A(n25563), .B(reg_file[1181]), .C(n25574), .D(
        reg_file[1053]), .Y(n33593) );
  NAND3X1 U20917 ( .A(n33598), .B(n33599), .C(n33600), .Y(n33591) );
  NOR2X1 U20918 ( .A(n33601), .B(n33602), .Y(n33600) );
  OAI22X1 U20919 ( .A(n29422), .B(n25585), .C(n29423), .D(n25595), .Y(n33602)
         );
  OAI22X1 U20920 ( .A(n29424), .B(n25606), .C(n29425), .D(n25616), .Y(n33601)
         );
  AOI22X1 U20921 ( .A(n25627), .B(reg_file[541]), .C(n25638), .D(reg_file[669]), .Y(n33599) );
  AOI22X1 U20922 ( .A(n25649), .B(reg_file[797]), .C(n25660), .D(reg_file[925]), .Y(n33598) );
  NOR2X1 U20923 ( .A(n33603), .B(n33604), .Y(n33589) );
  NAND3X1 U20924 ( .A(n33605), .B(n33606), .C(n33607), .Y(n33604) );
  NOR2X1 U20925 ( .A(n33608), .B(n33609), .Y(n33607) );
  OAI22X1 U20926 ( .A(n29433), .B(n25671), .C(n29434), .D(n25681), .Y(n33609)
         );
  OAI22X1 U20927 ( .A(n29435), .B(n25692), .C(n29436), .D(n25702), .Y(n33608)
         );
  AOI22X1 U20928 ( .A(n25713), .B(reg_file[3485]), .C(n25724), .D(
        reg_file[3357]), .Y(n33606) );
  AOI22X1 U20929 ( .A(n25735), .B(reg_file[3229]), .C(n25746), .D(
        reg_file[3101]), .Y(n33605) );
  NAND3X1 U20930 ( .A(n33610), .B(n33611), .C(n33612), .Y(n33603) );
  NOR2X1 U20931 ( .A(n33613), .B(n33614), .Y(n33612) );
  OAI22X1 U20932 ( .A(n29442), .B(n25757), .C(n29443), .D(n25767), .Y(n33614)
         );
  OAI22X1 U20933 ( .A(n29444), .B(n25778), .C(n29445), .D(n25788), .Y(n33613)
         );
  AOI22X1 U20934 ( .A(n25799), .B(reg_file[2461]), .C(n25810), .D(
        reg_file[2333]), .Y(n33611) );
  AOI22X1 U20935 ( .A(n25821), .B(reg_file[2205]), .C(n25832), .D(
        reg_file[2077]), .Y(n33610) );
  AOI21X1 U20936 ( .A(n33615), .B(n33616), .C(n25488), .Y(rd1data1033_28_) );
  NOR2X1 U20937 ( .A(n33617), .B(n33618), .Y(n33616) );
  NAND3X1 U20938 ( .A(n33619), .B(n33620), .C(n33621), .Y(n33618) );
  NOR2X1 U20939 ( .A(n33622), .B(n33623), .Y(n33621) );
  OAI22X1 U20940 ( .A(n29455), .B(n25499), .C(n29456), .D(n25509), .Y(n33623)
         );
  OAI22X1 U20941 ( .A(n29457), .B(n25520), .C(n29458), .D(n25530), .Y(n33622)
         );
  AOI22X1 U20942 ( .A(n25541), .B(reg_file[1436]), .C(n25552), .D(
        reg_file[1308]), .Y(n33620) );
  AOI22X1 U20943 ( .A(n25563), .B(reg_file[1180]), .C(n25574), .D(
        reg_file[1052]), .Y(n33619) );
  NAND3X1 U20944 ( .A(n33624), .B(n33625), .C(n33626), .Y(n33617) );
  NOR2X1 U20945 ( .A(n33627), .B(n33628), .Y(n33626) );
  OAI22X1 U20946 ( .A(n29464), .B(n25585), .C(n29465), .D(n25595), .Y(n33628)
         );
  OAI22X1 U20947 ( .A(n29466), .B(n25606), .C(n29467), .D(n25616), .Y(n33627)
         );
  AOI22X1 U20948 ( .A(n25627), .B(reg_file[540]), .C(n25638), .D(reg_file[668]), .Y(n33625) );
  AOI22X1 U20949 ( .A(n25649), .B(reg_file[796]), .C(n25660), .D(reg_file[924]), .Y(n33624) );
  NOR2X1 U20950 ( .A(n33629), .B(n33630), .Y(n33615) );
  NAND3X1 U20951 ( .A(n33631), .B(n33632), .C(n33633), .Y(n33630) );
  NOR2X1 U20952 ( .A(n33634), .B(n33635), .Y(n33633) );
  OAI22X1 U20953 ( .A(n29475), .B(n25671), .C(n29476), .D(n25681), .Y(n33635)
         );
  OAI22X1 U20954 ( .A(n29477), .B(n25692), .C(n29478), .D(n25702), .Y(n33634)
         );
  AOI22X1 U20955 ( .A(n25713), .B(reg_file[3484]), .C(n25724), .D(
        reg_file[3356]), .Y(n33632) );
  AOI22X1 U20956 ( .A(n25735), .B(reg_file[3228]), .C(n25746), .D(
        reg_file[3100]), .Y(n33631) );
  NAND3X1 U20957 ( .A(n33636), .B(n33637), .C(n33638), .Y(n33629) );
  NOR2X1 U20958 ( .A(n33639), .B(n33640), .Y(n33638) );
  OAI22X1 U20959 ( .A(n29484), .B(n25757), .C(n29485), .D(n25767), .Y(n33640)
         );
  OAI22X1 U20960 ( .A(n29486), .B(n25778), .C(n29487), .D(n25788), .Y(n33639)
         );
  AOI22X1 U20961 ( .A(n25799), .B(reg_file[2460]), .C(n25810), .D(
        reg_file[2332]), .Y(n33637) );
  AOI22X1 U20962 ( .A(n25821), .B(reg_file[2204]), .C(n25832), .D(
        reg_file[2076]), .Y(n33636) );
  AOI21X1 U20963 ( .A(n33641), .B(n33642), .C(n25487), .Y(rd1data1033_27_) );
  NOR2X1 U20964 ( .A(n33643), .B(n33644), .Y(n33642) );
  NAND3X1 U20965 ( .A(n33645), .B(n33646), .C(n33647), .Y(n33644) );
  NOR2X1 U20966 ( .A(n33648), .B(n33649), .Y(n33647) );
  OAI22X1 U20967 ( .A(n29497), .B(n25498), .C(n29498), .D(n25509), .Y(n33649)
         );
  OAI22X1 U20968 ( .A(n29499), .B(n25519), .C(n29500), .D(n25530), .Y(n33648)
         );
  AOI22X1 U20969 ( .A(n25540), .B(reg_file[1435]), .C(n25551), .D(
        reg_file[1307]), .Y(n33646) );
  AOI22X1 U20970 ( .A(n25562), .B(reg_file[1179]), .C(n25573), .D(
        reg_file[1051]), .Y(n33645) );
  NAND3X1 U20971 ( .A(n33650), .B(n33651), .C(n33652), .Y(n33643) );
  NOR2X1 U20972 ( .A(n33653), .B(n33654), .Y(n33652) );
  OAI22X1 U20973 ( .A(n29506), .B(n25584), .C(n29507), .D(n25595), .Y(n33654)
         );
  OAI22X1 U20974 ( .A(n29508), .B(n25605), .C(n29509), .D(n25616), .Y(n33653)
         );
  AOI22X1 U20975 ( .A(n25626), .B(reg_file[539]), .C(n25637), .D(reg_file[667]), .Y(n33651) );
  AOI22X1 U20976 ( .A(n25648), .B(reg_file[795]), .C(n25659), .D(reg_file[923]), .Y(n33650) );
  NOR2X1 U20977 ( .A(n33655), .B(n33656), .Y(n33641) );
  NAND3X1 U20978 ( .A(n33657), .B(n33658), .C(n33659), .Y(n33656) );
  NOR2X1 U20979 ( .A(n33660), .B(n33661), .Y(n33659) );
  OAI22X1 U20980 ( .A(n29517), .B(n25670), .C(n29518), .D(n25681), .Y(n33661)
         );
  OAI22X1 U20981 ( .A(n29519), .B(n25691), .C(n29520), .D(n25702), .Y(n33660)
         );
  AOI22X1 U20982 ( .A(n25712), .B(reg_file[3483]), .C(n25723), .D(
        reg_file[3355]), .Y(n33658) );
  AOI22X1 U20983 ( .A(n25734), .B(reg_file[3227]), .C(n25745), .D(
        reg_file[3099]), .Y(n33657) );
  NAND3X1 U20984 ( .A(n33662), .B(n33663), .C(n33664), .Y(n33655) );
  NOR2X1 U20985 ( .A(n33665), .B(n33666), .Y(n33664) );
  OAI22X1 U20986 ( .A(n29526), .B(n25756), .C(n29527), .D(n25767), .Y(n33666)
         );
  OAI22X1 U20987 ( .A(n29528), .B(n25777), .C(n29529), .D(n25788), .Y(n33665)
         );
  AOI22X1 U20988 ( .A(n25798), .B(reg_file[2459]), .C(n25809), .D(
        reg_file[2331]), .Y(n33663) );
  AOI22X1 U20989 ( .A(n25820), .B(reg_file[2203]), .C(n25831), .D(
        reg_file[2075]), .Y(n33662) );
  AOI21X1 U20990 ( .A(n33667), .B(n33668), .C(n25487), .Y(rd1data1033_26_) );
  NOR2X1 U20991 ( .A(n33669), .B(n33670), .Y(n33668) );
  NAND3X1 U20992 ( .A(n33671), .B(n33672), .C(n33673), .Y(n33670) );
  NOR2X1 U20993 ( .A(n33674), .B(n33675), .Y(n33673) );
  OAI22X1 U20994 ( .A(n29539), .B(n25498), .C(n29540), .D(n25509), .Y(n33675)
         );
  OAI22X1 U20995 ( .A(n29541), .B(n25519), .C(n29542), .D(n25530), .Y(n33674)
         );
  AOI22X1 U20996 ( .A(n25540), .B(reg_file[1434]), .C(n25551), .D(
        reg_file[1306]), .Y(n33672) );
  AOI22X1 U20997 ( .A(n25562), .B(reg_file[1178]), .C(n25573), .D(
        reg_file[1050]), .Y(n33671) );
  NAND3X1 U20998 ( .A(n33676), .B(n33677), .C(n33678), .Y(n33669) );
  NOR2X1 U20999 ( .A(n33679), .B(n33680), .Y(n33678) );
  OAI22X1 U21000 ( .A(n29548), .B(n25584), .C(n29549), .D(n25595), .Y(n33680)
         );
  OAI22X1 U21001 ( .A(n29550), .B(n25605), .C(n29551), .D(n25616), .Y(n33679)
         );
  AOI22X1 U21002 ( .A(n25626), .B(reg_file[538]), .C(n25637), .D(reg_file[666]), .Y(n33677) );
  AOI22X1 U21003 ( .A(n25648), .B(reg_file[794]), .C(n25659), .D(reg_file[922]), .Y(n33676) );
  NOR2X1 U21004 ( .A(n33681), .B(n33682), .Y(n33667) );
  NAND3X1 U21005 ( .A(n33683), .B(n33684), .C(n33685), .Y(n33682) );
  NOR2X1 U21006 ( .A(n33686), .B(n33687), .Y(n33685) );
  OAI22X1 U21007 ( .A(n29559), .B(n25670), .C(n29560), .D(n25681), .Y(n33687)
         );
  OAI22X1 U21008 ( .A(n29561), .B(n25691), .C(n29562), .D(n25702), .Y(n33686)
         );
  AOI22X1 U21009 ( .A(n25712), .B(reg_file[3482]), .C(n25723), .D(
        reg_file[3354]), .Y(n33684) );
  AOI22X1 U21010 ( .A(n25734), .B(reg_file[3226]), .C(n25745), .D(
        reg_file[3098]), .Y(n33683) );
  NAND3X1 U21011 ( .A(n33688), .B(n33689), .C(n33690), .Y(n33681) );
  NOR2X1 U21012 ( .A(n33691), .B(n33692), .Y(n33690) );
  OAI22X1 U21013 ( .A(n29568), .B(n25756), .C(n29569), .D(n25767), .Y(n33692)
         );
  OAI22X1 U21014 ( .A(n29570), .B(n25777), .C(n29571), .D(n25788), .Y(n33691)
         );
  AOI22X1 U21015 ( .A(n25798), .B(reg_file[2458]), .C(n25809), .D(
        reg_file[2330]), .Y(n33689) );
  AOI22X1 U21016 ( .A(n25820), .B(reg_file[2202]), .C(n25831), .D(
        reg_file[2074]), .Y(n33688) );
  AOI21X1 U21017 ( .A(n33693), .B(n33694), .C(n25487), .Y(rd1data1033_25_) );
  NOR2X1 U21018 ( .A(n33695), .B(n33696), .Y(n33694) );
  NAND3X1 U21019 ( .A(n33697), .B(n33698), .C(n33699), .Y(n33696) );
  NOR2X1 U21020 ( .A(n33700), .B(n33701), .Y(n33699) );
  OAI22X1 U21021 ( .A(n29581), .B(n25498), .C(n29582), .D(n25509), .Y(n33701)
         );
  OAI22X1 U21022 ( .A(n29583), .B(n25519), .C(n29584), .D(n25530), .Y(n33700)
         );
  AOI22X1 U21023 ( .A(n25540), .B(reg_file[1433]), .C(n25551), .D(
        reg_file[1305]), .Y(n33698) );
  AOI22X1 U21024 ( .A(n25562), .B(reg_file[1177]), .C(n25573), .D(
        reg_file[1049]), .Y(n33697) );
  NAND3X1 U21025 ( .A(n33702), .B(n33703), .C(n33704), .Y(n33695) );
  NOR2X1 U21026 ( .A(n33705), .B(n33706), .Y(n33704) );
  OAI22X1 U21027 ( .A(n29590), .B(n25584), .C(n29591), .D(n25595), .Y(n33706)
         );
  OAI22X1 U21028 ( .A(n29592), .B(n25605), .C(n29593), .D(n25616), .Y(n33705)
         );
  AOI22X1 U21029 ( .A(n25626), .B(reg_file[537]), .C(n25637), .D(reg_file[665]), .Y(n33703) );
  AOI22X1 U21030 ( .A(n25648), .B(reg_file[793]), .C(n25659), .D(reg_file[921]), .Y(n33702) );
  NOR2X1 U21031 ( .A(n33707), .B(n33708), .Y(n33693) );
  NAND3X1 U21032 ( .A(n33709), .B(n33710), .C(n33711), .Y(n33708) );
  NOR2X1 U21033 ( .A(n33712), .B(n33713), .Y(n33711) );
  OAI22X1 U21034 ( .A(n29601), .B(n25670), .C(n29602), .D(n25681), .Y(n33713)
         );
  OAI22X1 U21035 ( .A(n29603), .B(n25691), .C(n29604), .D(n25702), .Y(n33712)
         );
  AOI22X1 U21036 ( .A(n25712), .B(reg_file[3481]), .C(n25723), .D(
        reg_file[3353]), .Y(n33710) );
  AOI22X1 U21037 ( .A(n25734), .B(reg_file[3225]), .C(n25745), .D(
        reg_file[3097]), .Y(n33709) );
  NAND3X1 U21038 ( .A(n33714), .B(n33715), .C(n33716), .Y(n33707) );
  NOR2X1 U21039 ( .A(n33717), .B(n33718), .Y(n33716) );
  OAI22X1 U21040 ( .A(n29610), .B(n25756), .C(n29611), .D(n25767), .Y(n33718)
         );
  OAI22X1 U21041 ( .A(n29612), .B(n25777), .C(n29613), .D(n25788), .Y(n33717)
         );
  AOI22X1 U21042 ( .A(n25798), .B(reg_file[2457]), .C(n25809), .D(
        reg_file[2329]), .Y(n33715) );
  AOI22X1 U21043 ( .A(n25820), .B(reg_file[2201]), .C(n25831), .D(
        reg_file[2073]), .Y(n33714) );
  AOI21X1 U21044 ( .A(n33719), .B(n33720), .C(n25487), .Y(rd1data1033_24_) );
  NOR2X1 U21045 ( .A(n33721), .B(n33722), .Y(n33720) );
  NAND3X1 U21046 ( .A(n33723), .B(n33724), .C(n33725), .Y(n33722) );
  NOR2X1 U21047 ( .A(n33726), .B(n33727), .Y(n33725) );
  OAI22X1 U21048 ( .A(n29623), .B(n25498), .C(n29624), .D(n25509), .Y(n33727)
         );
  OAI22X1 U21049 ( .A(n29625), .B(n25519), .C(n29626), .D(n25530), .Y(n33726)
         );
  AOI22X1 U21050 ( .A(n25540), .B(reg_file[1432]), .C(n25551), .D(
        reg_file[1304]), .Y(n33724) );
  AOI22X1 U21051 ( .A(n25562), .B(reg_file[1176]), .C(n25573), .D(
        reg_file[1048]), .Y(n33723) );
  NAND3X1 U21052 ( .A(n33728), .B(n33729), .C(n33730), .Y(n33721) );
  NOR2X1 U21053 ( .A(n33731), .B(n33732), .Y(n33730) );
  OAI22X1 U21054 ( .A(n29632), .B(n25584), .C(n29633), .D(n25595), .Y(n33732)
         );
  OAI22X1 U21055 ( .A(n29634), .B(n25605), .C(n29635), .D(n25616), .Y(n33731)
         );
  AOI22X1 U21056 ( .A(n25626), .B(reg_file[536]), .C(n25637), .D(reg_file[664]), .Y(n33729) );
  AOI22X1 U21057 ( .A(n25648), .B(reg_file[792]), .C(n25659), .D(reg_file[920]), .Y(n33728) );
  NOR2X1 U21058 ( .A(n33733), .B(n33734), .Y(n33719) );
  NAND3X1 U21059 ( .A(n33735), .B(n33736), .C(n33737), .Y(n33734) );
  NOR2X1 U21060 ( .A(n33738), .B(n33739), .Y(n33737) );
  OAI22X1 U21061 ( .A(n29643), .B(n25670), .C(n29644), .D(n25681), .Y(n33739)
         );
  OAI22X1 U21062 ( .A(n29645), .B(n25691), .C(n29646), .D(n25702), .Y(n33738)
         );
  AOI22X1 U21063 ( .A(n25712), .B(reg_file[3480]), .C(n25723), .D(
        reg_file[3352]), .Y(n33736) );
  AOI22X1 U21064 ( .A(n25734), .B(reg_file[3224]), .C(n25745), .D(
        reg_file[3096]), .Y(n33735) );
  NAND3X1 U21065 ( .A(n33740), .B(n33741), .C(n33742), .Y(n33733) );
  NOR2X1 U21066 ( .A(n33743), .B(n33744), .Y(n33742) );
  OAI22X1 U21067 ( .A(n29652), .B(n25756), .C(n29653), .D(n25767), .Y(n33744)
         );
  OAI22X1 U21068 ( .A(n29654), .B(n25777), .C(n29655), .D(n25788), .Y(n33743)
         );
  AOI22X1 U21069 ( .A(n25798), .B(reg_file[2456]), .C(n25809), .D(
        reg_file[2328]), .Y(n33741) );
  AOI22X1 U21070 ( .A(n25820), .B(reg_file[2200]), .C(n25831), .D(
        reg_file[2072]), .Y(n33740) );
  AOI21X1 U21071 ( .A(n33745), .B(n33746), .C(n25487), .Y(rd1data1033_23_) );
  NOR2X1 U21072 ( .A(n33747), .B(n33748), .Y(n33746) );
  NAND3X1 U21073 ( .A(n33749), .B(n33750), .C(n33751), .Y(n33748) );
  NOR2X1 U21074 ( .A(n33752), .B(n33753), .Y(n33751) );
  OAI22X1 U21075 ( .A(n29665), .B(n25498), .C(n29666), .D(n25509), .Y(n33753)
         );
  OAI22X1 U21076 ( .A(n29667), .B(n25519), .C(n29668), .D(n25530), .Y(n33752)
         );
  AOI22X1 U21077 ( .A(n25540), .B(reg_file[1431]), .C(n25551), .D(
        reg_file[1303]), .Y(n33750) );
  AOI22X1 U21078 ( .A(n25562), .B(reg_file[1175]), .C(n25573), .D(
        reg_file[1047]), .Y(n33749) );
  NAND3X1 U21079 ( .A(n33754), .B(n33755), .C(n33756), .Y(n33747) );
  NOR2X1 U21080 ( .A(n33757), .B(n33758), .Y(n33756) );
  OAI22X1 U21081 ( .A(n29674), .B(n25584), .C(n29675), .D(n25595), .Y(n33758)
         );
  OAI22X1 U21082 ( .A(n29676), .B(n25605), .C(n29677), .D(n25616), .Y(n33757)
         );
  AOI22X1 U21083 ( .A(n25626), .B(reg_file[535]), .C(n25637), .D(reg_file[663]), .Y(n33755) );
  AOI22X1 U21084 ( .A(n25648), .B(reg_file[791]), .C(n25659), .D(reg_file[919]), .Y(n33754) );
  NOR2X1 U21085 ( .A(n33759), .B(n33760), .Y(n33745) );
  NAND3X1 U21086 ( .A(n33761), .B(n33762), .C(n33763), .Y(n33760) );
  NOR2X1 U21087 ( .A(n33764), .B(n33765), .Y(n33763) );
  OAI22X1 U21088 ( .A(n29685), .B(n25670), .C(n29686), .D(n25681), .Y(n33765)
         );
  OAI22X1 U21089 ( .A(n29687), .B(n25691), .C(n29688), .D(n25702), .Y(n33764)
         );
  AOI22X1 U21090 ( .A(n25712), .B(reg_file[3479]), .C(n25723), .D(
        reg_file[3351]), .Y(n33762) );
  AOI22X1 U21091 ( .A(n25734), .B(reg_file[3223]), .C(n25745), .D(
        reg_file[3095]), .Y(n33761) );
  NAND3X1 U21092 ( .A(n33766), .B(n33767), .C(n33768), .Y(n33759) );
  NOR2X1 U21093 ( .A(n33769), .B(n33770), .Y(n33768) );
  OAI22X1 U21094 ( .A(n29694), .B(n25756), .C(n29695), .D(n25767), .Y(n33770)
         );
  OAI22X1 U21095 ( .A(n29696), .B(n25777), .C(n29697), .D(n25788), .Y(n33769)
         );
  AOI22X1 U21096 ( .A(n25798), .B(reg_file[2455]), .C(n25809), .D(
        reg_file[2327]), .Y(n33767) );
  AOI22X1 U21097 ( .A(n25820), .B(reg_file[2199]), .C(n25831), .D(
        reg_file[2071]), .Y(n33766) );
  AOI21X1 U21098 ( .A(n33771), .B(n33772), .C(n25487), .Y(rd1data1033_22_) );
  NOR2X1 U21099 ( .A(n33773), .B(n33774), .Y(n33772) );
  NAND3X1 U21100 ( .A(n33775), .B(n33776), .C(n33777), .Y(n33774) );
  NOR2X1 U21101 ( .A(n33778), .B(n33779), .Y(n33777) );
  OAI22X1 U21102 ( .A(n29707), .B(n25498), .C(n29708), .D(n25509), .Y(n33779)
         );
  OAI22X1 U21103 ( .A(n29709), .B(n25519), .C(n29710), .D(n25530), .Y(n33778)
         );
  AOI22X1 U21104 ( .A(n25540), .B(reg_file[1430]), .C(n25551), .D(
        reg_file[1302]), .Y(n33776) );
  AOI22X1 U21105 ( .A(n25562), .B(reg_file[1174]), .C(n25573), .D(
        reg_file[1046]), .Y(n33775) );
  NAND3X1 U21106 ( .A(n33780), .B(n33781), .C(n33782), .Y(n33773) );
  NOR2X1 U21107 ( .A(n33783), .B(n33784), .Y(n33782) );
  OAI22X1 U21108 ( .A(n29716), .B(n25584), .C(n29717), .D(n25595), .Y(n33784)
         );
  OAI22X1 U21109 ( .A(n29718), .B(n25605), .C(n29719), .D(n25616), .Y(n33783)
         );
  AOI22X1 U21110 ( .A(n25626), .B(reg_file[534]), .C(n25637), .D(reg_file[662]), .Y(n33781) );
  AOI22X1 U21111 ( .A(n25648), .B(reg_file[790]), .C(n25659), .D(reg_file[918]), .Y(n33780) );
  NOR2X1 U21112 ( .A(n33785), .B(n33786), .Y(n33771) );
  NAND3X1 U21113 ( .A(n33787), .B(n33788), .C(n33789), .Y(n33786) );
  NOR2X1 U21114 ( .A(n33790), .B(n33791), .Y(n33789) );
  OAI22X1 U21115 ( .A(n29727), .B(n25670), .C(n29728), .D(n25681), .Y(n33791)
         );
  OAI22X1 U21116 ( .A(n29729), .B(n25691), .C(n29730), .D(n25702), .Y(n33790)
         );
  AOI22X1 U21117 ( .A(n25712), .B(reg_file[3478]), .C(n25723), .D(
        reg_file[3350]), .Y(n33788) );
  AOI22X1 U21118 ( .A(n25734), .B(reg_file[3222]), .C(n25745), .D(
        reg_file[3094]), .Y(n33787) );
  NAND3X1 U21119 ( .A(n33792), .B(n33793), .C(n33794), .Y(n33785) );
  NOR2X1 U21120 ( .A(n33795), .B(n33796), .Y(n33794) );
  OAI22X1 U21121 ( .A(n29736), .B(n25756), .C(n29737), .D(n25767), .Y(n33796)
         );
  OAI22X1 U21122 ( .A(n29738), .B(n25777), .C(n29739), .D(n25788), .Y(n33795)
         );
  AOI22X1 U21123 ( .A(n25798), .B(reg_file[2454]), .C(n25809), .D(
        reg_file[2326]), .Y(n33793) );
  AOI22X1 U21124 ( .A(n25820), .B(reg_file[2198]), .C(n25831), .D(
        reg_file[2070]), .Y(n33792) );
  AOI21X1 U21125 ( .A(n33797), .B(n33798), .C(n25487), .Y(rd1data1033_21_) );
  NOR2X1 U21126 ( .A(n33799), .B(n33800), .Y(n33798) );
  NAND3X1 U21127 ( .A(n33801), .B(n33802), .C(n33803), .Y(n33800) );
  NOR2X1 U21128 ( .A(n33804), .B(n33805), .Y(n33803) );
  OAI22X1 U21129 ( .A(n29749), .B(n25498), .C(n29750), .D(n25509), .Y(n33805)
         );
  OAI22X1 U21130 ( .A(n29751), .B(n25519), .C(n29752), .D(n25530), .Y(n33804)
         );
  AOI22X1 U21131 ( .A(n25540), .B(reg_file[1429]), .C(n25551), .D(
        reg_file[1301]), .Y(n33802) );
  AOI22X1 U21132 ( .A(n25562), .B(reg_file[1173]), .C(n25573), .D(
        reg_file[1045]), .Y(n33801) );
  NAND3X1 U21133 ( .A(n33806), .B(n33807), .C(n33808), .Y(n33799) );
  NOR2X1 U21134 ( .A(n33809), .B(n33810), .Y(n33808) );
  OAI22X1 U21135 ( .A(n29758), .B(n25584), .C(n29759), .D(n25595), .Y(n33810)
         );
  OAI22X1 U21136 ( .A(n29760), .B(n25605), .C(n29761), .D(n25616), .Y(n33809)
         );
  AOI22X1 U21137 ( .A(n25626), .B(reg_file[533]), .C(n25637), .D(reg_file[661]), .Y(n33807) );
  AOI22X1 U21138 ( .A(n25648), .B(reg_file[789]), .C(n25659), .D(reg_file[917]), .Y(n33806) );
  NOR2X1 U21139 ( .A(n33811), .B(n33812), .Y(n33797) );
  NAND3X1 U21140 ( .A(n33813), .B(n33814), .C(n33815), .Y(n33812) );
  NOR2X1 U21141 ( .A(n33816), .B(n33817), .Y(n33815) );
  OAI22X1 U21142 ( .A(n29769), .B(n25670), .C(n29770), .D(n25681), .Y(n33817)
         );
  OAI22X1 U21143 ( .A(n29771), .B(n25691), .C(n29772), .D(n25702), .Y(n33816)
         );
  AOI22X1 U21144 ( .A(n25712), .B(reg_file[3477]), .C(n25723), .D(
        reg_file[3349]), .Y(n33814) );
  AOI22X1 U21145 ( .A(n25734), .B(reg_file[3221]), .C(n25745), .D(
        reg_file[3093]), .Y(n33813) );
  NAND3X1 U21146 ( .A(n33818), .B(n33819), .C(n33820), .Y(n33811) );
  NOR2X1 U21147 ( .A(n33821), .B(n33822), .Y(n33820) );
  OAI22X1 U21148 ( .A(n29778), .B(n25756), .C(n29779), .D(n25767), .Y(n33822)
         );
  OAI22X1 U21149 ( .A(n29780), .B(n25777), .C(n29781), .D(n25788), .Y(n33821)
         );
  AOI22X1 U21150 ( .A(n25798), .B(reg_file[2453]), .C(n25809), .D(
        reg_file[2325]), .Y(n33819) );
  AOI22X1 U21151 ( .A(n25820), .B(reg_file[2197]), .C(n25831), .D(
        reg_file[2069]), .Y(n33818) );
  AOI21X1 U21152 ( .A(n33823), .B(n33824), .C(n25487), .Y(rd1data1033_20_) );
  NOR2X1 U21153 ( .A(n33825), .B(n33826), .Y(n33824) );
  NAND3X1 U21154 ( .A(n33827), .B(n33828), .C(n33829), .Y(n33826) );
  NOR2X1 U21155 ( .A(n33830), .B(n33831), .Y(n33829) );
  OAI22X1 U21156 ( .A(n29791), .B(n25498), .C(n29792), .D(n25509), .Y(n33831)
         );
  OAI22X1 U21157 ( .A(n29793), .B(n25519), .C(n29794), .D(n25530), .Y(n33830)
         );
  AOI22X1 U21158 ( .A(n25540), .B(reg_file[1428]), .C(n25551), .D(
        reg_file[1300]), .Y(n33828) );
  AOI22X1 U21159 ( .A(n25562), .B(reg_file[1172]), .C(n25573), .D(
        reg_file[1044]), .Y(n33827) );
  NAND3X1 U21160 ( .A(n33832), .B(n33833), .C(n33834), .Y(n33825) );
  NOR2X1 U21161 ( .A(n33835), .B(n33836), .Y(n33834) );
  OAI22X1 U21162 ( .A(n29800), .B(n25584), .C(n29801), .D(n25595), .Y(n33836)
         );
  OAI22X1 U21163 ( .A(n29802), .B(n25605), .C(n29803), .D(n25616), .Y(n33835)
         );
  AOI22X1 U21164 ( .A(n25626), .B(reg_file[532]), .C(n25637), .D(reg_file[660]), .Y(n33833) );
  AOI22X1 U21165 ( .A(n25648), .B(reg_file[788]), .C(n25659), .D(reg_file[916]), .Y(n33832) );
  NOR2X1 U21166 ( .A(n33837), .B(n33838), .Y(n33823) );
  NAND3X1 U21167 ( .A(n33839), .B(n33840), .C(n33841), .Y(n33838) );
  NOR2X1 U21168 ( .A(n33842), .B(n33843), .Y(n33841) );
  OAI22X1 U21169 ( .A(n29811), .B(n25670), .C(n29812), .D(n25681), .Y(n33843)
         );
  OAI22X1 U21170 ( .A(n29813), .B(n25691), .C(n29814), .D(n25702), .Y(n33842)
         );
  AOI22X1 U21171 ( .A(n25712), .B(reg_file[3476]), .C(n25723), .D(
        reg_file[3348]), .Y(n33840) );
  AOI22X1 U21172 ( .A(n25734), .B(reg_file[3220]), .C(n25745), .D(
        reg_file[3092]), .Y(n33839) );
  NAND3X1 U21173 ( .A(n33844), .B(n33845), .C(n33846), .Y(n33837) );
  NOR2X1 U21174 ( .A(n33847), .B(n33848), .Y(n33846) );
  OAI22X1 U21175 ( .A(n29820), .B(n25756), .C(n29821), .D(n25767), .Y(n33848)
         );
  OAI22X1 U21176 ( .A(n29822), .B(n25777), .C(n29823), .D(n25788), .Y(n33847)
         );
  AOI22X1 U21177 ( .A(n25798), .B(reg_file[2452]), .C(n25809), .D(
        reg_file[2324]), .Y(n33845) );
  AOI22X1 U21178 ( .A(n25820), .B(reg_file[2196]), .C(n25831), .D(
        reg_file[2068]), .Y(n33844) );
  AOI21X1 U21179 ( .A(n33849), .B(n33850), .C(n25487), .Y(rd1data1033_1_) );
  NOR2X1 U21180 ( .A(n33851), .B(n33852), .Y(n33850) );
  NAND3X1 U21181 ( .A(n33853), .B(n33854), .C(n33855), .Y(n33852) );
  NOR2X1 U21182 ( .A(n33856), .B(n33857), .Y(n33855) );
  OAI22X1 U21183 ( .A(n29833), .B(n25498), .C(n29834), .D(n25509), .Y(n33857)
         );
  OAI22X1 U21184 ( .A(n29835), .B(n25519), .C(n29836), .D(n25530), .Y(n33856)
         );
  AOI22X1 U21185 ( .A(n25540), .B(reg_file[1409]), .C(n25551), .D(
        reg_file[1281]), .Y(n33854) );
  AOI22X1 U21186 ( .A(n25562), .B(reg_file[1153]), .C(n25573), .D(
        reg_file[1025]), .Y(n33853) );
  NAND3X1 U21187 ( .A(n33858), .B(n33859), .C(n33860), .Y(n33851) );
  NOR2X1 U21188 ( .A(n33861), .B(n33862), .Y(n33860) );
  OAI22X1 U21189 ( .A(n29842), .B(n25584), .C(n29843), .D(n25595), .Y(n33862)
         );
  OAI22X1 U21190 ( .A(n29844), .B(n25605), .C(n29845), .D(n25616), .Y(n33861)
         );
  AOI22X1 U21191 ( .A(n25626), .B(reg_file[513]), .C(n25637), .D(reg_file[641]), .Y(n33859) );
  AOI22X1 U21192 ( .A(n25648), .B(reg_file[769]), .C(n25659), .D(reg_file[897]), .Y(n33858) );
  NOR2X1 U21193 ( .A(n33863), .B(n33864), .Y(n33849) );
  NAND3X1 U21194 ( .A(n33865), .B(n33866), .C(n33867), .Y(n33864) );
  NOR2X1 U21195 ( .A(n33868), .B(n33869), .Y(n33867) );
  OAI22X1 U21196 ( .A(n29853), .B(n25670), .C(n29854), .D(n25681), .Y(n33869)
         );
  OAI22X1 U21197 ( .A(n29855), .B(n25691), .C(n29856), .D(n25702), .Y(n33868)
         );
  AOI22X1 U21198 ( .A(n25712), .B(reg_file[3457]), .C(n25723), .D(
        reg_file[3329]), .Y(n33866) );
  AOI22X1 U21199 ( .A(n25734), .B(reg_file[3201]), .C(n25745), .D(
        reg_file[3073]), .Y(n33865) );
  NAND3X1 U21200 ( .A(n33870), .B(n33871), .C(n33872), .Y(n33863) );
  NOR2X1 U21201 ( .A(n33873), .B(n33874), .Y(n33872) );
  OAI22X1 U21202 ( .A(n29862), .B(n25756), .C(n29863), .D(n25767), .Y(n33874)
         );
  OAI22X1 U21203 ( .A(n29864), .B(n25777), .C(n29865), .D(n25788), .Y(n33873)
         );
  AOI22X1 U21204 ( .A(n25798), .B(reg_file[2433]), .C(n25809), .D(
        reg_file[2305]), .Y(n33871) );
  AOI22X1 U21205 ( .A(n25820), .B(reg_file[2177]), .C(n25831), .D(
        reg_file[2049]), .Y(n33870) );
  AOI21X1 U21206 ( .A(n33875), .B(n33876), .C(n25487), .Y(rd1data1033_19_) );
  NOR2X1 U21207 ( .A(n33877), .B(n33878), .Y(n33876) );
  NAND3X1 U21208 ( .A(n33879), .B(n33880), .C(n33881), .Y(n33878) );
  NOR2X1 U21209 ( .A(n33882), .B(n33883), .Y(n33881) );
  OAI22X1 U21210 ( .A(n29875), .B(n25498), .C(n29876), .D(n25508), .Y(n33883)
         );
  OAI22X1 U21211 ( .A(n29877), .B(n25519), .C(n29878), .D(n25529), .Y(n33882)
         );
  AOI22X1 U21212 ( .A(n25540), .B(reg_file[1427]), .C(n25551), .D(
        reg_file[1299]), .Y(n33880) );
  AOI22X1 U21213 ( .A(n25562), .B(reg_file[1171]), .C(n25573), .D(
        reg_file[1043]), .Y(n33879) );
  NAND3X1 U21214 ( .A(n33884), .B(n33885), .C(n33886), .Y(n33877) );
  NOR2X1 U21215 ( .A(n33887), .B(n33888), .Y(n33886) );
  OAI22X1 U21216 ( .A(n29884), .B(n25584), .C(n29885), .D(n25594), .Y(n33888)
         );
  OAI22X1 U21217 ( .A(n29886), .B(n25605), .C(n29887), .D(n25615), .Y(n33887)
         );
  AOI22X1 U21218 ( .A(n25626), .B(reg_file[531]), .C(n25637), .D(reg_file[659]), .Y(n33885) );
  AOI22X1 U21219 ( .A(n25648), .B(reg_file[787]), .C(n25659), .D(reg_file[915]), .Y(n33884) );
  NOR2X1 U21220 ( .A(n33889), .B(n33890), .Y(n33875) );
  NAND3X1 U21221 ( .A(n33891), .B(n33892), .C(n33893), .Y(n33890) );
  NOR2X1 U21222 ( .A(n33894), .B(n33895), .Y(n33893) );
  OAI22X1 U21223 ( .A(n29895), .B(n25670), .C(n29896), .D(n25680), .Y(n33895)
         );
  OAI22X1 U21224 ( .A(n29897), .B(n25691), .C(n29898), .D(n25701), .Y(n33894)
         );
  AOI22X1 U21225 ( .A(n25712), .B(reg_file[3475]), .C(n25723), .D(
        reg_file[3347]), .Y(n33892) );
  AOI22X1 U21226 ( .A(n25734), .B(reg_file[3219]), .C(n25745), .D(
        reg_file[3091]), .Y(n33891) );
  NAND3X1 U21227 ( .A(n33896), .B(n33897), .C(n33898), .Y(n33889) );
  NOR2X1 U21228 ( .A(n33899), .B(n33900), .Y(n33898) );
  OAI22X1 U21229 ( .A(n29904), .B(n25756), .C(n29905), .D(n25766), .Y(n33900)
         );
  OAI22X1 U21230 ( .A(n29906), .B(n25777), .C(n29907), .D(n25787), .Y(n33899)
         );
  AOI22X1 U21231 ( .A(n25798), .B(reg_file[2451]), .C(n25809), .D(
        reg_file[2323]), .Y(n33897) );
  AOI22X1 U21232 ( .A(n25820), .B(reg_file[2195]), .C(n25831), .D(
        reg_file[2067]), .Y(n33896) );
  AOI21X1 U21233 ( .A(n33901), .B(n33902), .C(n25487), .Y(rd1data1033_18_) );
  NOR2X1 U21234 ( .A(n33903), .B(n33904), .Y(n33902) );
  NAND3X1 U21235 ( .A(n33905), .B(n33906), .C(n33907), .Y(n33904) );
  NOR2X1 U21236 ( .A(n33908), .B(n33909), .Y(n33907) );
  OAI22X1 U21237 ( .A(n29917), .B(n25498), .C(n29918), .D(n25508), .Y(n33909)
         );
  OAI22X1 U21238 ( .A(n29919), .B(n25519), .C(n29920), .D(n25529), .Y(n33908)
         );
  AOI22X1 U21239 ( .A(n25540), .B(reg_file[1426]), .C(n25551), .D(
        reg_file[1298]), .Y(n33906) );
  AOI22X1 U21240 ( .A(n25562), .B(reg_file[1170]), .C(n25573), .D(
        reg_file[1042]), .Y(n33905) );
  NAND3X1 U21241 ( .A(n33910), .B(n33911), .C(n33912), .Y(n33903) );
  NOR2X1 U21242 ( .A(n33913), .B(n33914), .Y(n33912) );
  OAI22X1 U21243 ( .A(n29926), .B(n25584), .C(n29927), .D(n25594), .Y(n33914)
         );
  OAI22X1 U21244 ( .A(n29928), .B(n25605), .C(n29929), .D(n25615), .Y(n33913)
         );
  AOI22X1 U21245 ( .A(n25626), .B(reg_file[530]), .C(n25637), .D(reg_file[658]), .Y(n33911) );
  AOI22X1 U21246 ( .A(n25648), .B(reg_file[786]), .C(n25659), .D(reg_file[914]), .Y(n33910) );
  NOR2X1 U21247 ( .A(n33915), .B(n33916), .Y(n33901) );
  NAND3X1 U21248 ( .A(n33917), .B(n33918), .C(n33919), .Y(n33916) );
  NOR2X1 U21249 ( .A(n33920), .B(n33921), .Y(n33919) );
  OAI22X1 U21250 ( .A(n29937), .B(n25670), .C(n29938), .D(n25680), .Y(n33921)
         );
  OAI22X1 U21251 ( .A(n29939), .B(n25691), .C(n29940), .D(n25701), .Y(n33920)
         );
  AOI22X1 U21252 ( .A(n25712), .B(reg_file[3474]), .C(n25723), .D(
        reg_file[3346]), .Y(n33918) );
  AOI22X1 U21253 ( .A(n25734), .B(reg_file[3218]), .C(n25745), .D(
        reg_file[3090]), .Y(n33917) );
  NAND3X1 U21254 ( .A(n33922), .B(n33923), .C(n33924), .Y(n33915) );
  NOR2X1 U21255 ( .A(n33925), .B(n33926), .Y(n33924) );
  OAI22X1 U21256 ( .A(n29946), .B(n25756), .C(n29947), .D(n25766), .Y(n33926)
         );
  OAI22X1 U21257 ( .A(n29948), .B(n25777), .C(n29949), .D(n25787), .Y(n33925)
         );
  AOI22X1 U21258 ( .A(n25798), .B(reg_file[2450]), .C(n25809), .D(
        reg_file[2322]), .Y(n33923) );
  AOI22X1 U21259 ( .A(n25820), .B(reg_file[2194]), .C(n25831), .D(
        reg_file[2066]), .Y(n33922) );
  AOI21X1 U21260 ( .A(n33927), .B(n33928), .C(n25487), .Y(rd1data1033_17_) );
  NOR2X1 U21261 ( .A(n33929), .B(n33930), .Y(n33928) );
  NAND3X1 U21262 ( .A(n33931), .B(n33932), .C(n33933), .Y(n33930) );
  NOR2X1 U21263 ( .A(n33934), .B(n33935), .Y(n33933) );
  OAI22X1 U21264 ( .A(n29959), .B(n25498), .C(n29960), .D(n25508), .Y(n33935)
         );
  OAI22X1 U21265 ( .A(n29961), .B(n25519), .C(n29962), .D(n25529), .Y(n33934)
         );
  AOI22X1 U21266 ( .A(n25540), .B(reg_file[1425]), .C(n25551), .D(
        reg_file[1297]), .Y(n33932) );
  AOI22X1 U21267 ( .A(n25562), .B(reg_file[1169]), .C(n25573), .D(
        reg_file[1041]), .Y(n33931) );
  NAND3X1 U21268 ( .A(n33936), .B(n33937), .C(n33938), .Y(n33929) );
  NOR2X1 U21269 ( .A(n33939), .B(n33940), .Y(n33938) );
  OAI22X1 U21270 ( .A(n29968), .B(n25584), .C(n29969), .D(n25594), .Y(n33940)
         );
  OAI22X1 U21271 ( .A(n29970), .B(n25605), .C(n29971), .D(n25615), .Y(n33939)
         );
  AOI22X1 U21272 ( .A(n25626), .B(reg_file[529]), .C(n25637), .D(reg_file[657]), .Y(n33937) );
  AOI22X1 U21273 ( .A(n25648), .B(reg_file[785]), .C(n25659), .D(reg_file[913]), .Y(n33936) );
  NOR2X1 U21274 ( .A(n33941), .B(n33942), .Y(n33927) );
  NAND3X1 U21275 ( .A(n33943), .B(n33944), .C(n33945), .Y(n33942) );
  NOR2X1 U21276 ( .A(n33946), .B(n33947), .Y(n33945) );
  OAI22X1 U21277 ( .A(n29979), .B(n25670), .C(n29980), .D(n25680), .Y(n33947)
         );
  OAI22X1 U21278 ( .A(n29981), .B(n25691), .C(n29982), .D(n25701), .Y(n33946)
         );
  AOI22X1 U21279 ( .A(n25712), .B(reg_file[3473]), .C(n25723), .D(
        reg_file[3345]), .Y(n33944) );
  AOI22X1 U21280 ( .A(n25734), .B(reg_file[3217]), .C(n25745), .D(
        reg_file[3089]), .Y(n33943) );
  NAND3X1 U21281 ( .A(n33948), .B(n33949), .C(n33950), .Y(n33941) );
  NOR2X1 U21282 ( .A(n33951), .B(n33952), .Y(n33950) );
  OAI22X1 U21283 ( .A(n29988), .B(n25756), .C(n29989), .D(n25766), .Y(n33952)
         );
  OAI22X1 U21284 ( .A(n29990), .B(n25777), .C(n29991), .D(n25787), .Y(n33951)
         );
  AOI22X1 U21285 ( .A(n25798), .B(reg_file[2449]), .C(n25809), .D(
        reg_file[2321]), .Y(n33949) );
  AOI22X1 U21286 ( .A(n25820), .B(reg_file[2193]), .C(n25831), .D(
        reg_file[2065]), .Y(n33948) );
  AOI21X1 U21287 ( .A(n33953), .B(n33954), .C(n25486), .Y(rd1data1033_16_) );
  NOR2X1 U21288 ( .A(n33955), .B(n33956), .Y(n33954) );
  NAND3X1 U21289 ( .A(n33957), .B(n33958), .C(n33959), .Y(n33956) );
  NOR2X1 U21290 ( .A(n33960), .B(n33961), .Y(n33959) );
  OAI22X1 U21291 ( .A(n30001), .B(n25497), .C(n30002), .D(n25508), .Y(n33961)
         );
  OAI22X1 U21292 ( .A(n30003), .B(n25518), .C(n30004), .D(n25529), .Y(n33960)
         );
  AOI22X1 U21293 ( .A(n25539), .B(reg_file[1424]), .C(n25550), .D(
        reg_file[1296]), .Y(n33958) );
  AOI22X1 U21294 ( .A(n25561), .B(reg_file[1168]), .C(n25572), .D(
        reg_file[1040]), .Y(n33957) );
  NAND3X1 U21295 ( .A(n33962), .B(n33963), .C(n33964), .Y(n33955) );
  NOR2X1 U21296 ( .A(n33965), .B(n33966), .Y(n33964) );
  OAI22X1 U21297 ( .A(n30010), .B(n25583), .C(n30011), .D(n25594), .Y(n33966)
         );
  OAI22X1 U21298 ( .A(n30012), .B(n25604), .C(n30013), .D(n25615), .Y(n33965)
         );
  AOI22X1 U21299 ( .A(n25625), .B(reg_file[528]), .C(n25636), .D(reg_file[656]), .Y(n33963) );
  AOI22X1 U21300 ( .A(n25647), .B(reg_file[784]), .C(n25658), .D(reg_file[912]), .Y(n33962) );
  NOR2X1 U21301 ( .A(n33967), .B(n33968), .Y(n33953) );
  NAND3X1 U21302 ( .A(n33969), .B(n33970), .C(n33971), .Y(n33968) );
  NOR2X1 U21303 ( .A(n33972), .B(n33973), .Y(n33971) );
  OAI22X1 U21304 ( .A(n30021), .B(n25669), .C(n30022), .D(n25680), .Y(n33973)
         );
  OAI22X1 U21305 ( .A(n30023), .B(n25690), .C(n30024), .D(n25701), .Y(n33972)
         );
  AOI22X1 U21306 ( .A(n25711), .B(reg_file[3472]), .C(n25722), .D(
        reg_file[3344]), .Y(n33970) );
  AOI22X1 U21307 ( .A(n25733), .B(reg_file[3216]), .C(n25744), .D(
        reg_file[3088]), .Y(n33969) );
  NAND3X1 U21308 ( .A(n33974), .B(n33975), .C(n33976), .Y(n33967) );
  NOR2X1 U21309 ( .A(n33977), .B(n33978), .Y(n33976) );
  OAI22X1 U21310 ( .A(n30030), .B(n25755), .C(n30031), .D(n25766), .Y(n33978)
         );
  OAI22X1 U21311 ( .A(n30032), .B(n25776), .C(n30033), .D(n25787), .Y(n33977)
         );
  AOI22X1 U21312 ( .A(n25797), .B(reg_file[2448]), .C(n25808), .D(
        reg_file[2320]), .Y(n33975) );
  AOI22X1 U21313 ( .A(n25819), .B(reg_file[2192]), .C(n25830), .D(
        reg_file[2064]), .Y(n33974) );
  AOI21X1 U21314 ( .A(n33979), .B(n33980), .C(n25486), .Y(rd1data1033_15_) );
  NOR2X1 U21315 ( .A(n33981), .B(n33982), .Y(n33980) );
  NAND3X1 U21316 ( .A(n33983), .B(n33984), .C(n33985), .Y(n33982) );
  NOR2X1 U21317 ( .A(n33986), .B(n33987), .Y(n33985) );
  OAI22X1 U21318 ( .A(n30043), .B(n25497), .C(n30044), .D(n25508), .Y(n33987)
         );
  OAI22X1 U21319 ( .A(n30045), .B(n25518), .C(n30046), .D(n25529), .Y(n33986)
         );
  AOI22X1 U21320 ( .A(n25539), .B(reg_file[1423]), .C(n25550), .D(
        reg_file[1295]), .Y(n33984) );
  AOI22X1 U21321 ( .A(n25561), .B(reg_file[1167]), .C(n25572), .D(
        reg_file[1039]), .Y(n33983) );
  NAND3X1 U21322 ( .A(n33988), .B(n33989), .C(n33990), .Y(n33981) );
  NOR2X1 U21323 ( .A(n33991), .B(n33992), .Y(n33990) );
  OAI22X1 U21324 ( .A(n30052), .B(n25583), .C(n30053), .D(n25594), .Y(n33992)
         );
  OAI22X1 U21325 ( .A(n30054), .B(n25604), .C(n30055), .D(n25615), .Y(n33991)
         );
  AOI22X1 U21326 ( .A(n25625), .B(reg_file[527]), .C(n25636), .D(reg_file[655]), .Y(n33989) );
  AOI22X1 U21327 ( .A(n25647), .B(reg_file[783]), .C(n25658), .D(reg_file[911]), .Y(n33988) );
  NOR2X1 U21328 ( .A(n33993), .B(n33994), .Y(n33979) );
  NAND3X1 U21329 ( .A(n33995), .B(n33996), .C(n33997), .Y(n33994) );
  NOR2X1 U21330 ( .A(n33998), .B(n33999), .Y(n33997) );
  OAI22X1 U21331 ( .A(n30063), .B(n25669), .C(n30064), .D(n25680), .Y(n33999)
         );
  OAI22X1 U21332 ( .A(n30065), .B(n25690), .C(n30066), .D(n25701), .Y(n33998)
         );
  AOI22X1 U21333 ( .A(n25711), .B(reg_file[3471]), .C(n25722), .D(
        reg_file[3343]), .Y(n33996) );
  AOI22X1 U21334 ( .A(n25733), .B(reg_file[3215]), .C(n25744), .D(
        reg_file[3087]), .Y(n33995) );
  NAND3X1 U21335 ( .A(n34000), .B(n34001), .C(n34002), .Y(n33993) );
  NOR2X1 U21336 ( .A(n34003), .B(n34004), .Y(n34002) );
  OAI22X1 U21337 ( .A(n30072), .B(n25755), .C(n30073), .D(n25766), .Y(n34004)
         );
  OAI22X1 U21338 ( .A(n30074), .B(n25776), .C(n30075), .D(n25787), .Y(n34003)
         );
  AOI22X1 U21339 ( .A(n25797), .B(reg_file[2447]), .C(n25808), .D(
        reg_file[2319]), .Y(n34001) );
  AOI22X1 U21340 ( .A(n25819), .B(reg_file[2191]), .C(n25830), .D(
        reg_file[2063]), .Y(n34000) );
  AOI21X1 U21341 ( .A(n34005), .B(n34006), .C(n25486), .Y(rd1data1033_14_) );
  NOR2X1 U21342 ( .A(n34007), .B(n34008), .Y(n34006) );
  NAND3X1 U21343 ( .A(n34009), .B(n34010), .C(n34011), .Y(n34008) );
  NOR2X1 U21344 ( .A(n34012), .B(n34013), .Y(n34011) );
  OAI22X1 U21345 ( .A(n30085), .B(n25497), .C(n30086), .D(n25508), .Y(n34013)
         );
  OAI22X1 U21346 ( .A(n30087), .B(n25518), .C(n30088), .D(n25529), .Y(n34012)
         );
  AOI22X1 U21347 ( .A(n25539), .B(reg_file[1422]), .C(n25550), .D(
        reg_file[1294]), .Y(n34010) );
  AOI22X1 U21348 ( .A(n25561), .B(reg_file[1166]), .C(n25572), .D(
        reg_file[1038]), .Y(n34009) );
  NAND3X1 U21349 ( .A(n34014), .B(n34015), .C(n34016), .Y(n34007) );
  NOR2X1 U21350 ( .A(n34017), .B(n34018), .Y(n34016) );
  OAI22X1 U21351 ( .A(n30094), .B(n25583), .C(n30095), .D(n25594), .Y(n34018)
         );
  OAI22X1 U21352 ( .A(n30096), .B(n25604), .C(n30097), .D(n25615), .Y(n34017)
         );
  AOI22X1 U21353 ( .A(n25625), .B(reg_file[526]), .C(n25636), .D(reg_file[654]), .Y(n34015) );
  AOI22X1 U21354 ( .A(n25647), .B(reg_file[782]), .C(n25658), .D(reg_file[910]), .Y(n34014) );
  NOR2X1 U21355 ( .A(n34019), .B(n34020), .Y(n34005) );
  NAND3X1 U21356 ( .A(n34021), .B(n34022), .C(n34023), .Y(n34020) );
  NOR2X1 U21357 ( .A(n34024), .B(n34025), .Y(n34023) );
  OAI22X1 U21358 ( .A(n30105), .B(n25669), .C(n30106), .D(n25680), .Y(n34025)
         );
  OAI22X1 U21359 ( .A(n30107), .B(n25690), .C(n30108), .D(n25701), .Y(n34024)
         );
  AOI22X1 U21360 ( .A(n25711), .B(reg_file[3470]), .C(n25722), .D(
        reg_file[3342]), .Y(n34022) );
  AOI22X1 U21361 ( .A(n25733), .B(reg_file[3214]), .C(n25744), .D(
        reg_file[3086]), .Y(n34021) );
  NAND3X1 U21362 ( .A(n34026), .B(n34027), .C(n34028), .Y(n34019) );
  NOR2X1 U21363 ( .A(n34029), .B(n34030), .Y(n34028) );
  OAI22X1 U21364 ( .A(n30114), .B(n25755), .C(n30115), .D(n25766), .Y(n34030)
         );
  OAI22X1 U21365 ( .A(n30116), .B(n25776), .C(n30117), .D(n25787), .Y(n34029)
         );
  AOI22X1 U21366 ( .A(n25797), .B(reg_file[2446]), .C(n25808), .D(
        reg_file[2318]), .Y(n34027) );
  AOI22X1 U21367 ( .A(n25819), .B(reg_file[2190]), .C(n25830), .D(
        reg_file[2062]), .Y(n34026) );
  AOI21X1 U21368 ( .A(n34031), .B(n34032), .C(n25486), .Y(rd1data1033_13_) );
  NOR2X1 U21369 ( .A(n34033), .B(n34034), .Y(n34032) );
  NAND3X1 U21370 ( .A(n34035), .B(n34036), .C(n34037), .Y(n34034) );
  NOR2X1 U21371 ( .A(n34038), .B(n34039), .Y(n34037) );
  OAI22X1 U21372 ( .A(n30127), .B(n25497), .C(n30128), .D(n25508), .Y(n34039)
         );
  OAI22X1 U21373 ( .A(n30129), .B(n25518), .C(n30130), .D(n25529), .Y(n34038)
         );
  AOI22X1 U21374 ( .A(n25539), .B(reg_file[1421]), .C(n25550), .D(
        reg_file[1293]), .Y(n34036) );
  AOI22X1 U21375 ( .A(n25561), .B(reg_file[1165]), .C(n25572), .D(
        reg_file[1037]), .Y(n34035) );
  NAND3X1 U21376 ( .A(n34040), .B(n34041), .C(n34042), .Y(n34033) );
  NOR2X1 U21377 ( .A(n34043), .B(n34044), .Y(n34042) );
  OAI22X1 U21378 ( .A(n30136), .B(n25583), .C(n30137), .D(n25594), .Y(n34044)
         );
  OAI22X1 U21379 ( .A(n30138), .B(n25604), .C(n30139), .D(n25615), .Y(n34043)
         );
  AOI22X1 U21380 ( .A(n25625), .B(reg_file[525]), .C(n25636), .D(reg_file[653]), .Y(n34041) );
  AOI22X1 U21381 ( .A(n25647), .B(reg_file[781]), .C(n25658), .D(reg_file[909]), .Y(n34040) );
  NOR2X1 U21382 ( .A(n34045), .B(n34046), .Y(n34031) );
  NAND3X1 U21383 ( .A(n34047), .B(n34048), .C(n34049), .Y(n34046) );
  NOR2X1 U21384 ( .A(n34050), .B(n34051), .Y(n34049) );
  OAI22X1 U21385 ( .A(n30147), .B(n25669), .C(n30148), .D(n25680), .Y(n34051)
         );
  OAI22X1 U21386 ( .A(n30149), .B(n25690), .C(n30150), .D(n25701), .Y(n34050)
         );
  AOI22X1 U21387 ( .A(n25711), .B(reg_file[3469]), .C(n25722), .D(
        reg_file[3341]), .Y(n34048) );
  AOI22X1 U21388 ( .A(n25733), .B(reg_file[3213]), .C(n25744), .D(
        reg_file[3085]), .Y(n34047) );
  NAND3X1 U21389 ( .A(n34052), .B(n34053), .C(n34054), .Y(n34045) );
  NOR2X1 U21390 ( .A(n34055), .B(n34056), .Y(n34054) );
  OAI22X1 U21391 ( .A(n30156), .B(n25755), .C(n30157), .D(n25766), .Y(n34056)
         );
  OAI22X1 U21392 ( .A(n30158), .B(n25776), .C(n30159), .D(n25787), .Y(n34055)
         );
  AOI22X1 U21393 ( .A(n25797), .B(reg_file[2445]), .C(n25808), .D(
        reg_file[2317]), .Y(n34053) );
  AOI22X1 U21394 ( .A(n25819), .B(reg_file[2189]), .C(n25830), .D(
        reg_file[2061]), .Y(n34052) );
  AOI21X1 U21395 ( .A(n34057), .B(n34058), .C(n25486), .Y(rd1data1033_12_) );
  NOR2X1 U21396 ( .A(n34059), .B(n34060), .Y(n34058) );
  NAND3X1 U21397 ( .A(n34061), .B(n34062), .C(n34063), .Y(n34060) );
  NOR2X1 U21398 ( .A(n34064), .B(n34065), .Y(n34063) );
  OAI22X1 U21399 ( .A(n30169), .B(n25497), .C(n30170), .D(n25508), .Y(n34065)
         );
  OAI22X1 U21400 ( .A(n30171), .B(n25518), .C(n30172), .D(n25529), .Y(n34064)
         );
  AOI22X1 U21401 ( .A(n25539), .B(reg_file[1420]), .C(n25550), .D(
        reg_file[1292]), .Y(n34062) );
  AOI22X1 U21402 ( .A(n25561), .B(reg_file[1164]), .C(n25572), .D(
        reg_file[1036]), .Y(n34061) );
  NAND3X1 U21403 ( .A(n34066), .B(n34067), .C(n34068), .Y(n34059) );
  NOR2X1 U21404 ( .A(n34069), .B(n34070), .Y(n34068) );
  OAI22X1 U21405 ( .A(n30178), .B(n25583), .C(n30179), .D(n25594), .Y(n34070)
         );
  OAI22X1 U21406 ( .A(n30180), .B(n25604), .C(n30181), .D(n25615), .Y(n34069)
         );
  AOI22X1 U21407 ( .A(n25625), .B(reg_file[524]), .C(n25636), .D(reg_file[652]), .Y(n34067) );
  AOI22X1 U21408 ( .A(n25647), .B(reg_file[780]), .C(n25658), .D(reg_file[908]), .Y(n34066) );
  NOR2X1 U21409 ( .A(n34071), .B(n34072), .Y(n34057) );
  NAND3X1 U21410 ( .A(n34073), .B(n34074), .C(n34075), .Y(n34072) );
  NOR2X1 U21411 ( .A(n34076), .B(n34077), .Y(n34075) );
  OAI22X1 U21412 ( .A(n30189), .B(n25669), .C(n30190), .D(n25680), .Y(n34077)
         );
  OAI22X1 U21413 ( .A(n30191), .B(n25690), .C(n30192), .D(n25701), .Y(n34076)
         );
  AOI22X1 U21414 ( .A(n25711), .B(reg_file[3468]), .C(n25722), .D(
        reg_file[3340]), .Y(n34074) );
  AOI22X1 U21415 ( .A(n25733), .B(reg_file[3212]), .C(n25744), .D(
        reg_file[3084]), .Y(n34073) );
  NAND3X1 U21416 ( .A(n34078), .B(n34079), .C(n34080), .Y(n34071) );
  NOR2X1 U21417 ( .A(n34081), .B(n34082), .Y(n34080) );
  OAI22X1 U21418 ( .A(n30198), .B(n25755), .C(n30199), .D(n25766), .Y(n34082)
         );
  OAI22X1 U21419 ( .A(n30200), .B(n25776), .C(n30201), .D(n25787), .Y(n34081)
         );
  AOI22X1 U21420 ( .A(n25797), .B(reg_file[2444]), .C(n25808), .D(
        reg_file[2316]), .Y(n34079) );
  AOI22X1 U21421 ( .A(n25819), .B(reg_file[2188]), .C(n25830), .D(
        reg_file[2060]), .Y(n34078) );
  AOI21X1 U21422 ( .A(n34083), .B(n34084), .C(n25486), .Y(rd1data1033_127_) );
  NOR2X1 U21423 ( .A(n34085), .B(n34086), .Y(n34084) );
  NAND3X1 U21424 ( .A(n34087), .B(n34088), .C(n34089), .Y(n34086) );
  NOR2X1 U21425 ( .A(n34090), .B(n34091), .Y(n34089) );
  OAI22X1 U21426 ( .A(n30211), .B(n25497), .C(n30212), .D(n25508), .Y(n34091)
         );
  OAI22X1 U21427 ( .A(n30213), .B(n25518), .C(n30214), .D(n25529), .Y(n34090)
         );
  AOI22X1 U21428 ( .A(n25539), .B(reg_file[1535]), .C(n25550), .D(
        reg_file[1407]), .Y(n34088) );
  AOI22X1 U21429 ( .A(n25561), .B(reg_file[1279]), .C(n25572), .D(
        reg_file[1151]), .Y(n34087) );
  NAND3X1 U21430 ( .A(n34092), .B(n34093), .C(n34094), .Y(n34085) );
  NOR2X1 U21431 ( .A(n34095), .B(n34096), .Y(n34094) );
  OAI22X1 U21432 ( .A(n30220), .B(n25583), .C(n30221), .D(n25594), .Y(n34096)
         );
  OAI22X1 U21433 ( .A(n30222), .B(n25604), .C(n30223), .D(n25615), .Y(n34095)
         );
  AOI22X1 U21434 ( .A(n25625), .B(reg_file[639]), .C(n25636), .D(reg_file[767]), .Y(n34093) );
  AOI22X1 U21435 ( .A(n25647), .B(reg_file[895]), .C(n25658), .D(
        reg_file[1023]), .Y(n34092) );
  NOR2X1 U21436 ( .A(n34097), .B(n34098), .Y(n34083) );
  NAND3X1 U21437 ( .A(n34099), .B(n34100), .C(n34101), .Y(n34098) );
  NOR2X1 U21438 ( .A(n34102), .B(n34103), .Y(n34101) );
  OAI22X1 U21439 ( .A(n30231), .B(n25669), .C(n30232), .D(n25680), .Y(n34103)
         );
  OAI22X1 U21440 ( .A(n30233), .B(n25690), .C(n30234), .D(n25701), .Y(n34102)
         );
  AOI22X1 U21441 ( .A(n25711), .B(reg_file[3583]), .C(n25722), .D(
        reg_file[3455]), .Y(n34100) );
  AOI22X1 U21442 ( .A(n25733), .B(reg_file[3327]), .C(n25744), .D(
        reg_file[3199]), .Y(n34099) );
  NAND3X1 U21443 ( .A(n34104), .B(n34105), .C(n34106), .Y(n34097) );
  NOR2X1 U21444 ( .A(n34107), .B(n34108), .Y(n34106) );
  OAI22X1 U21445 ( .A(n30240), .B(n25755), .C(n30241), .D(n25766), .Y(n34108)
         );
  OAI22X1 U21446 ( .A(n30242), .B(n25776), .C(n30243), .D(n25787), .Y(n34107)
         );
  AOI22X1 U21447 ( .A(n25797), .B(reg_file[2559]), .C(n25808), .D(
        reg_file[2431]), .Y(n34105) );
  AOI22X1 U21448 ( .A(n25819), .B(reg_file[2303]), .C(n25830), .D(
        reg_file[2175]), .Y(n34104) );
  AOI21X1 U21449 ( .A(n34109), .B(n34110), .C(n25486), .Y(rd1data1033_126_) );
  NOR2X1 U21450 ( .A(n34111), .B(n34112), .Y(n34110) );
  NAND3X1 U21451 ( .A(n34113), .B(n34114), .C(n34115), .Y(n34112) );
  NOR2X1 U21452 ( .A(n34116), .B(n34117), .Y(n34115) );
  OAI22X1 U21453 ( .A(n30253), .B(n25497), .C(n30254), .D(n25508), .Y(n34117)
         );
  OAI22X1 U21454 ( .A(n30255), .B(n25518), .C(n30256), .D(n25529), .Y(n34116)
         );
  AOI22X1 U21455 ( .A(n25539), .B(reg_file[1534]), .C(n25550), .D(
        reg_file[1406]), .Y(n34114) );
  AOI22X1 U21456 ( .A(n25561), .B(reg_file[1278]), .C(n25572), .D(
        reg_file[1150]), .Y(n34113) );
  NAND3X1 U21457 ( .A(n34118), .B(n34119), .C(n34120), .Y(n34111) );
  NOR2X1 U21458 ( .A(n34121), .B(n34122), .Y(n34120) );
  OAI22X1 U21459 ( .A(n30262), .B(n25583), .C(n30263), .D(n25594), .Y(n34122)
         );
  OAI22X1 U21460 ( .A(n30264), .B(n25604), .C(n30265), .D(n25615), .Y(n34121)
         );
  AOI22X1 U21461 ( .A(n25625), .B(reg_file[638]), .C(n25636), .D(reg_file[766]), .Y(n34119) );
  AOI22X1 U21462 ( .A(n25647), .B(reg_file[894]), .C(n25658), .D(
        reg_file[1022]), .Y(n34118) );
  NOR2X1 U21463 ( .A(n34123), .B(n34124), .Y(n34109) );
  NAND3X1 U21464 ( .A(n34125), .B(n34126), .C(n34127), .Y(n34124) );
  NOR2X1 U21465 ( .A(n34128), .B(n34129), .Y(n34127) );
  OAI22X1 U21466 ( .A(n30273), .B(n25669), .C(n30274), .D(n25680), .Y(n34129)
         );
  OAI22X1 U21467 ( .A(n30275), .B(n25690), .C(n30276), .D(n25701), .Y(n34128)
         );
  AOI22X1 U21468 ( .A(n25711), .B(reg_file[3582]), .C(n25722), .D(
        reg_file[3454]), .Y(n34126) );
  AOI22X1 U21469 ( .A(n25733), .B(reg_file[3326]), .C(n25744), .D(
        reg_file[3198]), .Y(n34125) );
  NAND3X1 U21470 ( .A(n34130), .B(n34131), .C(n34132), .Y(n34123) );
  NOR2X1 U21471 ( .A(n34133), .B(n34134), .Y(n34132) );
  OAI22X1 U21472 ( .A(n30282), .B(n25755), .C(n30283), .D(n25766), .Y(n34134)
         );
  OAI22X1 U21473 ( .A(n30284), .B(n25776), .C(n30285), .D(n25787), .Y(n34133)
         );
  AOI22X1 U21474 ( .A(n25797), .B(reg_file[2558]), .C(n25808), .D(
        reg_file[2430]), .Y(n34131) );
  AOI22X1 U21475 ( .A(n25819), .B(reg_file[2302]), .C(n25830), .D(
        reg_file[2174]), .Y(n34130) );
  AOI21X1 U21476 ( .A(n34135), .B(n34136), .C(n25486), .Y(rd1data1033_125_) );
  NOR2X1 U21477 ( .A(n34137), .B(n34138), .Y(n34136) );
  NAND3X1 U21478 ( .A(n34139), .B(n34140), .C(n34141), .Y(n34138) );
  NOR2X1 U21479 ( .A(n34142), .B(n34143), .Y(n34141) );
  OAI22X1 U21480 ( .A(n30295), .B(n25497), .C(n30296), .D(n25508), .Y(n34143)
         );
  OAI22X1 U21481 ( .A(n30297), .B(n25518), .C(n30298), .D(n25529), .Y(n34142)
         );
  AOI22X1 U21482 ( .A(n25539), .B(reg_file[1533]), .C(n25550), .D(
        reg_file[1405]), .Y(n34140) );
  AOI22X1 U21483 ( .A(n25561), .B(reg_file[1277]), .C(n25572), .D(
        reg_file[1149]), .Y(n34139) );
  NAND3X1 U21484 ( .A(n34144), .B(n34145), .C(n34146), .Y(n34137) );
  NOR2X1 U21485 ( .A(n34147), .B(n34148), .Y(n34146) );
  OAI22X1 U21486 ( .A(n30304), .B(n25583), .C(n30305), .D(n25594), .Y(n34148)
         );
  OAI22X1 U21487 ( .A(n30306), .B(n25604), .C(n30307), .D(n25615), .Y(n34147)
         );
  AOI22X1 U21488 ( .A(n25625), .B(reg_file[637]), .C(n25636), .D(reg_file[765]), .Y(n34145) );
  AOI22X1 U21489 ( .A(n25647), .B(reg_file[893]), .C(n25658), .D(
        reg_file[1021]), .Y(n34144) );
  NOR2X1 U21490 ( .A(n34149), .B(n34150), .Y(n34135) );
  NAND3X1 U21491 ( .A(n34151), .B(n34152), .C(n34153), .Y(n34150) );
  NOR2X1 U21492 ( .A(n34154), .B(n34155), .Y(n34153) );
  OAI22X1 U21493 ( .A(n30315), .B(n25669), .C(n30316), .D(n25680), .Y(n34155)
         );
  OAI22X1 U21494 ( .A(n30317), .B(n25690), .C(n30318), .D(n25701), .Y(n34154)
         );
  AOI22X1 U21495 ( .A(n25711), .B(reg_file[3581]), .C(n25722), .D(
        reg_file[3453]), .Y(n34152) );
  AOI22X1 U21496 ( .A(n25733), .B(reg_file[3325]), .C(n25744), .D(
        reg_file[3197]), .Y(n34151) );
  NAND3X1 U21497 ( .A(n34156), .B(n34157), .C(n34158), .Y(n34149) );
  NOR2X1 U21498 ( .A(n34159), .B(n34160), .Y(n34158) );
  OAI22X1 U21499 ( .A(n30324), .B(n25755), .C(n30325), .D(n25766), .Y(n34160)
         );
  OAI22X1 U21500 ( .A(n30326), .B(n25776), .C(n30327), .D(n25787), .Y(n34159)
         );
  AOI22X1 U21501 ( .A(n25797), .B(reg_file[2557]), .C(n25808), .D(
        reg_file[2429]), .Y(n34157) );
  AOI22X1 U21502 ( .A(n25819), .B(reg_file[2301]), .C(n25830), .D(
        reg_file[2173]), .Y(n34156) );
  AOI21X1 U21503 ( .A(n34161), .B(n34162), .C(n25486), .Y(rd1data1033_124_) );
  NOR2X1 U21504 ( .A(n34163), .B(n34164), .Y(n34162) );
  NAND3X1 U21505 ( .A(n34165), .B(n34166), .C(n34167), .Y(n34164) );
  NOR2X1 U21506 ( .A(n34168), .B(n34169), .Y(n34167) );
  OAI22X1 U21507 ( .A(n30337), .B(n25497), .C(n30338), .D(n25508), .Y(n34169)
         );
  OAI22X1 U21508 ( .A(n30339), .B(n25518), .C(n30340), .D(n25529), .Y(n34168)
         );
  AOI22X1 U21509 ( .A(n25539), .B(reg_file[1532]), .C(n25550), .D(
        reg_file[1404]), .Y(n34166) );
  AOI22X1 U21510 ( .A(n25561), .B(reg_file[1276]), .C(n25572), .D(
        reg_file[1148]), .Y(n34165) );
  NAND3X1 U21511 ( .A(n34170), .B(n34171), .C(n34172), .Y(n34163) );
  NOR2X1 U21512 ( .A(n34173), .B(n34174), .Y(n34172) );
  OAI22X1 U21513 ( .A(n30346), .B(n25583), .C(n30347), .D(n25594), .Y(n34174)
         );
  OAI22X1 U21514 ( .A(n30348), .B(n25604), .C(n30349), .D(n25615), .Y(n34173)
         );
  AOI22X1 U21515 ( .A(n25625), .B(reg_file[636]), .C(n25636), .D(reg_file[764]), .Y(n34171) );
  AOI22X1 U21516 ( .A(n25647), .B(reg_file[892]), .C(n25658), .D(
        reg_file[1020]), .Y(n34170) );
  NOR2X1 U21517 ( .A(n34175), .B(n34176), .Y(n34161) );
  NAND3X1 U21518 ( .A(n34177), .B(n34178), .C(n34179), .Y(n34176) );
  NOR2X1 U21519 ( .A(n34180), .B(n34181), .Y(n34179) );
  OAI22X1 U21520 ( .A(n30357), .B(n25669), .C(n30358), .D(n25680), .Y(n34181)
         );
  OAI22X1 U21521 ( .A(n30359), .B(n25690), .C(n30360), .D(n25701), .Y(n34180)
         );
  AOI22X1 U21522 ( .A(n25711), .B(reg_file[3580]), .C(n25722), .D(
        reg_file[3452]), .Y(n34178) );
  AOI22X1 U21523 ( .A(n25733), .B(reg_file[3324]), .C(n25744), .D(
        reg_file[3196]), .Y(n34177) );
  NAND3X1 U21524 ( .A(n34182), .B(n34183), .C(n34184), .Y(n34175) );
  NOR2X1 U21525 ( .A(n34185), .B(n34186), .Y(n34184) );
  OAI22X1 U21526 ( .A(n30366), .B(n25755), .C(n30367), .D(n25766), .Y(n34186)
         );
  OAI22X1 U21527 ( .A(n30368), .B(n25776), .C(n30369), .D(n25787), .Y(n34185)
         );
  AOI22X1 U21528 ( .A(n25797), .B(reg_file[2556]), .C(n25808), .D(
        reg_file[2428]), .Y(n34183) );
  AOI22X1 U21529 ( .A(n25819), .B(reg_file[2300]), .C(n25830), .D(
        reg_file[2172]), .Y(n34182) );
  AOI21X1 U21530 ( .A(n34187), .B(n34188), .C(n25486), .Y(rd1data1033_123_) );
  NOR2X1 U21531 ( .A(n34189), .B(n34190), .Y(n34188) );
  NAND3X1 U21532 ( .A(n34191), .B(n34192), .C(n34193), .Y(n34190) );
  NOR2X1 U21533 ( .A(n34194), .B(n34195), .Y(n34193) );
  OAI22X1 U21534 ( .A(n30379), .B(n25497), .C(n30380), .D(n25508), .Y(n34195)
         );
  OAI22X1 U21535 ( .A(n30381), .B(n25518), .C(n30382), .D(n25529), .Y(n34194)
         );
  AOI22X1 U21536 ( .A(n25539), .B(reg_file[1531]), .C(n25550), .D(
        reg_file[1403]), .Y(n34192) );
  AOI22X1 U21537 ( .A(n25561), .B(reg_file[1275]), .C(n25572), .D(
        reg_file[1147]), .Y(n34191) );
  NAND3X1 U21538 ( .A(n34196), .B(n34197), .C(n34198), .Y(n34189) );
  NOR2X1 U21539 ( .A(n34199), .B(n34200), .Y(n34198) );
  OAI22X1 U21540 ( .A(n30388), .B(n25583), .C(n30389), .D(n25594), .Y(n34200)
         );
  OAI22X1 U21541 ( .A(n30390), .B(n25604), .C(n30391), .D(n25615), .Y(n34199)
         );
  AOI22X1 U21542 ( .A(n25625), .B(reg_file[635]), .C(n25636), .D(reg_file[763]), .Y(n34197) );
  AOI22X1 U21543 ( .A(n25647), .B(reg_file[891]), .C(n25658), .D(
        reg_file[1019]), .Y(n34196) );
  NOR2X1 U21544 ( .A(n34201), .B(n34202), .Y(n34187) );
  NAND3X1 U21545 ( .A(n34203), .B(n34204), .C(n34205), .Y(n34202) );
  NOR2X1 U21546 ( .A(n34206), .B(n34207), .Y(n34205) );
  OAI22X1 U21547 ( .A(n30399), .B(n25669), .C(n30400), .D(n25680), .Y(n34207)
         );
  OAI22X1 U21548 ( .A(n30401), .B(n25690), .C(n30402), .D(n25701), .Y(n34206)
         );
  AOI22X1 U21549 ( .A(n25711), .B(reg_file[3579]), .C(n25722), .D(
        reg_file[3451]), .Y(n34204) );
  AOI22X1 U21550 ( .A(n25733), .B(reg_file[3323]), .C(n25744), .D(
        reg_file[3195]), .Y(n34203) );
  NAND3X1 U21551 ( .A(n34208), .B(n34209), .C(n34210), .Y(n34201) );
  NOR2X1 U21552 ( .A(n34211), .B(n34212), .Y(n34210) );
  OAI22X1 U21553 ( .A(n30408), .B(n25755), .C(n30409), .D(n25766), .Y(n34212)
         );
  OAI22X1 U21554 ( .A(n30410), .B(n25776), .C(n30411), .D(n25787), .Y(n34211)
         );
  AOI22X1 U21555 ( .A(n25797), .B(reg_file[2555]), .C(n25808), .D(
        reg_file[2427]), .Y(n34209) );
  AOI22X1 U21556 ( .A(n25819), .B(reg_file[2299]), .C(n25830), .D(
        reg_file[2171]), .Y(n34208) );
  AOI21X1 U21557 ( .A(n34213), .B(n34214), .C(n25486), .Y(rd1data1033_122_) );
  NOR2X1 U21558 ( .A(n34215), .B(n34216), .Y(n34214) );
  NAND3X1 U21559 ( .A(n34217), .B(n34218), .C(n34219), .Y(n34216) );
  NOR2X1 U21560 ( .A(n34220), .B(n34221), .Y(n34219) );
  OAI22X1 U21561 ( .A(n30421), .B(n25497), .C(n30422), .D(n25507), .Y(n34221)
         );
  OAI22X1 U21562 ( .A(n30423), .B(n25518), .C(n30424), .D(n25528), .Y(n34220)
         );
  AOI22X1 U21563 ( .A(n25539), .B(reg_file[1530]), .C(n25550), .D(
        reg_file[1402]), .Y(n34218) );
  AOI22X1 U21564 ( .A(n25561), .B(reg_file[1274]), .C(n25572), .D(
        reg_file[1146]), .Y(n34217) );
  NAND3X1 U21565 ( .A(n34222), .B(n34223), .C(n34224), .Y(n34215) );
  NOR2X1 U21566 ( .A(n34225), .B(n34226), .Y(n34224) );
  OAI22X1 U21567 ( .A(n30430), .B(n25583), .C(n30431), .D(n25593), .Y(n34226)
         );
  OAI22X1 U21568 ( .A(n30432), .B(n25604), .C(n30433), .D(n25614), .Y(n34225)
         );
  AOI22X1 U21569 ( .A(n25625), .B(reg_file[634]), .C(n25636), .D(reg_file[762]), .Y(n34223) );
  AOI22X1 U21570 ( .A(n25647), .B(reg_file[890]), .C(n25658), .D(
        reg_file[1018]), .Y(n34222) );
  NOR2X1 U21571 ( .A(n34227), .B(n34228), .Y(n34213) );
  NAND3X1 U21572 ( .A(n34229), .B(n34230), .C(n34231), .Y(n34228) );
  NOR2X1 U21573 ( .A(n34232), .B(n34233), .Y(n34231) );
  OAI22X1 U21574 ( .A(n30441), .B(n25669), .C(n30442), .D(n25679), .Y(n34233)
         );
  OAI22X1 U21575 ( .A(n30443), .B(n25690), .C(n30444), .D(n25700), .Y(n34232)
         );
  AOI22X1 U21576 ( .A(n25711), .B(reg_file[3578]), .C(n25722), .D(
        reg_file[3450]), .Y(n34230) );
  AOI22X1 U21577 ( .A(n25733), .B(reg_file[3322]), .C(n25744), .D(
        reg_file[3194]), .Y(n34229) );
  NAND3X1 U21578 ( .A(n34234), .B(n34235), .C(n34236), .Y(n34227) );
  NOR2X1 U21579 ( .A(n34237), .B(n34238), .Y(n34236) );
  OAI22X1 U21580 ( .A(n30450), .B(n25755), .C(n30451), .D(n25765), .Y(n34238)
         );
  OAI22X1 U21581 ( .A(n30452), .B(n25776), .C(n30453), .D(n25786), .Y(n34237)
         );
  AOI22X1 U21582 ( .A(n25797), .B(reg_file[2554]), .C(n25808), .D(
        reg_file[2426]), .Y(n34235) );
  AOI22X1 U21583 ( .A(n25819), .B(reg_file[2298]), .C(n25830), .D(
        reg_file[2170]), .Y(n34234) );
  AOI21X1 U21584 ( .A(n34239), .B(n34240), .C(n25486), .Y(rd1data1033_121_) );
  NOR2X1 U21585 ( .A(n34241), .B(n34242), .Y(n34240) );
  NAND3X1 U21586 ( .A(n34243), .B(n34244), .C(n34245), .Y(n34242) );
  NOR2X1 U21587 ( .A(n34246), .B(n34247), .Y(n34245) );
  OAI22X1 U21588 ( .A(n30463), .B(n25497), .C(n30464), .D(n25507), .Y(n34247)
         );
  OAI22X1 U21589 ( .A(n30465), .B(n25518), .C(n30466), .D(n25528), .Y(n34246)
         );
  AOI22X1 U21590 ( .A(n25539), .B(reg_file[1529]), .C(n25550), .D(
        reg_file[1401]), .Y(n34244) );
  AOI22X1 U21591 ( .A(n25561), .B(reg_file[1273]), .C(n25572), .D(
        reg_file[1145]), .Y(n34243) );
  NAND3X1 U21592 ( .A(n34248), .B(n34249), .C(n34250), .Y(n34241) );
  NOR2X1 U21593 ( .A(n34251), .B(n34252), .Y(n34250) );
  OAI22X1 U21594 ( .A(n30472), .B(n25583), .C(n30473), .D(n25593), .Y(n34252)
         );
  OAI22X1 U21595 ( .A(n30474), .B(n25604), .C(n30475), .D(n25614), .Y(n34251)
         );
  AOI22X1 U21596 ( .A(n25625), .B(reg_file[633]), .C(n25636), .D(reg_file[761]), .Y(n34249) );
  AOI22X1 U21597 ( .A(n25647), .B(reg_file[889]), .C(n25658), .D(
        reg_file[1017]), .Y(n34248) );
  NOR2X1 U21598 ( .A(n34253), .B(n34254), .Y(n34239) );
  NAND3X1 U21599 ( .A(n34255), .B(n34256), .C(n34257), .Y(n34254) );
  NOR2X1 U21600 ( .A(n34258), .B(n34259), .Y(n34257) );
  OAI22X1 U21601 ( .A(n30483), .B(n25669), .C(n30484), .D(n25679), .Y(n34259)
         );
  OAI22X1 U21602 ( .A(n30485), .B(n25690), .C(n30486), .D(n25700), .Y(n34258)
         );
  AOI22X1 U21603 ( .A(n25711), .B(reg_file[3577]), .C(n25722), .D(
        reg_file[3449]), .Y(n34256) );
  AOI22X1 U21604 ( .A(n25733), .B(reg_file[3321]), .C(n25744), .D(
        reg_file[3193]), .Y(n34255) );
  NAND3X1 U21605 ( .A(n34260), .B(n34261), .C(n34262), .Y(n34253) );
  NOR2X1 U21606 ( .A(n34263), .B(n34264), .Y(n34262) );
  OAI22X1 U21607 ( .A(n30492), .B(n25755), .C(n30493), .D(n25765), .Y(n34264)
         );
  OAI22X1 U21608 ( .A(n30494), .B(n25776), .C(n30495), .D(n25786), .Y(n34263)
         );
  AOI22X1 U21609 ( .A(n25797), .B(reg_file[2553]), .C(n25808), .D(
        reg_file[2425]), .Y(n34261) );
  AOI22X1 U21610 ( .A(n25819), .B(reg_file[2297]), .C(n25830), .D(
        reg_file[2169]), .Y(n34260) );
  AOI21X1 U21611 ( .A(n34265), .B(n34266), .C(n25485), .Y(rd1data1033_120_) );
  NOR2X1 U21612 ( .A(n34267), .B(n34268), .Y(n34266) );
  NAND3X1 U21613 ( .A(n34269), .B(n34270), .C(n34271), .Y(n34268) );
  NOR2X1 U21614 ( .A(n34272), .B(n34273), .Y(n34271) );
  OAI22X1 U21615 ( .A(n30505), .B(n25496), .C(n30506), .D(n25507), .Y(n34273)
         );
  OAI22X1 U21616 ( .A(n30507), .B(n25517), .C(n30508), .D(n25528), .Y(n34272)
         );
  AOI22X1 U21617 ( .A(n25538), .B(reg_file[1528]), .C(n25549), .D(
        reg_file[1400]), .Y(n34270) );
  AOI22X1 U21618 ( .A(n25560), .B(reg_file[1272]), .C(n25571), .D(
        reg_file[1144]), .Y(n34269) );
  NAND3X1 U21619 ( .A(n34274), .B(n34275), .C(n34276), .Y(n34267) );
  NOR2X1 U21620 ( .A(n34277), .B(n34278), .Y(n34276) );
  OAI22X1 U21621 ( .A(n30514), .B(n25582), .C(n30515), .D(n25593), .Y(n34278)
         );
  OAI22X1 U21622 ( .A(n30516), .B(n25603), .C(n30517), .D(n25614), .Y(n34277)
         );
  AOI22X1 U21623 ( .A(n25624), .B(reg_file[632]), .C(n25635), .D(reg_file[760]), .Y(n34275) );
  AOI22X1 U21624 ( .A(n25646), .B(reg_file[888]), .C(n25657), .D(
        reg_file[1016]), .Y(n34274) );
  NOR2X1 U21625 ( .A(n34279), .B(n34280), .Y(n34265) );
  NAND3X1 U21626 ( .A(n34281), .B(n34282), .C(n34283), .Y(n34280) );
  NOR2X1 U21627 ( .A(n34284), .B(n34285), .Y(n34283) );
  OAI22X1 U21628 ( .A(n30525), .B(n25668), .C(n30526), .D(n25679), .Y(n34285)
         );
  OAI22X1 U21629 ( .A(n30527), .B(n25689), .C(n30528), .D(n25700), .Y(n34284)
         );
  AOI22X1 U21630 ( .A(n25710), .B(reg_file[3576]), .C(n25721), .D(
        reg_file[3448]), .Y(n34282) );
  AOI22X1 U21631 ( .A(n25732), .B(reg_file[3320]), .C(n25743), .D(
        reg_file[3192]), .Y(n34281) );
  NAND3X1 U21632 ( .A(n34286), .B(n34287), .C(n34288), .Y(n34279) );
  NOR2X1 U21633 ( .A(n34289), .B(n34290), .Y(n34288) );
  OAI22X1 U21634 ( .A(n30534), .B(n25754), .C(n30535), .D(n25765), .Y(n34290)
         );
  OAI22X1 U21635 ( .A(n30536), .B(n25775), .C(n30537), .D(n25786), .Y(n34289)
         );
  AOI22X1 U21636 ( .A(n25796), .B(reg_file[2552]), .C(n25807), .D(
        reg_file[2424]), .Y(n34287) );
  AOI22X1 U21637 ( .A(n25818), .B(reg_file[2296]), .C(n25829), .D(
        reg_file[2168]), .Y(n34286) );
  AOI21X1 U21638 ( .A(n34291), .B(n34292), .C(n25485), .Y(rd1data1033_11_) );
  NOR2X1 U21639 ( .A(n34293), .B(n34294), .Y(n34292) );
  NAND3X1 U21640 ( .A(n34295), .B(n34296), .C(n34297), .Y(n34294) );
  NOR2X1 U21641 ( .A(n34298), .B(n34299), .Y(n34297) );
  OAI22X1 U21642 ( .A(n30547), .B(n25496), .C(n30548), .D(n25507), .Y(n34299)
         );
  OAI22X1 U21643 ( .A(n30549), .B(n25517), .C(n30550), .D(n25528), .Y(n34298)
         );
  AOI22X1 U21644 ( .A(n25538), .B(reg_file[1419]), .C(n25549), .D(
        reg_file[1291]), .Y(n34296) );
  AOI22X1 U21645 ( .A(n25560), .B(reg_file[1163]), .C(n25571), .D(
        reg_file[1035]), .Y(n34295) );
  NAND3X1 U21646 ( .A(n34300), .B(n34301), .C(n34302), .Y(n34293) );
  NOR2X1 U21647 ( .A(n34303), .B(n34304), .Y(n34302) );
  OAI22X1 U21648 ( .A(n30556), .B(n25582), .C(n30557), .D(n25593), .Y(n34304)
         );
  OAI22X1 U21649 ( .A(n30558), .B(n25603), .C(n30559), .D(n25614), .Y(n34303)
         );
  AOI22X1 U21650 ( .A(n25624), .B(reg_file[523]), .C(n25635), .D(reg_file[651]), .Y(n34301) );
  AOI22X1 U21651 ( .A(n25646), .B(reg_file[779]), .C(n25657), .D(reg_file[907]), .Y(n34300) );
  NOR2X1 U21652 ( .A(n34305), .B(n34306), .Y(n34291) );
  NAND3X1 U21653 ( .A(n34307), .B(n34308), .C(n34309), .Y(n34306) );
  NOR2X1 U21654 ( .A(n34310), .B(n34311), .Y(n34309) );
  OAI22X1 U21655 ( .A(n30567), .B(n25668), .C(n30568), .D(n25679), .Y(n34311)
         );
  OAI22X1 U21656 ( .A(n30569), .B(n25689), .C(n30570), .D(n25700), .Y(n34310)
         );
  AOI22X1 U21657 ( .A(n25710), .B(reg_file[3467]), .C(n25721), .D(
        reg_file[3339]), .Y(n34308) );
  AOI22X1 U21658 ( .A(n25732), .B(reg_file[3211]), .C(n25743), .D(
        reg_file[3083]), .Y(n34307) );
  NAND3X1 U21659 ( .A(n34312), .B(n34313), .C(n34314), .Y(n34305) );
  NOR2X1 U21660 ( .A(n34315), .B(n34316), .Y(n34314) );
  OAI22X1 U21661 ( .A(n30576), .B(n25754), .C(n30577), .D(n25765), .Y(n34316)
         );
  OAI22X1 U21662 ( .A(n30578), .B(n25775), .C(n30579), .D(n25786), .Y(n34315)
         );
  AOI22X1 U21663 ( .A(n25796), .B(reg_file[2443]), .C(n25807), .D(
        reg_file[2315]), .Y(n34313) );
  AOI22X1 U21664 ( .A(n25818), .B(reg_file[2187]), .C(n25829), .D(
        reg_file[2059]), .Y(n34312) );
  AOI21X1 U21665 ( .A(n34317), .B(n34318), .C(n25485), .Y(rd1data1033_119_) );
  NOR2X1 U21666 ( .A(n34319), .B(n34320), .Y(n34318) );
  NAND3X1 U21667 ( .A(n34321), .B(n34322), .C(n34323), .Y(n34320) );
  NOR2X1 U21668 ( .A(n34324), .B(n34325), .Y(n34323) );
  OAI22X1 U21669 ( .A(n30589), .B(n25496), .C(n30590), .D(n25507), .Y(n34325)
         );
  OAI22X1 U21670 ( .A(n30591), .B(n25517), .C(n30592), .D(n25528), .Y(n34324)
         );
  AOI22X1 U21671 ( .A(n25538), .B(reg_file[1527]), .C(n25549), .D(
        reg_file[1399]), .Y(n34322) );
  AOI22X1 U21672 ( .A(n25560), .B(reg_file[1271]), .C(n25571), .D(
        reg_file[1143]), .Y(n34321) );
  NAND3X1 U21673 ( .A(n34326), .B(n34327), .C(n34328), .Y(n34319) );
  NOR2X1 U21674 ( .A(n34329), .B(n34330), .Y(n34328) );
  OAI22X1 U21675 ( .A(n30598), .B(n25582), .C(n30599), .D(n25593), .Y(n34330)
         );
  OAI22X1 U21676 ( .A(n30600), .B(n25603), .C(n30601), .D(n25614), .Y(n34329)
         );
  AOI22X1 U21677 ( .A(n25624), .B(reg_file[631]), .C(n25635), .D(reg_file[759]), .Y(n34327) );
  AOI22X1 U21678 ( .A(n25646), .B(reg_file[887]), .C(n25657), .D(
        reg_file[1015]), .Y(n34326) );
  NOR2X1 U21679 ( .A(n34331), .B(n34332), .Y(n34317) );
  NAND3X1 U21680 ( .A(n34333), .B(n34334), .C(n34335), .Y(n34332) );
  NOR2X1 U21681 ( .A(n34336), .B(n34337), .Y(n34335) );
  OAI22X1 U21682 ( .A(n30609), .B(n25668), .C(n30610), .D(n25679), .Y(n34337)
         );
  OAI22X1 U21683 ( .A(n30611), .B(n25689), .C(n30612), .D(n25700), .Y(n34336)
         );
  AOI22X1 U21684 ( .A(n25710), .B(reg_file[3575]), .C(n25721), .D(
        reg_file[3447]), .Y(n34334) );
  AOI22X1 U21685 ( .A(n25732), .B(reg_file[3319]), .C(n25743), .D(
        reg_file[3191]), .Y(n34333) );
  NAND3X1 U21686 ( .A(n34338), .B(n34339), .C(n34340), .Y(n34331) );
  NOR2X1 U21687 ( .A(n34341), .B(n34342), .Y(n34340) );
  OAI22X1 U21688 ( .A(n30618), .B(n25754), .C(n30619), .D(n25765), .Y(n34342)
         );
  OAI22X1 U21689 ( .A(n30620), .B(n25775), .C(n30621), .D(n25786), .Y(n34341)
         );
  AOI22X1 U21690 ( .A(n25796), .B(reg_file[2551]), .C(n25807), .D(
        reg_file[2423]), .Y(n34339) );
  AOI22X1 U21691 ( .A(n25818), .B(reg_file[2295]), .C(n25829), .D(
        reg_file[2167]), .Y(n34338) );
  AOI21X1 U21692 ( .A(n34343), .B(n34344), .C(n25485), .Y(rd1data1033_118_) );
  NOR2X1 U21693 ( .A(n34345), .B(n34346), .Y(n34344) );
  NAND3X1 U21694 ( .A(n34347), .B(n34348), .C(n34349), .Y(n34346) );
  NOR2X1 U21695 ( .A(n34350), .B(n34351), .Y(n34349) );
  OAI22X1 U21696 ( .A(n30631), .B(n25496), .C(n30632), .D(n25507), .Y(n34351)
         );
  OAI22X1 U21697 ( .A(n30633), .B(n25517), .C(n30634), .D(n25528), .Y(n34350)
         );
  AOI22X1 U21698 ( .A(n25538), .B(reg_file[1526]), .C(n25549), .D(
        reg_file[1398]), .Y(n34348) );
  AOI22X1 U21699 ( .A(n25560), .B(reg_file[1270]), .C(n25571), .D(
        reg_file[1142]), .Y(n34347) );
  NAND3X1 U21700 ( .A(n34352), .B(n34353), .C(n34354), .Y(n34345) );
  NOR2X1 U21701 ( .A(n34355), .B(n34356), .Y(n34354) );
  OAI22X1 U21702 ( .A(n30640), .B(n25582), .C(n30641), .D(n25593), .Y(n34356)
         );
  OAI22X1 U21703 ( .A(n30642), .B(n25603), .C(n30643), .D(n25614), .Y(n34355)
         );
  AOI22X1 U21704 ( .A(n25624), .B(reg_file[630]), .C(n25635), .D(reg_file[758]), .Y(n34353) );
  AOI22X1 U21705 ( .A(n25646), .B(reg_file[886]), .C(n25657), .D(
        reg_file[1014]), .Y(n34352) );
  NOR2X1 U21706 ( .A(n34357), .B(n34358), .Y(n34343) );
  NAND3X1 U21707 ( .A(n34359), .B(n34360), .C(n34361), .Y(n34358) );
  NOR2X1 U21708 ( .A(n34362), .B(n34363), .Y(n34361) );
  OAI22X1 U21709 ( .A(n30651), .B(n25668), .C(n30652), .D(n25679), .Y(n34363)
         );
  OAI22X1 U21710 ( .A(n30653), .B(n25689), .C(n30654), .D(n25700), .Y(n34362)
         );
  AOI22X1 U21711 ( .A(n25710), .B(reg_file[3574]), .C(n25721), .D(
        reg_file[3446]), .Y(n34360) );
  AOI22X1 U21712 ( .A(n25732), .B(reg_file[3318]), .C(n25743), .D(
        reg_file[3190]), .Y(n34359) );
  NAND3X1 U21713 ( .A(n34364), .B(n34365), .C(n34366), .Y(n34357) );
  NOR2X1 U21714 ( .A(n34367), .B(n34368), .Y(n34366) );
  OAI22X1 U21715 ( .A(n30660), .B(n25754), .C(n30661), .D(n25765), .Y(n34368)
         );
  OAI22X1 U21716 ( .A(n30662), .B(n25775), .C(n30663), .D(n25786), .Y(n34367)
         );
  AOI22X1 U21717 ( .A(n25796), .B(reg_file[2550]), .C(n25807), .D(
        reg_file[2422]), .Y(n34365) );
  AOI22X1 U21718 ( .A(n25818), .B(reg_file[2294]), .C(n25829), .D(
        reg_file[2166]), .Y(n34364) );
  AOI21X1 U21719 ( .A(n34369), .B(n34370), .C(n25485), .Y(rd1data1033_117_) );
  NOR2X1 U21720 ( .A(n34371), .B(n34372), .Y(n34370) );
  NAND3X1 U21721 ( .A(n34373), .B(n34374), .C(n34375), .Y(n34372) );
  NOR2X1 U21722 ( .A(n34376), .B(n34377), .Y(n34375) );
  OAI22X1 U21723 ( .A(n30673), .B(n25496), .C(n30674), .D(n25507), .Y(n34377)
         );
  OAI22X1 U21724 ( .A(n30675), .B(n25517), .C(n30676), .D(n25528), .Y(n34376)
         );
  AOI22X1 U21725 ( .A(n25538), .B(reg_file[1525]), .C(n25549), .D(
        reg_file[1397]), .Y(n34374) );
  AOI22X1 U21726 ( .A(n25560), .B(reg_file[1269]), .C(n25571), .D(
        reg_file[1141]), .Y(n34373) );
  NAND3X1 U21727 ( .A(n34378), .B(n34379), .C(n34380), .Y(n34371) );
  NOR2X1 U21728 ( .A(n34381), .B(n34382), .Y(n34380) );
  OAI22X1 U21729 ( .A(n30682), .B(n25582), .C(n30683), .D(n25593), .Y(n34382)
         );
  OAI22X1 U21730 ( .A(n30684), .B(n25603), .C(n30685), .D(n25614), .Y(n34381)
         );
  AOI22X1 U21731 ( .A(n25624), .B(reg_file[629]), .C(n25635), .D(reg_file[757]), .Y(n34379) );
  AOI22X1 U21732 ( .A(n25646), .B(reg_file[885]), .C(n25657), .D(
        reg_file[1013]), .Y(n34378) );
  NOR2X1 U21733 ( .A(n34383), .B(n34384), .Y(n34369) );
  NAND3X1 U21734 ( .A(n34385), .B(n34386), .C(n34387), .Y(n34384) );
  NOR2X1 U21735 ( .A(n34388), .B(n34389), .Y(n34387) );
  OAI22X1 U21736 ( .A(n30693), .B(n25668), .C(n30694), .D(n25679), .Y(n34389)
         );
  OAI22X1 U21737 ( .A(n30695), .B(n25689), .C(n30696), .D(n25700), .Y(n34388)
         );
  AOI22X1 U21738 ( .A(n25710), .B(reg_file[3573]), .C(n25721), .D(
        reg_file[3445]), .Y(n34386) );
  AOI22X1 U21739 ( .A(n25732), .B(reg_file[3317]), .C(n25743), .D(
        reg_file[3189]), .Y(n34385) );
  NAND3X1 U21740 ( .A(n34390), .B(n34391), .C(n34392), .Y(n34383) );
  NOR2X1 U21741 ( .A(n34393), .B(n34394), .Y(n34392) );
  OAI22X1 U21742 ( .A(n30702), .B(n25754), .C(n30703), .D(n25765), .Y(n34394)
         );
  OAI22X1 U21743 ( .A(n30704), .B(n25775), .C(n30705), .D(n25786), .Y(n34393)
         );
  AOI22X1 U21744 ( .A(n25796), .B(reg_file[2549]), .C(n25807), .D(
        reg_file[2421]), .Y(n34391) );
  AOI22X1 U21745 ( .A(n25818), .B(reg_file[2293]), .C(n25829), .D(
        reg_file[2165]), .Y(n34390) );
  AOI21X1 U21746 ( .A(n34395), .B(n34396), .C(n25485), .Y(rd1data1033_116_) );
  NOR2X1 U21747 ( .A(n34397), .B(n34398), .Y(n34396) );
  NAND3X1 U21748 ( .A(n34399), .B(n34400), .C(n34401), .Y(n34398) );
  NOR2X1 U21749 ( .A(n34402), .B(n34403), .Y(n34401) );
  OAI22X1 U21750 ( .A(n30715), .B(n25496), .C(n30716), .D(n25507), .Y(n34403)
         );
  OAI22X1 U21751 ( .A(n30717), .B(n25517), .C(n30718), .D(n25528), .Y(n34402)
         );
  AOI22X1 U21752 ( .A(n25538), .B(reg_file[1524]), .C(n25549), .D(
        reg_file[1396]), .Y(n34400) );
  AOI22X1 U21753 ( .A(n25560), .B(reg_file[1268]), .C(n25571), .D(
        reg_file[1140]), .Y(n34399) );
  NAND3X1 U21754 ( .A(n34404), .B(n34405), .C(n34406), .Y(n34397) );
  NOR2X1 U21755 ( .A(n34407), .B(n34408), .Y(n34406) );
  OAI22X1 U21756 ( .A(n30724), .B(n25582), .C(n30725), .D(n25593), .Y(n34408)
         );
  OAI22X1 U21757 ( .A(n30726), .B(n25603), .C(n30727), .D(n25614), .Y(n34407)
         );
  AOI22X1 U21758 ( .A(n25624), .B(reg_file[628]), .C(n25635), .D(reg_file[756]), .Y(n34405) );
  AOI22X1 U21759 ( .A(n25646), .B(reg_file[884]), .C(n25657), .D(
        reg_file[1012]), .Y(n34404) );
  NOR2X1 U21760 ( .A(n34409), .B(n34410), .Y(n34395) );
  NAND3X1 U21761 ( .A(n34411), .B(n34412), .C(n34413), .Y(n34410) );
  NOR2X1 U21762 ( .A(n34414), .B(n34415), .Y(n34413) );
  OAI22X1 U21763 ( .A(n30735), .B(n25668), .C(n30736), .D(n25679), .Y(n34415)
         );
  OAI22X1 U21764 ( .A(n30737), .B(n25689), .C(n30738), .D(n25700), .Y(n34414)
         );
  AOI22X1 U21765 ( .A(n25710), .B(reg_file[3572]), .C(n25721), .D(
        reg_file[3444]), .Y(n34412) );
  AOI22X1 U21766 ( .A(n25732), .B(reg_file[3316]), .C(n25743), .D(
        reg_file[3188]), .Y(n34411) );
  NAND3X1 U21767 ( .A(n34416), .B(n34417), .C(n34418), .Y(n34409) );
  NOR2X1 U21768 ( .A(n34419), .B(n34420), .Y(n34418) );
  OAI22X1 U21769 ( .A(n30744), .B(n25754), .C(n30745), .D(n25765), .Y(n34420)
         );
  OAI22X1 U21770 ( .A(n30746), .B(n25775), .C(n30747), .D(n25786), .Y(n34419)
         );
  AOI22X1 U21771 ( .A(n25796), .B(reg_file[2548]), .C(n25807), .D(
        reg_file[2420]), .Y(n34417) );
  AOI22X1 U21772 ( .A(n25818), .B(reg_file[2292]), .C(n25829), .D(
        reg_file[2164]), .Y(n34416) );
  AOI21X1 U21773 ( .A(n34421), .B(n34422), .C(n25485), .Y(rd1data1033_115_) );
  NOR2X1 U21774 ( .A(n34423), .B(n34424), .Y(n34422) );
  NAND3X1 U21775 ( .A(n34425), .B(n34426), .C(n34427), .Y(n34424) );
  NOR2X1 U21776 ( .A(n34428), .B(n34429), .Y(n34427) );
  OAI22X1 U21777 ( .A(n30757), .B(n25496), .C(n30758), .D(n25507), .Y(n34429)
         );
  OAI22X1 U21778 ( .A(n30759), .B(n25517), .C(n30760), .D(n25528), .Y(n34428)
         );
  AOI22X1 U21779 ( .A(n25538), .B(reg_file[1523]), .C(n25549), .D(
        reg_file[1395]), .Y(n34426) );
  AOI22X1 U21780 ( .A(n25560), .B(reg_file[1267]), .C(n25571), .D(
        reg_file[1139]), .Y(n34425) );
  NAND3X1 U21781 ( .A(n34430), .B(n34431), .C(n34432), .Y(n34423) );
  NOR2X1 U21782 ( .A(n34433), .B(n34434), .Y(n34432) );
  OAI22X1 U21783 ( .A(n30766), .B(n25582), .C(n30767), .D(n25593), .Y(n34434)
         );
  OAI22X1 U21784 ( .A(n30768), .B(n25603), .C(n30769), .D(n25614), .Y(n34433)
         );
  AOI22X1 U21785 ( .A(n25624), .B(reg_file[627]), .C(n25635), .D(reg_file[755]), .Y(n34431) );
  AOI22X1 U21786 ( .A(n25646), .B(reg_file[883]), .C(n25657), .D(
        reg_file[1011]), .Y(n34430) );
  NOR2X1 U21787 ( .A(n34435), .B(n34436), .Y(n34421) );
  NAND3X1 U21788 ( .A(n34437), .B(n34438), .C(n34439), .Y(n34436) );
  NOR2X1 U21789 ( .A(n34440), .B(n34441), .Y(n34439) );
  OAI22X1 U21790 ( .A(n30777), .B(n25668), .C(n30778), .D(n25679), .Y(n34441)
         );
  OAI22X1 U21791 ( .A(n30779), .B(n25689), .C(n30780), .D(n25700), .Y(n34440)
         );
  AOI22X1 U21792 ( .A(n25710), .B(reg_file[3571]), .C(n25721), .D(
        reg_file[3443]), .Y(n34438) );
  AOI22X1 U21793 ( .A(n25732), .B(reg_file[3315]), .C(n25743), .D(
        reg_file[3187]), .Y(n34437) );
  NAND3X1 U21794 ( .A(n34442), .B(n34443), .C(n34444), .Y(n34435) );
  NOR2X1 U21795 ( .A(n34445), .B(n34446), .Y(n34444) );
  OAI22X1 U21796 ( .A(n30786), .B(n25754), .C(n30787), .D(n25765), .Y(n34446)
         );
  OAI22X1 U21797 ( .A(n30788), .B(n25775), .C(n30789), .D(n25786), .Y(n34445)
         );
  AOI22X1 U21798 ( .A(n25796), .B(reg_file[2547]), .C(n25807), .D(
        reg_file[2419]), .Y(n34443) );
  AOI22X1 U21799 ( .A(n25818), .B(reg_file[2291]), .C(n25829), .D(
        reg_file[2163]), .Y(n34442) );
  AOI21X1 U21800 ( .A(n34447), .B(n34448), .C(n25485), .Y(rd1data1033_114_) );
  NOR2X1 U21801 ( .A(n34449), .B(n34450), .Y(n34448) );
  NAND3X1 U21802 ( .A(n34451), .B(n34452), .C(n34453), .Y(n34450) );
  NOR2X1 U21803 ( .A(n34454), .B(n34455), .Y(n34453) );
  OAI22X1 U21804 ( .A(n30799), .B(n25496), .C(n30800), .D(n25507), .Y(n34455)
         );
  OAI22X1 U21805 ( .A(n30801), .B(n25517), .C(n30802), .D(n25528), .Y(n34454)
         );
  AOI22X1 U21806 ( .A(n25538), .B(reg_file[1522]), .C(n25549), .D(
        reg_file[1394]), .Y(n34452) );
  AOI22X1 U21807 ( .A(n25560), .B(reg_file[1266]), .C(n25571), .D(
        reg_file[1138]), .Y(n34451) );
  NAND3X1 U21808 ( .A(n34456), .B(n34457), .C(n34458), .Y(n34449) );
  NOR2X1 U21809 ( .A(n34459), .B(n34460), .Y(n34458) );
  OAI22X1 U21810 ( .A(n30808), .B(n25582), .C(n30809), .D(n25593), .Y(n34460)
         );
  OAI22X1 U21811 ( .A(n30810), .B(n25603), .C(n30811), .D(n25614), .Y(n34459)
         );
  AOI22X1 U21812 ( .A(n25624), .B(reg_file[626]), .C(n25635), .D(reg_file[754]), .Y(n34457) );
  AOI22X1 U21813 ( .A(n25646), .B(reg_file[882]), .C(n25657), .D(
        reg_file[1010]), .Y(n34456) );
  NOR2X1 U21814 ( .A(n34461), .B(n34462), .Y(n34447) );
  NAND3X1 U21815 ( .A(n34463), .B(n34464), .C(n34465), .Y(n34462) );
  NOR2X1 U21816 ( .A(n34466), .B(n34467), .Y(n34465) );
  OAI22X1 U21817 ( .A(n30819), .B(n25668), .C(n30820), .D(n25679), .Y(n34467)
         );
  OAI22X1 U21818 ( .A(n30821), .B(n25689), .C(n30822), .D(n25700), .Y(n34466)
         );
  AOI22X1 U21819 ( .A(n25710), .B(reg_file[3570]), .C(n25721), .D(
        reg_file[3442]), .Y(n34464) );
  AOI22X1 U21820 ( .A(n25732), .B(reg_file[3314]), .C(n25743), .D(
        reg_file[3186]), .Y(n34463) );
  NAND3X1 U21821 ( .A(n34468), .B(n34469), .C(n34470), .Y(n34461) );
  NOR2X1 U21822 ( .A(n34471), .B(n34472), .Y(n34470) );
  OAI22X1 U21823 ( .A(n30828), .B(n25754), .C(n30829), .D(n25765), .Y(n34472)
         );
  OAI22X1 U21824 ( .A(n30830), .B(n25775), .C(n30831), .D(n25786), .Y(n34471)
         );
  AOI22X1 U21825 ( .A(n25796), .B(reg_file[2546]), .C(n25807), .D(
        reg_file[2418]), .Y(n34469) );
  AOI22X1 U21826 ( .A(n25818), .B(reg_file[2290]), .C(n25829), .D(
        reg_file[2162]), .Y(n34468) );
  AOI21X1 U21827 ( .A(n34473), .B(n34474), .C(n25485), .Y(rd1data1033_113_) );
  NOR2X1 U21828 ( .A(n34475), .B(n34476), .Y(n34474) );
  NAND3X1 U21829 ( .A(n34477), .B(n34478), .C(n34479), .Y(n34476) );
  NOR2X1 U21830 ( .A(n34480), .B(n34481), .Y(n34479) );
  OAI22X1 U21831 ( .A(n30841), .B(n25496), .C(n30842), .D(n25507), .Y(n34481)
         );
  OAI22X1 U21832 ( .A(n30843), .B(n25517), .C(n30844), .D(n25528), .Y(n34480)
         );
  AOI22X1 U21833 ( .A(n25538), .B(reg_file[1521]), .C(n25549), .D(
        reg_file[1393]), .Y(n34478) );
  AOI22X1 U21834 ( .A(n25560), .B(reg_file[1265]), .C(n25571), .D(
        reg_file[1137]), .Y(n34477) );
  NAND3X1 U21835 ( .A(n34482), .B(n34483), .C(n34484), .Y(n34475) );
  NOR2X1 U21836 ( .A(n34485), .B(n34486), .Y(n34484) );
  OAI22X1 U21837 ( .A(n30850), .B(n25582), .C(n30851), .D(n25593), .Y(n34486)
         );
  OAI22X1 U21838 ( .A(n30852), .B(n25603), .C(n30853), .D(n25614), .Y(n34485)
         );
  AOI22X1 U21839 ( .A(n25624), .B(reg_file[625]), .C(n25635), .D(reg_file[753]), .Y(n34483) );
  AOI22X1 U21840 ( .A(n25646), .B(reg_file[881]), .C(n25657), .D(
        reg_file[1009]), .Y(n34482) );
  NOR2X1 U21841 ( .A(n34487), .B(n34488), .Y(n34473) );
  NAND3X1 U21842 ( .A(n34489), .B(n34490), .C(n34491), .Y(n34488) );
  NOR2X1 U21843 ( .A(n34492), .B(n34493), .Y(n34491) );
  OAI22X1 U21844 ( .A(n30861), .B(n25668), .C(n30862), .D(n25679), .Y(n34493)
         );
  OAI22X1 U21845 ( .A(n30863), .B(n25689), .C(n30864), .D(n25700), .Y(n34492)
         );
  AOI22X1 U21846 ( .A(n25710), .B(reg_file[3569]), .C(n25721), .D(
        reg_file[3441]), .Y(n34490) );
  AOI22X1 U21847 ( .A(n25732), .B(reg_file[3313]), .C(n25743), .D(
        reg_file[3185]), .Y(n34489) );
  NAND3X1 U21848 ( .A(n34494), .B(n34495), .C(n34496), .Y(n34487) );
  NOR2X1 U21849 ( .A(n34497), .B(n34498), .Y(n34496) );
  OAI22X1 U21850 ( .A(n30870), .B(n25754), .C(n30871), .D(n25765), .Y(n34498)
         );
  OAI22X1 U21851 ( .A(n30872), .B(n25775), .C(n30873), .D(n25786), .Y(n34497)
         );
  AOI22X1 U21852 ( .A(n25796), .B(reg_file[2545]), .C(n25807), .D(
        reg_file[2417]), .Y(n34495) );
  AOI22X1 U21853 ( .A(n25818), .B(reg_file[2289]), .C(n25829), .D(
        reg_file[2161]), .Y(n34494) );
  AOI21X1 U21854 ( .A(n34499), .B(n34500), .C(n25485), .Y(rd1data1033_112_) );
  NOR2X1 U21855 ( .A(n34501), .B(n34502), .Y(n34500) );
  NAND3X1 U21856 ( .A(n34503), .B(n34504), .C(n34505), .Y(n34502) );
  NOR2X1 U21857 ( .A(n34506), .B(n34507), .Y(n34505) );
  OAI22X1 U21858 ( .A(n30883), .B(n25496), .C(n30884), .D(n25507), .Y(n34507)
         );
  OAI22X1 U21859 ( .A(n30885), .B(n25517), .C(n30886), .D(n25528), .Y(n34506)
         );
  AOI22X1 U21860 ( .A(n25538), .B(reg_file[1520]), .C(n25549), .D(
        reg_file[1392]), .Y(n34504) );
  AOI22X1 U21861 ( .A(n25560), .B(reg_file[1264]), .C(n25571), .D(
        reg_file[1136]), .Y(n34503) );
  NAND3X1 U21862 ( .A(n34508), .B(n34509), .C(n34510), .Y(n34501) );
  NOR2X1 U21863 ( .A(n34511), .B(n34512), .Y(n34510) );
  OAI22X1 U21864 ( .A(n30892), .B(n25582), .C(n30893), .D(n25593), .Y(n34512)
         );
  OAI22X1 U21865 ( .A(n30894), .B(n25603), .C(n30895), .D(n25614), .Y(n34511)
         );
  AOI22X1 U21866 ( .A(n25624), .B(reg_file[624]), .C(n25635), .D(reg_file[752]), .Y(n34509) );
  AOI22X1 U21867 ( .A(n25646), .B(reg_file[880]), .C(n25657), .D(
        reg_file[1008]), .Y(n34508) );
  NOR2X1 U21868 ( .A(n34513), .B(n34514), .Y(n34499) );
  NAND3X1 U21869 ( .A(n34515), .B(n34516), .C(n34517), .Y(n34514) );
  NOR2X1 U21870 ( .A(n34518), .B(n34519), .Y(n34517) );
  OAI22X1 U21871 ( .A(n30903), .B(n25668), .C(n30904), .D(n25679), .Y(n34519)
         );
  OAI22X1 U21872 ( .A(n30905), .B(n25689), .C(n30906), .D(n25700), .Y(n34518)
         );
  AOI22X1 U21873 ( .A(n25710), .B(reg_file[3568]), .C(n25721), .D(
        reg_file[3440]), .Y(n34516) );
  AOI22X1 U21874 ( .A(n25732), .B(reg_file[3312]), .C(n25743), .D(
        reg_file[3184]), .Y(n34515) );
  NAND3X1 U21875 ( .A(n34520), .B(n34521), .C(n34522), .Y(n34513) );
  NOR2X1 U21876 ( .A(n34523), .B(n34524), .Y(n34522) );
  OAI22X1 U21877 ( .A(n30912), .B(n25754), .C(n30913), .D(n25765), .Y(n34524)
         );
  OAI22X1 U21878 ( .A(n30914), .B(n25775), .C(n30915), .D(n25786), .Y(n34523)
         );
  AOI22X1 U21879 ( .A(n25796), .B(reg_file[2544]), .C(n25807), .D(
        reg_file[2416]), .Y(n34521) );
  AOI22X1 U21880 ( .A(n25818), .B(reg_file[2288]), .C(n25829), .D(
        reg_file[2160]), .Y(n34520) );
  AOI21X1 U21881 ( .A(n34525), .B(n34526), .C(n25485), .Y(rd1data1033_111_) );
  NOR2X1 U21882 ( .A(n34527), .B(n34528), .Y(n34526) );
  NAND3X1 U21883 ( .A(n34529), .B(n34530), .C(n34531), .Y(n34528) );
  NOR2X1 U21884 ( .A(n34532), .B(n34533), .Y(n34531) );
  OAI22X1 U21885 ( .A(n30925), .B(n25496), .C(n30926), .D(n25507), .Y(n34533)
         );
  OAI22X1 U21886 ( .A(n30927), .B(n25517), .C(n30928), .D(n25528), .Y(n34532)
         );
  AOI22X1 U21887 ( .A(n25538), .B(reg_file[1519]), .C(n25549), .D(
        reg_file[1391]), .Y(n34530) );
  AOI22X1 U21888 ( .A(n25560), .B(reg_file[1263]), .C(n25571), .D(
        reg_file[1135]), .Y(n34529) );
  NAND3X1 U21889 ( .A(n34534), .B(n34535), .C(n34536), .Y(n34527) );
  NOR2X1 U21890 ( .A(n34537), .B(n34538), .Y(n34536) );
  OAI22X1 U21891 ( .A(n30934), .B(n25582), .C(n30935), .D(n25593), .Y(n34538)
         );
  OAI22X1 U21892 ( .A(n30936), .B(n25603), .C(n30937), .D(n25614), .Y(n34537)
         );
  AOI22X1 U21893 ( .A(n25624), .B(reg_file[623]), .C(n25635), .D(reg_file[751]), .Y(n34535) );
  AOI22X1 U21894 ( .A(n25646), .B(reg_file[879]), .C(n25657), .D(
        reg_file[1007]), .Y(n34534) );
  NOR2X1 U21895 ( .A(n34539), .B(n34540), .Y(n34525) );
  NAND3X1 U21896 ( .A(n34541), .B(n34542), .C(n34543), .Y(n34540) );
  NOR2X1 U21897 ( .A(n34544), .B(n34545), .Y(n34543) );
  OAI22X1 U21898 ( .A(n30945), .B(n25668), .C(n30946), .D(n25679), .Y(n34545)
         );
  OAI22X1 U21899 ( .A(n30947), .B(n25689), .C(n30948), .D(n25700), .Y(n34544)
         );
  AOI22X1 U21900 ( .A(n25710), .B(reg_file[3567]), .C(n25721), .D(
        reg_file[3439]), .Y(n34542) );
  AOI22X1 U21901 ( .A(n25732), .B(reg_file[3311]), .C(n25743), .D(
        reg_file[3183]), .Y(n34541) );
  NAND3X1 U21902 ( .A(n34546), .B(n34547), .C(n34548), .Y(n34539) );
  NOR2X1 U21903 ( .A(n34549), .B(n34550), .Y(n34548) );
  OAI22X1 U21904 ( .A(n30954), .B(n25754), .C(n30955), .D(n25765), .Y(n34550)
         );
  OAI22X1 U21905 ( .A(n30956), .B(n25775), .C(n30957), .D(n25786), .Y(n34549)
         );
  AOI22X1 U21906 ( .A(n25796), .B(reg_file[2543]), .C(n25807), .D(
        reg_file[2415]), .Y(n34547) );
  AOI22X1 U21907 ( .A(n25818), .B(reg_file[2287]), .C(n25829), .D(
        reg_file[2159]), .Y(n34546) );
  AOI21X1 U21908 ( .A(n34551), .B(n34552), .C(n25485), .Y(rd1data1033_110_) );
  NOR2X1 U21909 ( .A(n34553), .B(n34554), .Y(n34552) );
  NAND3X1 U21910 ( .A(n34555), .B(n34556), .C(n34557), .Y(n34554) );
  NOR2X1 U21911 ( .A(n34558), .B(n34559), .Y(n34557) );
  OAI22X1 U21912 ( .A(n30967), .B(n25496), .C(n30968), .D(n25506), .Y(n34559)
         );
  OAI22X1 U21913 ( .A(n30969), .B(n25517), .C(n30970), .D(n25527), .Y(n34558)
         );
  AOI22X1 U21914 ( .A(n25538), .B(reg_file[1518]), .C(n25549), .D(
        reg_file[1390]), .Y(n34556) );
  AOI22X1 U21915 ( .A(n25560), .B(reg_file[1262]), .C(n25571), .D(
        reg_file[1134]), .Y(n34555) );
  NAND3X1 U21916 ( .A(n34560), .B(n34561), .C(n34562), .Y(n34553) );
  NOR2X1 U21917 ( .A(n34563), .B(n34564), .Y(n34562) );
  OAI22X1 U21918 ( .A(n30976), .B(n25582), .C(n30977), .D(n25592), .Y(n34564)
         );
  OAI22X1 U21919 ( .A(n30978), .B(n25603), .C(n30979), .D(n25613), .Y(n34563)
         );
  AOI22X1 U21920 ( .A(n25624), .B(reg_file[622]), .C(n25635), .D(reg_file[750]), .Y(n34561) );
  AOI22X1 U21921 ( .A(n25646), .B(reg_file[878]), .C(n25657), .D(
        reg_file[1006]), .Y(n34560) );
  NOR2X1 U21922 ( .A(n34565), .B(n34566), .Y(n34551) );
  NAND3X1 U21923 ( .A(n34567), .B(n34568), .C(n34569), .Y(n34566) );
  NOR2X1 U21924 ( .A(n34570), .B(n34571), .Y(n34569) );
  OAI22X1 U21925 ( .A(n30987), .B(n25668), .C(n30988), .D(n25678), .Y(n34571)
         );
  OAI22X1 U21926 ( .A(n30989), .B(n25689), .C(n30990), .D(n25699), .Y(n34570)
         );
  AOI22X1 U21927 ( .A(n25710), .B(reg_file[3566]), .C(n25721), .D(
        reg_file[3438]), .Y(n34568) );
  AOI22X1 U21928 ( .A(n25732), .B(reg_file[3310]), .C(n25743), .D(
        reg_file[3182]), .Y(n34567) );
  NAND3X1 U21929 ( .A(n34572), .B(n34573), .C(n34574), .Y(n34565) );
  NOR2X1 U21930 ( .A(n34575), .B(n34576), .Y(n34574) );
  OAI22X1 U21931 ( .A(n30996), .B(n25754), .C(n30997), .D(n25764), .Y(n34576)
         );
  OAI22X1 U21932 ( .A(n30998), .B(n25775), .C(n30999), .D(n25785), .Y(n34575)
         );
  AOI22X1 U21933 ( .A(n25796), .B(reg_file[2542]), .C(n25807), .D(
        reg_file[2414]), .Y(n34573) );
  AOI22X1 U21934 ( .A(n25818), .B(reg_file[2286]), .C(n25829), .D(
        reg_file[2158]), .Y(n34572) );
  AOI21X1 U21935 ( .A(n34577), .B(n34578), .C(n25484), .Y(rd1data1033_10_) );
  NOR2X1 U21936 ( .A(n34579), .B(n34580), .Y(n34578) );
  NAND3X1 U21937 ( .A(n34581), .B(n34582), .C(n34583), .Y(n34580) );
  NOR2X1 U21938 ( .A(n34584), .B(n34585), .Y(n34583) );
  OAI22X1 U21939 ( .A(n31009), .B(n25495), .C(n31010), .D(n25506), .Y(n34585)
         );
  OAI22X1 U21940 ( .A(n31011), .B(n25516), .C(n31012), .D(n25527), .Y(n34584)
         );
  AOI22X1 U21941 ( .A(n25537), .B(reg_file[1418]), .C(n25548), .D(
        reg_file[1290]), .Y(n34582) );
  AOI22X1 U21942 ( .A(n25559), .B(reg_file[1162]), .C(n25570), .D(
        reg_file[1034]), .Y(n34581) );
  NAND3X1 U21943 ( .A(n34586), .B(n34587), .C(n34588), .Y(n34579) );
  NOR2X1 U21944 ( .A(n34589), .B(n34590), .Y(n34588) );
  OAI22X1 U21945 ( .A(n31018), .B(n25581), .C(n31019), .D(n25592), .Y(n34590)
         );
  OAI22X1 U21946 ( .A(n31020), .B(n25602), .C(n31021), .D(n25613), .Y(n34589)
         );
  AOI22X1 U21947 ( .A(n25623), .B(reg_file[522]), .C(n25634), .D(reg_file[650]), .Y(n34587) );
  AOI22X1 U21948 ( .A(n25645), .B(reg_file[778]), .C(n25656), .D(reg_file[906]), .Y(n34586) );
  NOR2X1 U21949 ( .A(n34591), .B(n34592), .Y(n34577) );
  NAND3X1 U21950 ( .A(n34593), .B(n34594), .C(n34595), .Y(n34592) );
  NOR2X1 U21951 ( .A(n34596), .B(n34597), .Y(n34595) );
  OAI22X1 U21952 ( .A(n31029), .B(n25667), .C(n31030), .D(n25678), .Y(n34597)
         );
  OAI22X1 U21953 ( .A(n31031), .B(n25688), .C(n31032), .D(n25699), .Y(n34596)
         );
  AOI22X1 U21954 ( .A(n25709), .B(reg_file[3466]), .C(n25720), .D(
        reg_file[3338]), .Y(n34594) );
  AOI22X1 U21955 ( .A(n25731), .B(reg_file[3210]), .C(n25742), .D(
        reg_file[3082]), .Y(n34593) );
  NAND3X1 U21956 ( .A(n34598), .B(n34599), .C(n34600), .Y(n34591) );
  NOR2X1 U21957 ( .A(n34601), .B(n34602), .Y(n34600) );
  OAI22X1 U21958 ( .A(n31038), .B(n25753), .C(n31039), .D(n25764), .Y(n34602)
         );
  OAI22X1 U21959 ( .A(n31040), .B(n25774), .C(n31041), .D(n25785), .Y(n34601)
         );
  AOI22X1 U21960 ( .A(n25795), .B(reg_file[2442]), .C(n25806), .D(
        reg_file[2314]), .Y(n34599) );
  AOI22X1 U21961 ( .A(n25817), .B(reg_file[2186]), .C(n25828), .D(
        reg_file[2058]), .Y(n34598) );
  AOI21X1 U21962 ( .A(n34603), .B(n34604), .C(n25484), .Y(rd1data1033_109_) );
  NOR2X1 U21963 ( .A(n34605), .B(n34606), .Y(n34604) );
  NAND3X1 U21964 ( .A(n34607), .B(n34608), .C(n34609), .Y(n34606) );
  NOR2X1 U21965 ( .A(n34610), .B(n34611), .Y(n34609) );
  OAI22X1 U21966 ( .A(n31051), .B(n25495), .C(n31052), .D(n25506), .Y(n34611)
         );
  OAI22X1 U21967 ( .A(n31053), .B(n25516), .C(n31054), .D(n25527), .Y(n34610)
         );
  AOI22X1 U21968 ( .A(n25537), .B(reg_file[1517]), .C(n25548), .D(
        reg_file[1389]), .Y(n34608) );
  AOI22X1 U21969 ( .A(n25559), .B(reg_file[1261]), .C(n25570), .D(
        reg_file[1133]), .Y(n34607) );
  NAND3X1 U21970 ( .A(n34612), .B(n34613), .C(n34614), .Y(n34605) );
  NOR2X1 U21971 ( .A(n34615), .B(n34616), .Y(n34614) );
  OAI22X1 U21972 ( .A(n31060), .B(n25581), .C(n31061), .D(n25592), .Y(n34616)
         );
  OAI22X1 U21973 ( .A(n31062), .B(n25602), .C(n31063), .D(n25613), .Y(n34615)
         );
  AOI22X1 U21974 ( .A(n25623), .B(reg_file[621]), .C(n25634), .D(reg_file[749]), .Y(n34613) );
  AOI22X1 U21975 ( .A(n25645), .B(reg_file[877]), .C(n25656), .D(
        reg_file[1005]), .Y(n34612) );
  NOR2X1 U21976 ( .A(n34617), .B(n34618), .Y(n34603) );
  NAND3X1 U21977 ( .A(n34619), .B(n34620), .C(n34621), .Y(n34618) );
  NOR2X1 U21978 ( .A(n34622), .B(n34623), .Y(n34621) );
  OAI22X1 U21979 ( .A(n31071), .B(n25667), .C(n31072), .D(n25678), .Y(n34623)
         );
  OAI22X1 U21980 ( .A(n31073), .B(n25688), .C(n31074), .D(n25699), .Y(n34622)
         );
  AOI22X1 U21981 ( .A(n25709), .B(reg_file[3565]), .C(n25720), .D(
        reg_file[3437]), .Y(n34620) );
  AOI22X1 U21982 ( .A(n25731), .B(reg_file[3309]), .C(n25742), .D(
        reg_file[3181]), .Y(n34619) );
  NAND3X1 U21983 ( .A(n34624), .B(n34625), .C(n34626), .Y(n34617) );
  NOR2X1 U21984 ( .A(n34627), .B(n34628), .Y(n34626) );
  OAI22X1 U21985 ( .A(n31080), .B(n25753), .C(n31081), .D(n25764), .Y(n34628)
         );
  OAI22X1 U21986 ( .A(n31082), .B(n25774), .C(n31083), .D(n25785), .Y(n34627)
         );
  AOI22X1 U21987 ( .A(n25795), .B(reg_file[2541]), .C(n25806), .D(
        reg_file[2413]), .Y(n34625) );
  AOI22X1 U21988 ( .A(n25817), .B(reg_file[2285]), .C(n25828), .D(
        reg_file[2157]), .Y(n34624) );
  AOI21X1 U21989 ( .A(n34629), .B(n34630), .C(n25484), .Y(rd1data1033_108_) );
  NOR2X1 U21990 ( .A(n34631), .B(n34632), .Y(n34630) );
  NAND3X1 U21991 ( .A(n34633), .B(n34634), .C(n34635), .Y(n34632) );
  NOR2X1 U21992 ( .A(n34636), .B(n34637), .Y(n34635) );
  OAI22X1 U21993 ( .A(n31093), .B(n25495), .C(n31094), .D(n25506), .Y(n34637)
         );
  OAI22X1 U21994 ( .A(n31095), .B(n25516), .C(n31096), .D(n25527), .Y(n34636)
         );
  AOI22X1 U21995 ( .A(n25537), .B(reg_file[1516]), .C(n25548), .D(
        reg_file[1388]), .Y(n34634) );
  AOI22X1 U21996 ( .A(n25559), .B(reg_file[1260]), .C(n25570), .D(
        reg_file[1132]), .Y(n34633) );
  NAND3X1 U21997 ( .A(n34638), .B(n34639), .C(n34640), .Y(n34631) );
  NOR2X1 U21998 ( .A(n34641), .B(n34642), .Y(n34640) );
  OAI22X1 U21999 ( .A(n31102), .B(n25581), .C(n31103), .D(n25592), .Y(n34642)
         );
  OAI22X1 U22000 ( .A(n31104), .B(n25602), .C(n31105), .D(n25613), .Y(n34641)
         );
  AOI22X1 U22001 ( .A(n25623), .B(reg_file[620]), .C(n25634), .D(reg_file[748]), .Y(n34639) );
  AOI22X1 U22002 ( .A(n25645), .B(reg_file[876]), .C(n25656), .D(
        reg_file[1004]), .Y(n34638) );
  NOR2X1 U22003 ( .A(n34643), .B(n34644), .Y(n34629) );
  NAND3X1 U22004 ( .A(n34645), .B(n34646), .C(n34647), .Y(n34644) );
  NOR2X1 U22005 ( .A(n34648), .B(n34649), .Y(n34647) );
  OAI22X1 U22006 ( .A(n31113), .B(n25667), .C(n31114), .D(n25678), .Y(n34649)
         );
  OAI22X1 U22007 ( .A(n31115), .B(n25688), .C(n31116), .D(n25699), .Y(n34648)
         );
  AOI22X1 U22008 ( .A(n25709), .B(reg_file[3564]), .C(n25720), .D(
        reg_file[3436]), .Y(n34646) );
  AOI22X1 U22009 ( .A(n25731), .B(reg_file[3308]), .C(n25742), .D(
        reg_file[3180]), .Y(n34645) );
  NAND3X1 U22010 ( .A(n34650), .B(n34651), .C(n34652), .Y(n34643) );
  NOR2X1 U22011 ( .A(n34653), .B(n34654), .Y(n34652) );
  OAI22X1 U22012 ( .A(n31122), .B(n25753), .C(n31123), .D(n25764), .Y(n34654)
         );
  OAI22X1 U22013 ( .A(n31124), .B(n25774), .C(n31125), .D(n25785), .Y(n34653)
         );
  AOI22X1 U22014 ( .A(n25795), .B(reg_file[2540]), .C(n25806), .D(
        reg_file[2412]), .Y(n34651) );
  AOI22X1 U22015 ( .A(n25817), .B(reg_file[2284]), .C(n25828), .D(
        reg_file[2156]), .Y(n34650) );
  AOI21X1 U22016 ( .A(n34655), .B(n34656), .C(n25484), .Y(rd1data1033_107_) );
  NOR2X1 U22017 ( .A(n34657), .B(n34658), .Y(n34656) );
  NAND3X1 U22018 ( .A(n34659), .B(n34660), .C(n34661), .Y(n34658) );
  NOR2X1 U22019 ( .A(n34662), .B(n34663), .Y(n34661) );
  OAI22X1 U22020 ( .A(n31135), .B(n25495), .C(n31136), .D(n25506), .Y(n34663)
         );
  OAI22X1 U22021 ( .A(n31137), .B(n25516), .C(n31138), .D(n25527), .Y(n34662)
         );
  AOI22X1 U22022 ( .A(n25537), .B(reg_file[1515]), .C(n25548), .D(
        reg_file[1387]), .Y(n34660) );
  AOI22X1 U22023 ( .A(n25559), .B(reg_file[1259]), .C(n25570), .D(
        reg_file[1131]), .Y(n34659) );
  NAND3X1 U22024 ( .A(n34664), .B(n34665), .C(n34666), .Y(n34657) );
  NOR2X1 U22025 ( .A(n34667), .B(n34668), .Y(n34666) );
  OAI22X1 U22026 ( .A(n31144), .B(n25581), .C(n31145), .D(n25592), .Y(n34668)
         );
  OAI22X1 U22027 ( .A(n31146), .B(n25602), .C(n31147), .D(n25613), .Y(n34667)
         );
  AOI22X1 U22028 ( .A(n25623), .B(reg_file[619]), .C(n25634), .D(reg_file[747]), .Y(n34665) );
  AOI22X1 U22029 ( .A(n25645), .B(reg_file[875]), .C(n25656), .D(
        reg_file[1003]), .Y(n34664) );
  NOR2X1 U22030 ( .A(n34669), .B(n34670), .Y(n34655) );
  NAND3X1 U22031 ( .A(n34671), .B(n34672), .C(n34673), .Y(n34670) );
  NOR2X1 U22032 ( .A(n34674), .B(n34675), .Y(n34673) );
  OAI22X1 U22033 ( .A(n31155), .B(n25667), .C(n31156), .D(n25678), .Y(n34675)
         );
  OAI22X1 U22034 ( .A(n31157), .B(n25688), .C(n31158), .D(n25699), .Y(n34674)
         );
  AOI22X1 U22035 ( .A(n25709), .B(reg_file[3563]), .C(n25720), .D(
        reg_file[3435]), .Y(n34672) );
  AOI22X1 U22036 ( .A(n25731), .B(reg_file[3307]), .C(n25742), .D(
        reg_file[3179]), .Y(n34671) );
  NAND3X1 U22037 ( .A(n34676), .B(n34677), .C(n34678), .Y(n34669) );
  NOR2X1 U22038 ( .A(n34679), .B(n34680), .Y(n34678) );
  OAI22X1 U22039 ( .A(n31164), .B(n25753), .C(n31165), .D(n25764), .Y(n34680)
         );
  OAI22X1 U22040 ( .A(n31166), .B(n25774), .C(n31167), .D(n25785), .Y(n34679)
         );
  AOI22X1 U22041 ( .A(n25795), .B(reg_file[2539]), .C(n25806), .D(
        reg_file[2411]), .Y(n34677) );
  AOI22X1 U22042 ( .A(n25817), .B(reg_file[2283]), .C(n25828), .D(
        reg_file[2155]), .Y(n34676) );
  AOI21X1 U22043 ( .A(n34681), .B(n34682), .C(n25484), .Y(rd1data1033_106_) );
  NOR2X1 U22044 ( .A(n34683), .B(n34684), .Y(n34682) );
  NAND3X1 U22045 ( .A(n34685), .B(n34686), .C(n34687), .Y(n34684) );
  NOR2X1 U22046 ( .A(n34688), .B(n34689), .Y(n34687) );
  OAI22X1 U22047 ( .A(n31177), .B(n25495), .C(n31178), .D(n25506), .Y(n34689)
         );
  OAI22X1 U22048 ( .A(n31179), .B(n25516), .C(n31180), .D(n25527), .Y(n34688)
         );
  AOI22X1 U22049 ( .A(n25537), .B(reg_file[1514]), .C(n25548), .D(
        reg_file[1386]), .Y(n34686) );
  AOI22X1 U22050 ( .A(n25559), .B(reg_file[1258]), .C(n25570), .D(
        reg_file[1130]), .Y(n34685) );
  NAND3X1 U22051 ( .A(n34690), .B(n34691), .C(n34692), .Y(n34683) );
  NOR2X1 U22052 ( .A(n34693), .B(n34694), .Y(n34692) );
  OAI22X1 U22053 ( .A(n31186), .B(n25581), .C(n31187), .D(n25592), .Y(n34694)
         );
  OAI22X1 U22054 ( .A(n31188), .B(n25602), .C(n31189), .D(n25613), .Y(n34693)
         );
  AOI22X1 U22055 ( .A(n25623), .B(reg_file[618]), .C(n25634), .D(reg_file[746]), .Y(n34691) );
  AOI22X1 U22056 ( .A(n25645), .B(reg_file[874]), .C(n25656), .D(
        reg_file[1002]), .Y(n34690) );
  NOR2X1 U22057 ( .A(n34695), .B(n34696), .Y(n34681) );
  NAND3X1 U22058 ( .A(n34697), .B(n34698), .C(n34699), .Y(n34696) );
  NOR2X1 U22059 ( .A(n34700), .B(n34701), .Y(n34699) );
  OAI22X1 U22060 ( .A(n31197), .B(n25667), .C(n31198), .D(n25678), .Y(n34701)
         );
  OAI22X1 U22061 ( .A(n31199), .B(n25688), .C(n31200), .D(n25699), .Y(n34700)
         );
  AOI22X1 U22062 ( .A(n25709), .B(reg_file[3562]), .C(n25720), .D(
        reg_file[3434]), .Y(n34698) );
  AOI22X1 U22063 ( .A(n25731), .B(reg_file[3306]), .C(n25742), .D(
        reg_file[3178]), .Y(n34697) );
  NAND3X1 U22064 ( .A(n34702), .B(n34703), .C(n34704), .Y(n34695) );
  NOR2X1 U22065 ( .A(n34705), .B(n34706), .Y(n34704) );
  OAI22X1 U22066 ( .A(n31206), .B(n25753), .C(n31207), .D(n25764), .Y(n34706)
         );
  OAI22X1 U22067 ( .A(n31208), .B(n25774), .C(n31209), .D(n25785), .Y(n34705)
         );
  AOI22X1 U22068 ( .A(n25795), .B(reg_file[2538]), .C(n25806), .D(
        reg_file[2410]), .Y(n34703) );
  AOI22X1 U22069 ( .A(n25817), .B(reg_file[2282]), .C(n25828), .D(
        reg_file[2154]), .Y(n34702) );
  AOI21X1 U22070 ( .A(n34707), .B(n34708), .C(n25484), .Y(rd1data1033_105_) );
  NOR2X1 U22071 ( .A(n34709), .B(n34710), .Y(n34708) );
  NAND3X1 U22072 ( .A(n34711), .B(n34712), .C(n34713), .Y(n34710) );
  NOR2X1 U22073 ( .A(n34714), .B(n34715), .Y(n34713) );
  OAI22X1 U22074 ( .A(n31219), .B(n25495), .C(n31220), .D(n25506), .Y(n34715)
         );
  OAI22X1 U22075 ( .A(n31221), .B(n25516), .C(n31222), .D(n25527), .Y(n34714)
         );
  AOI22X1 U22076 ( .A(n25537), .B(reg_file[1513]), .C(n25548), .D(
        reg_file[1385]), .Y(n34712) );
  AOI22X1 U22077 ( .A(n25559), .B(reg_file[1257]), .C(n25570), .D(
        reg_file[1129]), .Y(n34711) );
  NAND3X1 U22078 ( .A(n34716), .B(n34717), .C(n34718), .Y(n34709) );
  NOR2X1 U22079 ( .A(n34719), .B(n34720), .Y(n34718) );
  OAI22X1 U22080 ( .A(n31228), .B(n25581), .C(n31229), .D(n25592), .Y(n34720)
         );
  OAI22X1 U22081 ( .A(n31230), .B(n25602), .C(n31231), .D(n25613), .Y(n34719)
         );
  AOI22X1 U22082 ( .A(n25623), .B(reg_file[617]), .C(n25634), .D(reg_file[745]), .Y(n34717) );
  AOI22X1 U22083 ( .A(n25645), .B(reg_file[873]), .C(n25656), .D(
        reg_file[1001]), .Y(n34716) );
  NOR2X1 U22084 ( .A(n34721), .B(n34722), .Y(n34707) );
  NAND3X1 U22085 ( .A(n34723), .B(n34724), .C(n34725), .Y(n34722) );
  NOR2X1 U22086 ( .A(n34726), .B(n34727), .Y(n34725) );
  OAI22X1 U22087 ( .A(n31239), .B(n25667), .C(n31240), .D(n25678), .Y(n34727)
         );
  OAI22X1 U22088 ( .A(n31241), .B(n25688), .C(n31242), .D(n25699), .Y(n34726)
         );
  AOI22X1 U22089 ( .A(n25709), .B(reg_file[3561]), .C(n25720), .D(
        reg_file[3433]), .Y(n34724) );
  AOI22X1 U22090 ( .A(n25731), .B(reg_file[3305]), .C(n25742), .D(
        reg_file[3177]), .Y(n34723) );
  NAND3X1 U22091 ( .A(n34728), .B(n34729), .C(n34730), .Y(n34721) );
  NOR2X1 U22092 ( .A(n34731), .B(n34732), .Y(n34730) );
  OAI22X1 U22093 ( .A(n31248), .B(n25753), .C(n31249), .D(n25764), .Y(n34732)
         );
  OAI22X1 U22094 ( .A(n31250), .B(n25774), .C(n31251), .D(n25785), .Y(n34731)
         );
  AOI22X1 U22095 ( .A(n25795), .B(reg_file[2537]), .C(n25806), .D(
        reg_file[2409]), .Y(n34729) );
  AOI22X1 U22096 ( .A(n25817), .B(reg_file[2281]), .C(n25828), .D(
        reg_file[2153]), .Y(n34728) );
  AOI21X1 U22097 ( .A(n34733), .B(n34734), .C(n25484), .Y(rd1data1033_104_) );
  NOR2X1 U22098 ( .A(n34735), .B(n34736), .Y(n34734) );
  NAND3X1 U22099 ( .A(n34737), .B(n34738), .C(n34739), .Y(n34736) );
  NOR2X1 U22100 ( .A(n34740), .B(n34741), .Y(n34739) );
  OAI22X1 U22101 ( .A(n31261), .B(n25495), .C(n31262), .D(n25506), .Y(n34741)
         );
  OAI22X1 U22102 ( .A(n31263), .B(n25516), .C(n31264), .D(n25527), .Y(n34740)
         );
  AOI22X1 U22103 ( .A(n25537), .B(reg_file[1512]), .C(n25548), .D(
        reg_file[1384]), .Y(n34738) );
  AOI22X1 U22104 ( .A(n25559), .B(reg_file[1256]), .C(n25570), .D(
        reg_file[1128]), .Y(n34737) );
  NAND3X1 U22105 ( .A(n34742), .B(n34743), .C(n34744), .Y(n34735) );
  NOR2X1 U22106 ( .A(n34745), .B(n34746), .Y(n34744) );
  OAI22X1 U22107 ( .A(n31270), .B(n25581), .C(n31271), .D(n25592), .Y(n34746)
         );
  OAI22X1 U22108 ( .A(n31272), .B(n25602), .C(n31273), .D(n25613), .Y(n34745)
         );
  AOI22X1 U22109 ( .A(n25623), .B(reg_file[616]), .C(n25634), .D(reg_file[744]), .Y(n34743) );
  AOI22X1 U22110 ( .A(n25645), .B(reg_file[872]), .C(n25656), .D(
        reg_file[1000]), .Y(n34742) );
  NOR2X1 U22111 ( .A(n34747), .B(n34748), .Y(n34733) );
  NAND3X1 U22112 ( .A(n34749), .B(n34750), .C(n34751), .Y(n34748) );
  NOR2X1 U22113 ( .A(n34752), .B(n34753), .Y(n34751) );
  OAI22X1 U22114 ( .A(n31281), .B(n25667), .C(n31282), .D(n25678), .Y(n34753)
         );
  OAI22X1 U22115 ( .A(n31283), .B(n25688), .C(n31284), .D(n25699), .Y(n34752)
         );
  AOI22X1 U22116 ( .A(n25709), .B(reg_file[3560]), .C(n25720), .D(
        reg_file[3432]), .Y(n34750) );
  AOI22X1 U22117 ( .A(n25731), .B(reg_file[3304]), .C(n25742), .D(
        reg_file[3176]), .Y(n34749) );
  NAND3X1 U22118 ( .A(n34754), .B(n34755), .C(n34756), .Y(n34747) );
  NOR2X1 U22119 ( .A(n34757), .B(n34758), .Y(n34756) );
  OAI22X1 U22120 ( .A(n31290), .B(n25753), .C(n31291), .D(n25764), .Y(n34758)
         );
  OAI22X1 U22121 ( .A(n31292), .B(n25774), .C(n31293), .D(n25785), .Y(n34757)
         );
  AOI22X1 U22122 ( .A(n25795), .B(reg_file[2536]), .C(n25806), .D(
        reg_file[2408]), .Y(n34755) );
  AOI22X1 U22123 ( .A(n25817), .B(reg_file[2280]), .C(n25828), .D(
        reg_file[2152]), .Y(n34754) );
  AOI21X1 U22124 ( .A(n34759), .B(n34760), .C(n25484), .Y(rd1data1033_103_) );
  NOR2X1 U22125 ( .A(n34761), .B(n34762), .Y(n34760) );
  NAND3X1 U22126 ( .A(n34763), .B(n34764), .C(n34765), .Y(n34762) );
  NOR2X1 U22127 ( .A(n34766), .B(n34767), .Y(n34765) );
  OAI22X1 U22128 ( .A(n31303), .B(n25495), .C(n31304), .D(n25506), .Y(n34767)
         );
  OAI22X1 U22129 ( .A(n31305), .B(n25516), .C(n31306), .D(n25527), .Y(n34766)
         );
  AOI22X1 U22130 ( .A(n25537), .B(reg_file[1511]), .C(n25548), .D(
        reg_file[1383]), .Y(n34764) );
  AOI22X1 U22131 ( .A(n25559), .B(reg_file[1255]), .C(n25570), .D(
        reg_file[1127]), .Y(n34763) );
  NAND3X1 U22132 ( .A(n34768), .B(n34769), .C(n34770), .Y(n34761) );
  NOR2X1 U22133 ( .A(n34771), .B(n34772), .Y(n34770) );
  OAI22X1 U22134 ( .A(n31312), .B(n25581), .C(n31313), .D(n25592), .Y(n34772)
         );
  OAI22X1 U22135 ( .A(n31314), .B(n25602), .C(n31315), .D(n25613), .Y(n34771)
         );
  AOI22X1 U22136 ( .A(n25623), .B(reg_file[615]), .C(n25634), .D(reg_file[743]), .Y(n34769) );
  AOI22X1 U22137 ( .A(n25645), .B(reg_file[871]), .C(n25656), .D(reg_file[999]), .Y(n34768) );
  NOR2X1 U22138 ( .A(n34773), .B(n34774), .Y(n34759) );
  NAND3X1 U22139 ( .A(n34775), .B(n34776), .C(n34777), .Y(n34774) );
  NOR2X1 U22140 ( .A(n34778), .B(n34779), .Y(n34777) );
  OAI22X1 U22141 ( .A(n31323), .B(n25667), .C(n31324), .D(n25678), .Y(n34779)
         );
  OAI22X1 U22142 ( .A(n31325), .B(n25688), .C(n31326), .D(n25699), .Y(n34778)
         );
  AOI22X1 U22143 ( .A(n25709), .B(reg_file[3559]), .C(n25720), .D(
        reg_file[3431]), .Y(n34776) );
  AOI22X1 U22144 ( .A(n25731), .B(reg_file[3303]), .C(n25742), .D(
        reg_file[3175]), .Y(n34775) );
  NAND3X1 U22145 ( .A(n34780), .B(n34781), .C(n34782), .Y(n34773) );
  NOR2X1 U22146 ( .A(n34783), .B(n34784), .Y(n34782) );
  OAI22X1 U22147 ( .A(n31332), .B(n25753), .C(n31333), .D(n25764), .Y(n34784)
         );
  OAI22X1 U22148 ( .A(n31334), .B(n25774), .C(n31335), .D(n25785), .Y(n34783)
         );
  AOI22X1 U22149 ( .A(n25795), .B(reg_file[2535]), .C(n25806), .D(
        reg_file[2407]), .Y(n34781) );
  AOI22X1 U22150 ( .A(n25817), .B(reg_file[2279]), .C(n25828), .D(
        reg_file[2151]), .Y(n34780) );
  AOI21X1 U22151 ( .A(n34785), .B(n34786), .C(n25484), .Y(rd1data1033_102_) );
  NOR2X1 U22152 ( .A(n34787), .B(n34788), .Y(n34786) );
  NAND3X1 U22153 ( .A(n34789), .B(n34790), .C(n34791), .Y(n34788) );
  NOR2X1 U22154 ( .A(n34792), .B(n34793), .Y(n34791) );
  OAI22X1 U22155 ( .A(n31345), .B(n25495), .C(n31346), .D(n25506), .Y(n34793)
         );
  OAI22X1 U22156 ( .A(n31347), .B(n25516), .C(n31348), .D(n25527), .Y(n34792)
         );
  AOI22X1 U22157 ( .A(n25537), .B(reg_file[1510]), .C(n25548), .D(
        reg_file[1382]), .Y(n34790) );
  AOI22X1 U22158 ( .A(n25559), .B(reg_file[1254]), .C(n25570), .D(
        reg_file[1126]), .Y(n34789) );
  NAND3X1 U22159 ( .A(n34794), .B(n34795), .C(n34796), .Y(n34787) );
  NOR2X1 U22160 ( .A(n34797), .B(n34798), .Y(n34796) );
  OAI22X1 U22161 ( .A(n31354), .B(n25581), .C(n31355), .D(n25592), .Y(n34798)
         );
  OAI22X1 U22162 ( .A(n31356), .B(n25602), .C(n31357), .D(n25613), .Y(n34797)
         );
  AOI22X1 U22163 ( .A(n25623), .B(reg_file[614]), .C(n25634), .D(reg_file[742]), .Y(n34795) );
  AOI22X1 U22164 ( .A(n25645), .B(reg_file[870]), .C(n25656), .D(reg_file[998]), .Y(n34794) );
  NOR2X1 U22165 ( .A(n34799), .B(n34800), .Y(n34785) );
  NAND3X1 U22166 ( .A(n34801), .B(n34802), .C(n34803), .Y(n34800) );
  NOR2X1 U22167 ( .A(n34804), .B(n34805), .Y(n34803) );
  OAI22X1 U22168 ( .A(n31365), .B(n25667), .C(n31366), .D(n25678), .Y(n34805)
         );
  OAI22X1 U22169 ( .A(n31367), .B(n25688), .C(n31368), .D(n25699), .Y(n34804)
         );
  AOI22X1 U22170 ( .A(n25709), .B(reg_file[3558]), .C(n25720), .D(
        reg_file[3430]), .Y(n34802) );
  AOI22X1 U22171 ( .A(n25731), .B(reg_file[3302]), .C(n25742), .D(
        reg_file[3174]), .Y(n34801) );
  NAND3X1 U22172 ( .A(n34806), .B(n34807), .C(n34808), .Y(n34799) );
  NOR2X1 U22173 ( .A(n34809), .B(n34810), .Y(n34808) );
  OAI22X1 U22174 ( .A(n31374), .B(n25753), .C(n31375), .D(n25764), .Y(n34810)
         );
  OAI22X1 U22175 ( .A(n31376), .B(n25774), .C(n31377), .D(n25785), .Y(n34809)
         );
  AOI22X1 U22176 ( .A(n25795), .B(reg_file[2534]), .C(n25806), .D(
        reg_file[2406]), .Y(n34807) );
  AOI22X1 U22177 ( .A(n25817), .B(reg_file[2278]), .C(n25828), .D(
        reg_file[2150]), .Y(n34806) );
  AOI21X1 U22178 ( .A(n34811), .B(n34812), .C(n25484), .Y(rd1data1033_101_) );
  NOR2X1 U22179 ( .A(n34813), .B(n34814), .Y(n34812) );
  NAND3X1 U22180 ( .A(n34815), .B(n34816), .C(n34817), .Y(n34814) );
  NOR2X1 U22181 ( .A(n34818), .B(n34819), .Y(n34817) );
  OAI22X1 U22182 ( .A(n31387), .B(n25495), .C(n31388), .D(n25506), .Y(n34819)
         );
  OAI22X1 U22183 ( .A(n31389), .B(n25516), .C(n31390), .D(n25527), .Y(n34818)
         );
  AOI22X1 U22184 ( .A(n25537), .B(reg_file[1509]), .C(n25548), .D(
        reg_file[1381]), .Y(n34816) );
  AOI22X1 U22185 ( .A(n25559), .B(reg_file[1253]), .C(n25570), .D(
        reg_file[1125]), .Y(n34815) );
  NAND3X1 U22186 ( .A(n34820), .B(n34821), .C(n34822), .Y(n34813) );
  NOR2X1 U22187 ( .A(n34823), .B(n34824), .Y(n34822) );
  OAI22X1 U22188 ( .A(n31396), .B(n25581), .C(n31397), .D(n25592), .Y(n34824)
         );
  OAI22X1 U22189 ( .A(n31398), .B(n25602), .C(n31399), .D(n25613), .Y(n34823)
         );
  AOI22X1 U22190 ( .A(n25623), .B(reg_file[613]), .C(n25634), .D(reg_file[741]), .Y(n34821) );
  AOI22X1 U22191 ( .A(n25645), .B(reg_file[869]), .C(n25656), .D(reg_file[997]), .Y(n34820) );
  NOR2X1 U22192 ( .A(n34825), .B(n34826), .Y(n34811) );
  NAND3X1 U22193 ( .A(n34827), .B(n34828), .C(n34829), .Y(n34826) );
  NOR2X1 U22194 ( .A(n34830), .B(n34831), .Y(n34829) );
  OAI22X1 U22195 ( .A(n31407), .B(n25667), .C(n31408), .D(n25678), .Y(n34831)
         );
  OAI22X1 U22196 ( .A(n31409), .B(n25688), .C(n31410), .D(n25699), .Y(n34830)
         );
  AOI22X1 U22197 ( .A(n25709), .B(reg_file[3557]), .C(n25720), .D(
        reg_file[3429]), .Y(n34828) );
  AOI22X1 U22198 ( .A(n25731), .B(reg_file[3301]), .C(n25742), .D(
        reg_file[3173]), .Y(n34827) );
  NAND3X1 U22199 ( .A(n34832), .B(n34833), .C(n34834), .Y(n34825) );
  NOR2X1 U22200 ( .A(n34835), .B(n34836), .Y(n34834) );
  OAI22X1 U22201 ( .A(n31416), .B(n25753), .C(n31417), .D(n25764), .Y(n34836)
         );
  OAI22X1 U22202 ( .A(n31418), .B(n25774), .C(n31419), .D(n25785), .Y(n34835)
         );
  AOI22X1 U22203 ( .A(n25795), .B(reg_file[2533]), .C(n25806), .D(
        reg_file[2405]), .Y(n34833) );
  AOI22X1 U22204 ( .A(n25817), .B(reg_file[2277]), .C(n25828), .D(
        reg_file[2149]), .Y(n34832) );
  AOI21X1 U22205 ( .A(n34837), .B(n34838), .C(n25484), .Y(rd1data1033_100_) );
  NOR2X1 U22206 ( .A(n34839), .B(n34840), .Y(n34838) );
  NAND3X1 U22207 ( .A(n34841), .B(n34842), .C(n34843), .Y(n34840) );
  NOR2X1 U22208 ( .A(n34844), .B(n34845), .Y(n34843) );
  OAI22X1 U22209 ( .A(n31429), .B(n25495), .C(n31430), .D(n25506), .Y(n34845)
         );
  OAI22X1 U22210 ( .A(n31431), .B(n25516), .C(n31432), .D(n25527), .Y(n34844)
         );
  AOI22X1 U22211 ( .A(n25537), .B(reg_file[1508]), .C(n25548), .D(
        reg_file[1380]), .Y(n34842) );
  AOI22X1 U22212 ( .A(n25559), .B(reg_file[1252]), .C(n25570), .D(
        reg_file[1124]), .Y(n34841) );
  NAND3X1 U22213 ( .A(n34846), .B(n34847), .C(n34848), .Y(n34839) );
  NOR2X1 U22214 ( .A(n34849), .B(n34850), .Y(n34848) );
  OAI22X1 U22215 ( .A(n31438), .B(n25581), .C(n31439), .D(n25592), .Y(n34850)
         );
  OAI22X1 U22216 ( .A(n31440), .B(n25602), .C(n31441), .D(n25613), .Y(n34849)
         );
  AOI22X1 U22217 ( .A(n25623), .B(reg_file[612]), .C(n25634), .D(reg_file[740]), .Y(n34847) );
  AOI22X1 U22218 ( .A(n25645), .B(reg_file[868]), .C(n25656), .D(reg_file[996]), .Y(n34846) );
  NOR2X1 U22219 ( .A(n34851), .B(n34852), .Y(n34837) );
  NAND3X1 U22220 ( .A(n34853), .B(n34854), .C(n34855), .Y(n34852) );
  NOR2X1 U22221 ( .A(n34856), .B(n34857), .Y(n34855) );
  OAI22X1 U22222 ( .A(n31449), .B(n25667), .C(n31450), .D(n25678), .Y(n34857)
         );
  OAI22X1 U22223 ( .A(n31451), .B(n25688), .C(n31452), .D(n25699), .Y(n34856)
         );
  AOI22X1 U22224 ( .A(n25709), .B(reg_file[3556]), .C(n25720), .D(
        reg_file[3428]), .Y(n34854) );
  AOI22X1 U22225 ( .A(n25731), .B(reg_file[3300]), .C(n25742), .D(
        reg_file[3172]), .Y(n34853) );
  NAND3X1 U22226 ( .A(n34858), .B(n34859), .C(n34860), .Y(n34851) );
  NOR2X1 U22227 ( .A(n34861), .B(n34862), .Y(n34860) );
  OAI22X1 U22228 ( .A(n31458), .B(n25753), .C(n31459), .D(n25764), .Y(n34862)
         );
  OAI22X1 U22229 ( .A(n31460), .B(n25774), .C(n31461), .D(n25785), .Y(n34861)
         );
  AOI22X1 U22230 ( .A(n25795), .B(reg_file[2532]), .C(n25806), .D(
        reg_file[2404]), .Y(n34859) );
  AOI22X1 U22231 ( .A(n25817), .B(reg_file[2276]), .C(n25828), .D(
        reg_file[2148]), .Y(n34858) );
  AOI21X1 U22232 ( .A(n34863), .B(n34864), .C(n25484), .Y(rd1data1033_0_) );
  INVX1 U22233 ( .A(rd1en), .Y(n31530) );
  NOR2X1 U22234 ( .A(n34865), .B(n34866), .Y(n34864) );
  NAND3X1 U22235 ( .A(n34867), .B(n34868), .C(n34869), .Y(n34866) );
  NOR2X1 U22236 ( .A(n34870), .B(n34871), .Y(n34869) );
  OAI22X1 U22237 ( .A(n31471), .B(n25495), .C(n31472), .D(n25506), .Y(n34871)
         );
  NAND2X1 U22238 ( .A(n34872), .B(n34873), .Y(n31539) );
  NAND2X1 U22239 ( .A(n34874), .B(n34873), .Y(n31538) );
  OAI22X1 U22240 ( .A(n31476), .B(n25516), .C(n31477), .D(n25527), .Y(n34870)
         );
  NAND2X1 U22241 ( .A(n34872), .B(n34875), .Y(n31541) );
  NAND2X1 U22242 ( .A(n34874), .B(n34875), .Y(n31540) );
  AOI22X1 U22243 ( .A(n25537), .B(reg_file[1408]), .C(n25548), .D(
        reg_file[1280]), .Y(n34868) );
  AND2X1 U22244 ( .A(n34874), .B(n34876), .Y(n31543) );
  AND2X1 U22245 ( .A(n34872), .B(n34876), .Y(n31542) );
  AOI22X1 U22246 ( .A(n25559), .B(reg_file[1152]), .C(n25570), .D(
        reg_file[1024]), .Y(n34867) );
  AND2X1 U22247 ( .A(n34874), .B(n34877), .Y(n31545) );
  INVX1 U22248 ( .A(n34878), .Y(n34874) );
  NAND3X1 U22249 ( .A(n34879), .B(n34880), .C(rd1addr[3]), .Y(n34878) );
  AND2X1 U22250 ( .A(n34872), .B(n34877), .Y(n31544) );
  INVX1 U22251 ( .A(n34881), .Y(n34872) );
  NAND3X1 U22252 ( .A(rd1addr[0]), .B(n34880), .C(rd1addr[3]), .Y(n34881) );
  NAND3X1 U22253 ( .A(n34882), .B(n34883), .C(n34884), .Y(n34865) );
  NOR2X1 U22254 ( .A(n34885), .B(n34886), .Y(n34884) );
  OAI22X1 U22255 ( .A(n31490), .B(n25581), .C(n31491), .D(n25592), .Y(n34886)
         );
  NAND2X1 U22256 ( .A(n34876), .B(n34887), .Y(n31552) );
  NAND2X1 U22257 ( .A(n34876), .B(n34888), .Y(n31551) );
  OAI22X1 U22258 ( .A(n31494), .B(n25602), .C(n31495), .D(n25613), .Y(n34885)
         );
  NAND2X1 U22259 ( .A(n34877), .B(n34887), .Y(n31554) );
  NAND2X1 U22260 ( .A(n34888), .B(n34877), .Y(n31553) );
  AOI22X1 U22261 ( .A(n25623), .B(reg_file[512]), .C(n25634), .D(reg_file[640]), .Y(n34883) );
  AND2X1 U22262 ( .A(n34873), .B(n34888), .Y(n31556) );
  AND2X1 U22263 ( .A(n34873), .B(n34887), .Y(n31555) );
  AOI22X1 U22264 ( .A(n25645), .B(reg_file[768]), .C(n25656), .D(reg_file[896]), .Y(n34882) );
  AND2X1 U22265 ( .A(n34875), .B(n34888), .Y(n31558) );
  INVX1 U22266 ( .A(n34889), .Y(n34888) );
  NAND3X1 U22267 ( .A(n34890), .B(n34880), .C(rd1addr[0]), .Y(n34889) );
  AND2X1 U22268 ( .A(n34875), .B(n34887), .Y(n31557) );
  INVX1 U22269 ( .A(n34891), .Y(n34887) );
  NAND3X1 U22270 ( .A(n34890), .B(n34880), .C(n34879), .Y(n34891) );
  INVX1 U22271 ( .A(rd1addr[4]), .Y(n34880) );
  NOR2X1 U22272 ( .A(n34892), .B(n34893), .Y(n34863) );
  NAND3X1 U22273 ( .A(n34894), .B(n34895), .C(n34896), .Y(n34893) );
  NOR2X1 U22274 ( .A(n34897), .B(n34898), .Y(n34896) );
  OAI22X1 U22275 ( .A(n31506), .B(n25667), .C(n31507), .D(n25678), .Y(n34898)
         );
  NAND2X1 U22276 ( .A(n34899), .B(n34873), .Y(n31567) );
  NAND2X1 U22277 ( .A(n34900), .B(n34873), .Y(n31566) );
  OAI22X1 U22278 ( .A(n31510), .B(n25688), .C(n31511), .D(n25699), .Y(n34897)
         );
  NAND2X1 U22279 ( .A(n34899), .B(n34875), .Y(n31569) );
  NAND2X1 U22280 ( .A(n34900), .B(n34875), .Y(n31568) );
  AOI22X1 U22281 ( .A(n25709), .B(reg_file[3456]), .C(n25720), .D(
        reg_file[3328]), .Y(n34895) );
  AND2X1 U22282 ( .A(n34900), .B(n34876), .Y(n31571) );
  AND2X1 U22283 ( .A(n34899), .B(n34876), .Y(n31570) );
  AOI22X1 U22284 ( .A(n25731), .B(reg_file[3200]), .C(n25742), .D(
        reg_file[3072]), .Y(n34894) );
  AND2X1 U22285 ( .A(n34900), .B(n34877), .Y(n31573) );
  INVX1 U22286 ( .A(n34901), .Y(n34900) );
  NAND3X1 U22287 ( .A(rd1addr[3]), .B(n34879), .C(rd1addr[4]), .Y(n34901) );
  AND2X1 U22288 ( .A(n34899), .B(n34877), .Y(n31572) );
  INVX1 U22289 ( .A(n34902), .Y(n34899) );
  NAND3X1 U22290 ( .A(rd1addr[3]), .B(rd1addr[0]), .C(rd1addr[4]), .Y(n34902)
         );
  NAND3X1 U22291 ( .A(n34903), .B(n34904), .C(n34905), .Y(n34892) );
  NOR2X1 U22292 ( .A(n34906), .B(n34907), .Y(n34905) );
  OAI22X1 U22293 ( .A(n31519), .B(n25753), .C(n31520), .D(n25764), .Y(n34907)
         );
  NAND2X1 U22294 ( .A(n34908), .B(n34873), .Y(n31580) );
  NAND2X1 U22295 ( .A(n34909), .B(n34873), .Y(n31579) );
  AND2X1 U22296 ( .A(rd1addr[2]), .B(n34910), .Y(n34873) );
  OAI22X1 U22297 ( .A(n31524), .B(n25774), .C(n31525), .D(n25785), .Y(n34906)
         );
  NAND2X1 U22298 ( .A(n34908), .B(n34875), .Y(n31582) );
  NAND2X1 U22299 ( .A(n34909), .B(n34875), .Y(n31581) );
  AND2X1 U22300 ( .A(rd1addr[2]), .B(rd1addr[1]), .Y(n34875) );
  AOI22X1 U22301 ( .A(n25795), .B(reg_file[2432]), .C(n25806), .D(
        reg_file[2304]), .Y(n34904) );
  AND2X1 U22302 ( .A(n34909), .B(n34876), .Y(n31584) );
  AND2X1 U22303 ( .A(n34908), .B(n34876), .Y(n31583) );
  NOR2X1 U22304 ( .A(n34910), .B(rd1addr[2]), .Y(n34876) );
  INVX1 U22305 ( .A(rd1addr[1]), .Y(n34910) );
  AOI22X1 U22306 ( .A(n25817), .B(reg_file[2176]), .C(n25828), .D(
        reg_file[2048]), .Y(n34903) );
  AND2X1 U22307 ( .A(n34909), .B(n34877), .Y(n31586) );
  INVX1 U22308 ( .A(n34911), .Y(n34909) );
  NAND3X1 U22309 ( .A(n34879), .B(n34890), .C(rd1addr[4]), .Y(n34911) );
  INVX1 U22310 ( .A(rd1addr[0]), .Y(n34879) );
  AND2X1 U22311 ( .A(n34908), .B(n34877), .Y(n31585) );
  NOR2X1 U22312 ( .A(rd1addr[1]), .B(rd1addr[2]), .Y(n34877) );
  INVX1 U22313 ( .A(n34912), .Y(n34908) );
  NAND3X1 U22314 ( .A(rd1addr[0]), .B(n34890), .C(rd1addr[4]), .Y(n34912) );
  INVX1 U22315 ( .A(rd1addr[3]), .Y(n34890) );
  MUX2X1 U22316 ( .B(n31495), .A(n25129), .S(n25839), .Y(n25128) );
  INVX1 U22317 ( .A(reg_file[0]), .Y(n31495) );
  MUX2X1 U22318 ( .B(n29845), .A(n25130), .S(n25839), .Y(n25127) );
  INVX1 U22319 ( .A(reg_file[1]), .Y(n29845) );
  MUX2X1 U22320 ( .B(n29383), .A(n25131), .S(n25839), .Y(n25126) );
  INVX1 U22321 ( .A(reg_file[2]), .Y(n29383) );
  MUX2X1 U22322 ( .B(n28921), .A(n25132), .S(n25839), .Y(n25125) );
  INVX1 U22323 ( .A(reg_file[3]), .Y(n28921) );
  MUX2X1 U22324 ( .B(n28459), .A(n25133), .S(n25839), .Y(n25124) );
  INVX1 U22325 ( .A(reg_file[4]), .Y(n28459) );
  MUX2X1 U22326 ( .B(n27997), .A(n25134), .S(n25839), .Y(n25123) );
  INVX1 U22327 ( .A(reg_file[5]), .Y(n27997) );
  MUX2X1 U22328 ( .B(n27535), .A(n25135), .S(n25839), .Y(n25122) );
  INVX1 U22329 ( .A(reg_file[6]), .Y(n27535) );
  MUX2X1 U22330 ( .B(n27073), .A(n25136), .S(n25839), .Y(n25121) );
  INVX1 U22331 ( .A(reg_file[7]), .Y(n27073) );
  NOR2X1 U22332 ( .A(n25839), .B(n26611), .Y(n25120) );
  INVX1 U22333 ( .A(reg_file[8]), .Y(n26611) );
  NOR2X1 U22334 ( .A(n25839), .B(n26129), .Y(n25119) );
  INVX1 U22335 ( .A(reg_file[9]), .Y(n26129) );
  NOR2X1 U22336 ( .A(n25839), .B(n31021), .Y(n25118) );
  INVX1 U22337 ( .A(reg_file[10]), .Y(n31021) );
  NOR2X1 U22338 ( .A(n25839), .B(n30559), .Y(n25117) );
  INVX1 U22339 ( .A(reg_file[11]), .Y(n30559) );
  NOR2X1 U22340 ( .A(n25839), .B(n30181), .Y(n25116) );
  INVX1 U22341 ( .A(reg_file[12]), .Y(n30181) );
  NOR2X1 U22342 ( .A(n25839), .B(n30139), .Y(n25115) );
  INVX1 U22343 ( .A(reg_file[13]), .Y(n30139) );
  NOR2X1 U22344 ( .A(n25840), .B(n30097), .Y(n25114) );
  INVX1 U22345 ( .A(reg_file[14]), .Y(n30097) );
  NOR2X1 U22346 ( .A(n25840), .B(n30055), .Y(n25113) );
  INVX1 U22347 ( .A(reg_file[15]), .Y(n30055) );
  NOR2X1 U22348 ( .A(n25840), .B(n30013), .Y(n25112) );
  INVX1 U22349 ( .A(reg_file[16]), .Y(n30013) );
  NOR2X1 U22350 ( .A(n25840), .B(n29971), .Y(n25111) );
  INVX1 U22351 ( .A(reg_file[17]), .Y(n29971) );
  NOR2X1 U22352 ( .A(n25840), .B(n29929), .Y(n25110) );
  INVX1 U22353 ( .A(reg_file[18]), .Y(n29929) );
  NOR2X1 U22354 ( .A(n25840), .B(n29887), .Y(n25109) );
  INVX1 U22355 ( .A(reg_file[19]), .Y(n29887) );
  NOR2X1 U22356 ( .A(n25840), .B(n29803), .Y(n25108) );
  INVX1 U22357 ( .A(reg_file[20]), .Y(n29803) );
  NOR2X1 U22358 ( .A(n25840), .B(n29761), .Y(n25107) );
  INVX1 U22359 ( .A(reg_file[21]), .Y(n29761) );
  NOR2X1 U22360 ( .A(n25840), .B(n29719), .Y(n25106) );
  INVX1 U22361 ( .A(reg_file[22]), .Y(n29719) );
  NOR2X1 U22362 ( .A(n25840), .B(n29677), .Y(n25105) );
  INVX1 U22363 ( .A(reg_file[23]), .Y(n29677) );
  NOR2X1 U22364 ( .A(n25840), .B(n29635), .Y(n25104) );
  INVX1 U22365 ( .A(reg_file[24]), .Y(n29635) );
  NOR2X1 U22366 ( .A(n25840), .B(n29593), .Y(n25103) );
  INVX1 U22367 ( .A(reg_file[25]), .Y(n29593) );
  NOR2X1 U22368 ( .A(n25840), .B(n29551), .Y(n25102) );
  INVX1 U22369 ( .A(reg_file[26]), .Y(n29551) );
  NOR2X1 U22370 ( .A(n25840), .B(n29509), .Y(n25101) );
  INVX1 U22371 ( .A(reg_file[27]), .Y(n29509) );
  NOR2X1 U22372 ( .A(n25840), .B(n29467), .Y(n25100) );
  INVX1 U22373 ( .A(reg_file[28]), .Y(n29467) );
  NOR2X1 U22374 ( .A(n25840), .B(n29425), .Y(n25099) );
  INVX1 U22375 ( .A(reg_file[29]), .Y(n29425) );
  NOR2X1 U22376 ( .A(n25840), .B(n29341), .Y(n25098) );
  INVX1 U22377 ( .A(reg_file[30]), .Y(n29341) );
  NOR2X1 U22378 ( .A(n25841), .B(n29299), .Y(n25097) );
  INVX1 U22379 ( .A(reg_file[31]), .Y(n29299) );
  NOR2X1 U22380 ( .A(n25841), .B(n29257), .Y(n25096) );
  INVX1 U22381 ( .A(reg_file[32]), .Y(n29257) );
  NOR2X1 U22382 ( .A(n25841), .B(n29215), .Y(n25095) );
  INVX1 U22383 ( .A(reg_file[33]), .Y(n29215) );
  NOR2X1 U22384 ( .A(n25841), .B(n29173), .Y(n25094) );
  INVX1 U22385 ( .A(reg_file[34]), .Y(n29173) );
  NOR2X1 U22386 ( .A(n25841), .B(n29131), .Y(n25093) );
  INVX1 U22387 ( .A(reg_file[35]), .Y(n29131) );
  NOR2X1 U22388 ( .A(n25841), .B(n29089), .Y(n25092) );
  INVX1 U22389 ( .A(reg_file[36]), .Y(n29089) );
  NOR2X1 U22390 ( .A(n25841), .B(n29047), .Y(n25091) );
  INVX1 U22391 ( .A(reg_file[37]), .Y(n29047) );
  NOR2X1 U22392 ( .A(n25841), .B(n29005), .Y(n25090) );
  INVX1 U22393 ( .A(reg_file[38]), .Y(n29005) );
  NOR2X1 U22394 ( .A(n25841), .B(n28963), .Y(n25089) );
  INVX1 U22395 ( .A(reg_file[39]), .Y(n28963) );
  NOR2X1 U22396 ( .A(n25841), .B(n28879), .Y(n25088) );
  INVX1 U22397 ( .A(reg_file[40]), .Y(n28879) );
  NOR2X1 U22398 ( .A(n25841), .B(n28837), .Y(n25087) );
  INVX1 U22399 ( .A(reg_file[41]), .Y(n28837) );
  NOR2X1 U22400 ( .A(n25841), .B(n28795), .Y(n25086) );
  INVX1 U22401 ( .A(reg_file[42]), .Y(n28795) );
  NOR2X1 U22402 ( .A(n25841), .B(n28753), .Y(n25085) );
  INVX1 U22403 ( .A(reg_file[43]), .Y(n28753) );
  NOR2X1 U22404 ( .A(n25841), .B(n28711), .Y(n25084) );
  INVX1 U22405 ( .A(reg_file[44]), .Y(n28711) );
  NOR2X1 U22406 ( .A(n25841), .B(n28669), .Y(n25083) );
  INVX1 U22407 ( .A(reg_file[45]), .Y(n28669) );
  NOR2X1 U22408 ( .A(n25841), .B(n28627), .Y(n25082) );
  INVX1 U22409 ( .A(reg_file[46]), .Y(n28627) );
  NOR2X1 U22410 ( .A(n25841), .B(n28585), .Y(n25081) );
  INVX1 U22411 ( .A(reg_file[47]), .Y(n28585) );
  NOR2X1 U22412 ( .A(n25842), .B(n28543), .Y(n25080) );
  INVX1 U22413 ( .A(reg_file[48]), .Y(n28543) );
  NOR2X1 U22414 ( .A(n25842), .B(n28501), .Y(n25079) );
  INVX1 U22415 ( .A(reg_file[49]), .Y(n28501) );
  NOR2X1 U22416 ( .A(n25842), .B(n28417), .Y(n25078) );
  INVX1 U22417 ( .A(reg_file[50]), .Y(n28417) );
  NOR2X1 U22418 ( .A(n25842), .B(n28375), .Y(n25077) );
  INVX1 U22419 ( .A(reg_file[51]), .Y(n28375) );
  NOR2X1 U22420 ( .A(n25842), .B(n28333), .Y(n25076) );
  INVX1 U22421 ( .A(reg_file[52]), .Y(n28333) );
  NOR2X1 U22422 ( .A(n25842), .B(n28291), .Y(n25075) );
  INVX1 U22423 ( .A(reg_file[53]), .Y(n28291) );
  NOR2X1 U22424 ( .A(n25842), .B(n28249), .Y(n25074) );
  INVX1 U22425 ( .A(reg_file[54]), .Y(n28249) );
  NOR2X1 U22426 ( .A(n25842), .B(n28207), .Y(n25073) );
  INVX1 U22427 ( .A(reg_file[55]), .Y(n28207) );
  NOR2X1 U22428 ( .A(n25842), .B(n28165), .Y(n25072) );
  INVX1 U22429 ( .A(reg_file[56]), .Y(n28165) );
  NOR2X1 U22430 ( .A(n25842), .B(n28123), .Y(n25071) );
  INVX1 U22431 ( .A(reg_file[57]), .Y(n28123) );
  NOR2X1 U22432 ( .A(n25842), .B(n28081), .Y(n25070) );
  INVX1 U22433 ( .A(reg_file[58]), .Y(n28081) );
  NOR2X1 U22434 ( .A(n25842), .B(n28039), .Y(n25069) );
  INVX1 U22435 ( .A(reg_file[59]), .Y(n28039) );
  NOR2X1 U22436 ( .A(n25842), .B(n27955), .Y(n25068) );
  INVX1 U22437 ( .A(reg_file[60]), .Y(n27955) );
  NOR2X1 U22438 ( .A(n25842), .B(n27913), .Y(n25067) );
  INVX1 U22439 ( .A(reg_file[61]), .Y(n27913) );
  NOR2X1 U22440 ( .A(n25842), .B(n27871), .Y(n25066) );
  INVX1 U22441 ( .A(reg_file[62]), .Y(n27871) );
  NOR2X1 U22442 ( .A(n25842), .B(n27829), .Y(n25065) );
  INVX1 U22443 ( .A(reg_file[63]), .Y(n27829) );
  NOR2X1 U22444 ( .A(n25842), .B(n27787), .Y(n25064) );
  INVX1 U22445 ( .A(reg_file[64]), .Y(n27787) );
  NOR2X1 U22446 ( .A(n25843), .B(n27745), .Y(n25063) );
  INVX1 U22447 ( .A(reg_file[65]), .Y(n27745) );
  NOR2X1 U22448 ( .A(n25843), .B(n27703), .Y(n25062) );
  INVX1 U22449 ( .A(reg_file[66]), .Y(n27703) );
  NOR2X1 U22450 ( .A(n25843), .B(n27661), .Y(n25061) );
  INVX1 U22451 ( .A(reg_file[67]), .Y(n27661) );
  NOR2X1 U22452 ( .A(n25843), .B(n27619), .Y(n25060) );
  INVX1 U22453 ( .A(reg_file[68]), .Y(n27619) );
  NOR2X1 U22454 ( .A(n25843), .B(n27577), .Y(n25059) );
  INVX1 U22455 ( .A(reg_file[69]), .Y(n27577) );
  NOR2X1 U22456 ( .A(n25843), .B(n27493), .Y(n25058) );
  INVX1 U22457 ( .A(reg_file[70]), .Y(n27493) );
  NOR2X1 U22458 ( .A(n25843), .B(n27451), .Y(n25057) );
  INVX1 U22459 ( .A(reg_file[71]), .Y(n27451) );
  NOR2X1 U22460 ( .A(n25843), .B(n27409), .Y(n25056) );
  INVX1 U22461 ( .A(reg_file[72]), .Y(n27409) );
  NOR2X1 U22462 ( .A(n25843), .B(n27367), .Y(n25055) );
  INVX1 U22463 ( .A(reg_file[73]), .Y(n27367) );
  NOR2X1 U22464 ( .A(n25843), .B(n27325), .Y(n25054) );
  INVX1 U22465 ( .A(reg_file[74]), .Y(n27325) );
  NOR2X1 U22466 ( .A(n25843), .B(n27283), .Y(n25053) );
  INVX1 U22467 ( .A(reg_file[75]), .Y(n27283) );
  NOR2X1 U22468 ( .A(n25843), .B(n27241), .Y(n25052) );
  INVX1 U22469 ( .A(reg_file[76]), .Y(n27241) );
  NOR2X1 U22470 ( .A(n25843), .B(n27199), .Y(n25051) );
  INVX1 U22471 ( .A(reg_file[77]), .Y(n27199) );
  NOR2X1 U22472 ( .A(n25843), .B(n27157), .Y(n25050) );
  INVX1 U22473 ( .A(reg_file[78]), .Y(n27157) );
  NOR2X1 U22474 ( .A(n25843), .B(n27115), .Y(n25049) );
  INVX1 U22475 ( .A(reg_file[79]), .Y(n27115) );
  NOR2X1 U22476 ( .A(n25843), .B(n27031), .Y(n25048) );
  INVX1 U22477 ( .A(reg_file[80]), .Y(n27031) );
  NOR2X1 U22478 ( .A(n25843), .B(n26989), .Y(n25047) );
  INVX1 U22479 ( .A(reg_file[81]), .Y(n26989) );
  NOR2X1 U22480 ( .A(n25844), .B(n26947), .Y(n25046) );
  INVX1 U22481 ( .A(reg_file[82]), .Y(n26947) );
  NOR2X1 U22482 ( .A(n25844), .B(n26905), .Y(n25045) );
  INVX1 U22483 ( .A(reg_file[83]), .Y(n26905) );
  NOR2X1 U22484 ( .A(n25844), .B(n26863), .Y(n25044) );
  INVX1 U22485 ( .A(reg_file[84]), .Y(n26863) );
  NOR2X1 U22486 ( .A(n25844), .B(n26821), .Y(n25043) );
  INVX1 U22487 ( .A(reg_file[85]), .Y(n26821) );
  NOR2X1 U22488 ( .A(n25844), .B(n26779), .Y(n25042) );
  INVX1 U22489 ( .A(reg_file[86]), .Y(n26779) );
  NOR2X1 U22490 ( .A(n25844), .B(n26737), .Y(n25041) );
  INVX1 U22491 ( .A(reg_file[87]), .Y(n26737) );
  NOR2X1 U22492 ( .A(n25844), .B(n26695), .Y(n25040) );
  INVX1 U22493 ( .A(reg_file[88]), .Y(n26695) );
  NOR2X1 U22494 ( .A(n25844), .B(n26653), .Y(n25039) );
  INVX1 U22495 ( .A(reg_file[89]), .Y(n26653) );
  NOR2X1 U22496 ( .A(n25844), .B(n26569), .Y(n25038) );
  INVX1 U22497 ( .A(reg_file[90]), .Y(n26569) );
  NOR2X1 U22498 ( .A(n25844), .B(n26527), .Y(n25037) );
  INVX1 U22499 ( .A(reg_file[91]), .Y(n26527) );
  NOR2X1 U22500 ( .A(n25844), .B(n26485), .Y(n25036) );
  INVX1 U22501 ( .A(reg_file[92]), .Y(n26485) );
  NOR2X1 U22502 ( .A(n25844), .B(n26443), .Y(n25035) );
  INVX1 U22503 ( .A(reg_file[93]), .Y(n26443) );
  NOR2X1 U22504 ( .A(n25844), .B(n26401), .Y(n25034) );
  INVX1 U22505 ( .A(reg_file[94]), .Y(n26401) );
  NOR2X1 U22506 ( .A(n25844), .B(n26359), .Y(n25033) );
  INVX1 U22507 ( .A(reg_file[95]), .Y(n26359) );
  NOR2X1 U22508 ( .A(n25844), .B(n26317), .Y(n25032) );
  INVX1 U22509 ( .A(reg_file[96]), .Y(n26317) );
  NOR2X1 U22510 ( .A(n25844), .B(n26275), .Y(n25031) );
  INVX1 U22511 ( .A(reg_file[97]), .Y(n26275) );
  NOR2X1 U22512 ( .A(n25844), .B(n26233), .Y(n25030) );
  INVX1 U22513 ( .A(reg_file[98]), .Y(n26233) );
  NOR2X1 U22514 ( .A(n25845), .B(n26191), .Y(n25029) );
  INVX1 U22515 ( .A(reg_file[99]), .Y(n26191) );
  NOR2X1 U22516 ( .A(n25845), .B(n31441), .Y(n25028) );
  INVX1 U22517 ( .A(reg_file[100]), .Y(n31441) );
  NOR2X1 U22518 ( .A(n25845), .B(n31399), .Y(n25027) );
  INVX1 U22519 ( .A(reg_file[101]), .Y(n31399) );
  NOR2X1 U22520 ( .A(n25845), .B(n31357), .Y(n25026) );
  INVX1 U22521 ( .A(reg_file[102]), .Y(n31357) );
  NOR2X1 U22522 ( .A(n25845), .B(n31315), .Y(n25025) );
  INVX1 U22523 ( .A(reg_file[103]), .Y(n31315) );
  NOR2X1 U22524 ( .A(n25845), .B(n31273), .Y(n25024) );
  INVX1 U22525 ( .A(reg_file[104]), .Y(n31273) );
  NOR2X1 U22526 ( .A(n25845), .B(n31231), .Y(n25023) );
  INVX1 U22527 ( .A(reg_file[105]), .Y(n31231) );
  NOR2X1 U22528 ( .A(n25845), .B(n31189), .Y(n25022) );
  INVX1 U22529 ( .A(reg_file[106]), .Y(n31189) );
  NOR2X1 U22530 ( .A(n25845), .B(n31147), .Y(n25021) );
  INVX1 U22531 ( .A(reg_file[107]), .Y(n31147) );
  NOR2X1 U22532 ( .A(n25845), .B(n31105), .Y(n25020) );
  INVX1 U22533 ( .A(reg_file[108]), .Y(n31105) );
  NOR2X1 U22534 ( .A(n25845), .B(n31063), .Y(n25019) );
  INVX1 U22535 ( .A(reg_file[109]), .Y(n31063) );
  NOR2X1 U22536 ( .A(n25845), .B(n30979), .Y(n25018) );
  INVX1 U22537 ( .A(reg_file[110]), .Y(n30979) );
  NOR2X1 U22538 ( .A(n25845), .B(n30937), .Y(n25017) );
  INVX1 U22539 ( .A(reg_file[111]), .Y(n30937) );
  NOR2X1 U22540 ( .A(n25845), .B(n30895), .Y(n25016) );
  INVX1 U22541 ( .A(reg_file[112]), .Y(n30895) );
  NOR2X1 U22542 ( .A(n25845), .B(n30853), .Y(n25015) );
  INVX1 U22543 ( .A(reg_file[113]), .Y(n30853) );
  NOR2X1 U22544 ( .A(n25845), .B(n30811), .Y(n25014) );
  INVX1 U22545 ( .A(reg_file[114]), .Y(n30811) );
  NOR2X1 U22546 ( .A(n25845), .B(n30769), .Y(n25013) );
  INVX1 U22547 ( .A(reg_file[115]), .Y(n30769) );
  NOR2X1 U22548 ( .A(n25846), .B(n30727), .Y(n25012) );
  INVX1 U22549 ( .A(reg_file[116]), .Y(n30727) );
  NOR2X1 U22550 ( .A(n25846), .B(n30685), .Y(n25011) );
  INVX1 U22551 ( .A(reg_file[117]), .Y(n30685) );
  NOR2X1 U22552 ( .A(n25846), .B(n30643), .Y(n25010) );
  INVX1 U22553 ( .A(reg_file[118]), .Y(n30643) );
  NOR2X1 U22554 ( .A(n25846), .B(n30601), .Y(n25009) );
  INVX1 U22555 ( .A(reg_file[119]), .Y(n30601) );
  NOR2X1 U22556 ( .A(n25846), .B(n30517), .Y(n25008) );
  INVX1 U22557 ( .A(reg_file[120]), .Y(n30517) );
  NOR2X1 U22558 ( .A(n25846), .B(n30475), .Y(n25007) );
  INVX1 U22559 ( .A(reg_file[121]), .Y(n30475) );
  NOR2X1 U22560 ( .A(n25846), .B(n30433), .Y(n25006) );
  INVX1 U22561 ( .A(reg_file[122]), .Y(n30433) );
  NOR2X1 U22562 ( .A(n25846), .B(n30391), .Y(n25005) );
  INVX1 U22563 ( .A(reg_file[123]), .Y(n30391) );
  NOR2X1 U22564 ( .A(n25846), .B(n30349), .Y(n25004) );
  INVX1 U22565 ( .A(reg_file[124]), .Y(n30349) );
  NOR2X1 U22566 ( .A(n25846), .B(n30307), .Y(n25003) );
  INVX1 U22567 ( .A(reg_file[125]), .Y(n30307) );
  NOR2X1 U22568 ( .A(n25846), .B(n30265), .Y(n25002) );
  INVX1 U22569 ( .A(reg_file[126]), .Y(n30265) );
  NOR2X1 U22570 ( .A(n25846), .B(n30223), .Y(n25001) );
  INVX1 U22571 ( .A(reg_file[127]), .Y(n30223) );
  NOR2X1 U22572 ( .A(n34922), .B(n34923), .Y(n34914) );
  MUX2X1 U22573 ( .B(n31494), .A(n25129), .S(n25847), .Y(n25000) );
  INVX1 U22574 ( .A(reg_file[128]), .Y(n31494) );
  MUX2X1 U22575 ( .B(n29844), .A(n25130), .S(n25847), .Y(n24999) );
  INVX1 U22576 ( .A(reg_file[129]), .Y(n29844) );
  MUX2X1 U22577 ( .B(n29382), .A(n25131), .S(n25847), .Y(n24998) );
  INVX1 U22578 ( .A(reg_file[130]), .Y(n29382) );
  MUX2X1 U22579 ( .B(n28920), .A(n25132), .S(n25847), .Y(n24997) );
  INVX1 U22580 ( .A(reg_file[131]), .Y(n28920) );
  MUX2X1 U22581 ( .B(n28458), .A(n25133), .S(n25847), .Y(n24996) );
  INVX1 U22582 ( .A(reg_file[132]), .Y(n28458) );
  MUX2X1 U22583 ( .B(n27996), .A(n25134), .S(n25847), .Y(n24995) );
  INVX1 U22584 ( .A(reg_file[133]), .Y(n27996) );
  MUX2X1 U22585 ( .B(n27534), .A(n25135), .S(n25847), .Y(n24994) );
  INVX1 U22586 ( .A(reg_file[134]), .Y(n27534) );
  MUX2X1 U22587 ( .B(n27072), .A(n25136), .S(n25847), .Y(n24993) );
  INVX1 U22588 ( .A(reg_file[135]), .Y(n27072) );
  NOR2X1 U22589 ( .A(n25847), .B(n26610), .Y(n24992) );
  INVX1 U22590 ( .A(reg_file[136]), .Y(n26610) );
  NOR2X1 U22591 ( .A(n25847), .B(n26127), .Y(n24991) );
  INVX1 U22592 ( .A(reg_file[137]), .Y(n26127) );
  NOR2X1 U22593 ( .A(n25847), .B(n31020), .Y(n24990) );
  INVX1 U22594 ( .A(reg_file[138]), .Y(n31020) );
  NOR2X1 U22595 ( .A(n25847), .B(n30558), .Y(n24989) );
  INVX1 U22596 ( .A(reg_file[139]), .Y(n30558) );
  NOR2X1 U22597 ( .A(n25847), .B(n30180), .Y(n24988) );
  INVX1 U22598 ( .A(reg_file[140]), .Y(n30180) );
  NOR2X1 U22599 ( .A(n25847), .B(n30138), .Y(n24987) );
  INVX1 U22600 ( .A(reg_file[141]), .Y(n30138) );
  NOR2X1 U22601 ( .A(n25848), .B(n30096), .Y(n24986) );
  INVX1 U22602 ( .A(reg_file[142]), .Y(n30096) );
  NOR2X1 U22603 ( .A(n25848), .B(n30054), .Y(n24985) );
  INVX1 U22604 ( .A(reg_file[143]), .Y(n30054) );
  NOR2X1 U22605 ( .A(n25848), .B(n30012), .Y(n24984) );
  INVX1 U22606 ( .A(reg_file[144]), .Y(n30012) );
  NOR2X1 U22607 ( .A(n25848), .B(n29970), .Y(n24983) );
  INVX1 U22608 ( .A(reg_file[145]), .Y(n29970) );
  NOR2X1 U22609 ( .A(n25848), .B(n29928), .Y(n24982) );
  INVX1 U22610 ( .A(reg_file[146]), .Y(n29928) );
  NOR2X1 U22611 ( .A(n25848), .B(n29886), .Y(n24981) );
  INVX1 U22612 ( .A(reg_file[147]), .Y(n29886) );
  NOR2X1 U22613 ( .A(n25848), .B(n29802), .Y(n24980) );
  INVX1 U22614 ( .A(reg_file[148]), .Y(n29802) );
  NOR2X1 U22615 ( .A(n25848), .B(n29760), .Y(n24979) );
  INVX1 U22616 ( .A(reg_file[149]), .Y(n29760) );
  NOR2X1 U22617 ( .A(n25848), .B(n29718), .Y(n24978) );
  INVX1 U22618 ( .A(reg_file[150]), .Y(n29718) );
  NOR2X1 U22619 ( .A(n25848), .B(n29676), .Y(n24977) );
  INVX1 U22620 ( .A(reg_file[151]), .Y(n29676) );
  NOR2X1 U22621 ( .A(n25848), .B(n29634), .Y(n24976) );
  INVX1 U22622 ( .A(reg_file[152]), .Y(n29634) );
  NOR2X1 U22623 ( .A(n25848), .B(n29592), .Y(n24975) );
  INVX1 U22624 ( .A(reg_file[153]), .Y(n29592) );
  NOR2X1 U22625 ( .A(n25848), .B(n29550), .Y(n24974) );
  INVX1 U22626 ( .A(reg_file[154]), .Y(n29550) );
  NOR2X1 U22627 ( .A(n25848), .B(n29508), .Y(n24973) );
  INVX1 U22628 ( .A(reg_file[155]), .Y(n29508) );
  NOR2X1 U22629 ( .A(n25848), .B(n29466), .Y(n24972) );
  INVX1 U22630 ( .A(reg_file[156]), .Y(n29466) );
  NOR2X1 U22631 ( .A(n25848), .B(n29424), .Y(n24971) );
  INVX1 U22632 ( .A(reg_file[157]), .Y(n29424) );
  NOR2X1 U22633 ( .A(n25848), .B(n29340), .Y(n24970) );
  INVX1 U22634 ( .A(reg_file[158]), .Y(n29340) );
  NOR2X1 U22635 ( .A(n25849), .B(n29298), .Y(n24969) );
  INVX1 U22636 ( .A(reg_file[159]), .Y(n29298) );
  NOR2X1 U22637 ( .A(n25849), .B(n29256), .Y(n24968) );
  INVX1 U22638 ( .A(reg_file[160]), .Y(n29256) );
  NOR2X1 U22639 ( .A(n25849), .B(n29214), .Y(n24967) );
  INVX1 U22640 ( .A(reg_file[161]), .Y(n29214) );
  NOR2X1 U22641 ( .A(n25849), .B(n29172), .Y(n24966) );
  INVX1 U22642 ( .A(reg_file[162]), .Y(n29172) );
  NOR2X1 U22643 ( .A(n25849), .B(n29130), .Y(n24965) );
  INVX1 U22644 ( .A(reg_file[163]), .Y(n29130) );
  NOR2X1 U22645 ( .A(n25849), .B(n29088), .Y(n24964) );
  INVX1 U22646 ( .A(reg_file[164]), .Y(n29088) );
  NOR2X1 U22647 ( .A(n25849), .B(n29046), .Y(n24963) );
  INVX1 U22648 ( .A(reg_file[165]), .Y(n29046) );
  NOR2X1 U22649 ( .A(n25849), .B(n29004), .Y(n24962) );
  INVX1 U22650 ( .A(reg_file[166]), .Y(n29004) );
  NOR2X1 U22651 ( .A(n25849), .B(n28962), .Y(n24961) );
  INVX1 U22652 ( .A(reg_file[167]), .Y(n28962) );
  NOR2X1 U22653 ( .A(n25849), .B(n28878), .Y(n24960) );
  INVX1 U22654 ( .A(reg_file[168]), .Y(n28878) );
  NOR2X1 U22655 ( .A(n25849), .B(n28836), .Y(n24959) );
  INVX1 U22656 ( .A(reg_file[169]), .Y(n28836) );
  NOR2X1 U22657 ( .A(n25849), .B(n28794), .Y(n24958) );
  INVX1 U22658 ( .A(reg_file[170]), .Y(n28794) );
  NOR2X1 U22659 ( .A(n25849), .B(n28752), .Y(n24957) );
  INVX1 U22660 ( .A(reg_file[171]), .Y(n28752) );
  NOR2X1 U22661 ( .A(n25849), .B(n28710), .Y(n24956) );
  INVX1 U22662 ( .A(reg_file[172]), .Y(n28710) );
  NOR2X1 U22663 ( .A(n25849), .B(n28668), .Y(n24955) );
  INVX1 U22664 ( .A(reg_file[173]), .Y(n28668) );
  NOR2X1 U22665 ( .A(n25849), .B(n28626), .Y(n24954) );
  INVX1 U22666 ( .A(reg_file[174]), .Y(n28626) );
  NOR2X1 U22667 ( .A(n25849), .B(n28584), .Y(n24953) );
  INVX1 U22668 ( .A(reg_file[175]), .Y(n28584) );
  NOR2X1 U22669 ( .A(n25850), .B(n28542), .Y(n24952) );
  INVX1 U22670 ( .A(reg_file[176]), .Y(n28542) );
  NOR2X1 U22671 ( .A(n25850), .B(n28500), .Y(n24951) );
  INVX1 U22672 ( .A(reg_file[177]), .Y(n28500) );
  NOR2X1 U22673 ( .A(n25850), .B(n28416), .Y(n24950) );
  INVX1 U22674 ( .A(reg_file[178]), .Y(n28416) );
  NOR2X1 U22675 ( .A(n25850), .B(n28374), .Y(n24949) );
  INVX1 U22676 ( .A(reg_file[179]), .Y(n28374) );
  NOR2X1 U22677 ( .A(n25850), .B(n28332), .Y(n24948) );
  INVX1 U22678 ( .A(reg_file[180]), .Y(n28332) );
  NOR2X1 U22679 ( .A(n25850), .B(n28290), .Y(n24947) );
  INVX1 U22680 ( .A(reg_file[181]), .Y(n28290) );
  NOR2X1 U22681 ( .A(n25850), .B(n28248), .Y(n24946) );
  INVX1 U22682 ( .A(reg_file[182]), .Y(n28248) );
  NOR2X1 U22683 ( .A(n25850), .B(n28206), .Y(n24945) );
  INVX1 U22684 ( .A(reg_file[183]), .Y(n28206) );
  NOR2X1 U22685 ( .A(n25850), .B(n28164), .Y(n24944) );
  INVX1 U22686 ( .A(reg_file[184]), .Y(n28164) );
  NOR2X1 U22687 ( .A(n25850), .B(n28122), .Y(n24943) );
  INVX1 U22688 ( .A(reg_file[185]), .Y(n28122) );
  NOR2X1 U22689 ( .A(n25850), .B(n28080), .Y(n24942) );
  INVX1 U22690 ( .A(reg_file[186]), .Y(n28080) );
  NOR2X1 U22691 ( .A(n25850), .B(n28038), .Y(n24941) );
  INVX1 U22692 ( .A(reg_file[187]), .Y(n28038) );
  NOR2X1 U22693 ( .A(n25850), .B(n27954), .Y(n24940) );
  INVX1 U22694 ( .A(reg_file[188]), .Y(n27954) );
  NOR2X1 U22695 ( .A(n25850), .B(n27912), .Y(n24939) );
  INVX1 U22696 ( .A(reg_file[189]), .Y(n27912) );
  NOR2X1 U22697 ( .A(n25850), .B(n27870), .Y(n24938) );
  INVX1 U22698 ( .A(reg_file[190]), .Y(n27870) );
  NOR2X1 U22699 ( .A(n25850), .B(n27828), .Y(n24937) );
  INVX1 U22700 ( .A(reg_file[191]), .Y(n27828) );
  NOR2X1 U22701 ( .A(n25850), .B(n27786), .Y(n24936) );
  INVX1 U22702 ( .A(reg_file[192]), .Y(n27786) );
  NOR2X1 U22703 ( .A(n25851), .B(n27744), .Y(n24935) );
  INVX1 U22704 ( .A(reg_file[193]), .Y(n27744) );
  NOR2X1 U22705 ( .A(n25851), .B(n27702), .Y(n24934) );
  INVX1 U22706 ( .A(reg_file[194]), .Y(n27702) );
  NOR2X1 U22707 ( .A(n25851), .B(n27660), .Y(n24933) );
  INVX1 U22708 ( .A(reg_file[195]), .Y(n27660) );
  NOR2X1 U22709 ( .A(n25851), .B(n27618), .Y(n24932) );
  INVX1 U22710 ( .A(reg_file[196]), .Y(n27618) );
  NOR2X1 U22711 ( .A(n25851), .B(n27576), .Y(n24931) );
  INVX1 U22712 ( .A(reg_file[197]), .Y(n27576) );
  NOR2X1 U22713 ( .A(n25851), .B(n27492), .Y(n24930) );
  INVX1 U22714 ( .A(reg_file[198]), .Y(n27492) );
  NOR2X1 U22715 ( .A(n25851), .B(n27450), .Y(n24929) );
  INVX1 U22716 ( .A(reg_file[199]), .Y(n27450) );
  NOR2X1 U22717 ( .A(n25851), .B(n27408), .Y(n24928) );
  INVX1 U22718 ( .A(reg_file[200]), .Y(n27408) );
  NOR2X1 U22719 ( .A(n25851), .B(n27366), .Y(n24927) );
  INVX1 U22720 ( .A(reg_file[201]), .Y(n27366) );
  NOR2X1 U22721 ( .A(n25851), .B(n27324), .Y(n24926) );
  INVX1 U22722 ( .A(reg_file[202]), .Y(n27324) );
  NOR2X1 U22723 ( .A(n25851), .B(n27282), .Y(n24925) );
  INVX1 U22724 ( .A(reg_file[203]), .Y(n27282) );
  NOR2X1 U22725 ( .A(n25851), .B(n27240), .Y(n24924) );
  INVX1 U22726 ( .A(reg_file[204]), .Y(n27240) );
  NOR2X1 U22727 ( .A(n25851), .B(n27198), .Y(n24923) );
  INVX1 U22728 ( .A(reg_file[205]), .Y(n27198) );
  NOR2X1 U22729 ( .A(n25851), .B(n27156), .Y(n24922) );
  INVX1 U22730 ( .A(reg_file[206]), .Y(n27156) );
  NOR2X1 U22731 ( .A(n25851), .B(n27114), .Y(n24921) );
  INVX1 U22732 ( .A(reg_file[207]), .Y(n27114) );
  NOR2X1 U22733 ( .A(n25851), .B(n27030), .Y(n24920) );
  INVX1 U22734 ( .A(reg_file[208]), .Y(n27030) );
  NOR2X1 U22735 ( .A(n25851), .B(n26988), .Y(n24919) );
  INVX1 U22736 ( .A(reg_file[209]), .Y(n26988) );
  NOR2X1 U22737 ( .A(n25852), .B(n26946), .Y(n24918) );
  INVX1 U22738 ( .A(reg_file[210]), .Y(n26946) );
  NOR2X1 U22739 ( .A(n25852), .B(n26904), .Y(n24917) );
  INVX1 U22740 ( .A(reg_file[211]), .Y(n26904) );
  NOR2X1 U22741 ( .A(n25852), .B(n26862), .Y(n24916) );
  INVX1 U22742 ( .A(reg_file[212]), .Y(n26862) );
  NOR2X1 U22743 ( .A(n25852), .B(n26820), .Y(n24915) );
  INVX1 U22744 ( .A(reg_file[213]), .Y(n26820) );
  NOR2X1 U22745 ( .A(n25852), .B(n26778), .Y(n24914) );
  INVX1 U22746 ( .A(reg_file[214]), .Y(n26778) );
  NOR2X1 U22747 ( .A(n25852), .B(n26736), .Y(n24913) );
  INVX1 U22748 ( .A(reg_file[215]), .Y(n26736) );
  NOR2X1 U22749 ( .A(n25852), .B(n26694), .Y(n24912) );
  INVX1 U22750 ( .A(reg_file[216]), .Y(n26694) );
  NOR2X1 U22751 ( .A(n25852), .B(n26652), .Y(n24911) );
  INVX1 U22752 ( .A(reg_file[217]), .Y(n26652) );
  NOR2X1 U22753 ( .A(n25852), .B(n26568), .Y(n24910) );
  INVX1 U22754 ( .A(reg_file[218]), .Y(n26568) );
  NOR2X1 U22755 ( .A(n25852), .B(n26526), .Y(n24909) );
  INVX1 U22756 ( .A(reg_file[219]), .Y(n26526) );
  NOR2X1 U22757 ( .A(n25852), .B(n26484), .Y(n24908) );
  INVX1 U22758 ( .A(reg_file[220]), .Y(n26484) );
  NOR2X1 U22759 ( .A(n25852), .B(n26442), .Y(n24907) );
  INVX1 U22760 ( .A(reg_file[221]), .Y(n26442) );
  NOR2X1 U22761 ( .A(n25852), .B(n26400), .Y(n24906) );
  INVX1 U22762 ( .A(reg_file[222]), .Y(n26400) );
  NOR2X1 U22763 ( .A(n25852), .B(n26358), .Y(n24905) );
  INVX1 U22764 ( .A(reg_file[223]), .Y(n26358) );
  NOR2X1 U22765 ( .A(n25852), .B(n26316), .Y(n24904) );
  INVX1 U22766 ( .A(reg_file[224]), .Y(n26316) );
  NOR2X1 U22767 ( .A(n25852), .B(n26274), .Y(n24903) );
  INVX1 U22768 ( .A(reg_file[225]), .Y(n26274) );
  NOR2X1 U22769 ( .A(n25852), .B(n26232), .Y(n24902) );
  INVX1 U22770 ( .A(reg_file[226]), .Y(n26232) );
  NOR2X1 U22771 ( .A(n25853), .B(n26190), .Y(n24901) );
  INVX1 U22772 ( .A(reg_file[227]), .Y(n26190) );
  NOR2X1 U22773 ( .A(n25853), .B(n31440), .Y(n24900) );
  INVX1 U22774 ( .A(reg_file[228]), .Y(n31440) );
  NOR2X1 U22775 ( .A(n25853), .B(n31398), .Y(n24899) );
  INVX1 U22776 ( .A(reg_file[229]), .Y(n31398) );
  NOR2X1 U22777 ( .A(n25853), .B(n31356), .Y(n24898) );
  INVX1 U22778 ( .A(reg_file[230]), .Y(n31356) );
  NOR2X1 U22779 ( .A(n25853), .B(n31314), .Y(n24897) );
  INVX1 U22780 ( .A(reg_file[231]), .Y(n31314) );
  NOR2X1 U22781 ( .A(n25853), .B(n31272), .Y(n24896) );
  INVX1 U22782 ( .A(reg_file[232]), .Y(n31272) );
  NOR2X1 U22783 ( .A(n25853), .B(n31230), .Y(n24895) );
  INVX1 U22784 ( .A(reg_file[233]), .Y(n31230) );
  NOR2X1 U22785 ( .A(n25853), .B(n31188), .Y(n24894) );
  INVX1 U22786 ( .A(reg_file[234]), .Y(n31188) );
  NOR2X1 U22787 ( .A(n25853), .B(n31146), .Y(n24893) );
  INVX1 U22788 ( .A(reg_file[235]), .Y(n31146) );
  NOR2X1 U22789 ( .A(n25853), .B(n31104), .Y(n24892) );
  INVX1 U22790 ( .A(reg_file[236]), .Y(n31104) );
  NOR2X1 U22791 ( .A(n25853), .B(n31062), .Y(n24891) );
  INVX1 U22792 ( .A(reg_file[237]), .Y(n31062) );
  NOR2X1 U22793 ( .A(n25853), .B(n30978), .Y(n24890) );
  INVX1 U22794 ( .A(reg_file[238]), .Y(n30978) );
  NOR2X1 U22795 ( .A(n25853), .B(n30936), .Y(n24889) );
  INVX1 U22796 ( .A(reg_file[239]), .Y(n30936) );
  NOR2X1 U22797 ( .A(n25853), .B(n30894), .Y(n24888) );
  INVX1 U22798 ( .A(reg_file[240]), .Y(n30894) );
  NOR2X1 U22799 ( .A(n25853), .B(n30852), .Y(n24887) );
  INVX1 U22800 ( .A(reg_file[241]), .Y(n30852) );
  NOR2X1 U22801 ( .A(n25853), .B(n30810), .Y(n24886) );
  INVX1 U22802 ( .A(reg_file[242]), .Y(n30810) );
  NOR2X1 U22803 ( .A(n25853), .B(n30768), .Y(n24885) );
  INVX1 U22804 ( .A(reg_file[243]), .Y(n30768) );
  NOR2X1 U22805 ( .A(n25854), .B(n30726), .Y(n24884) );
  INVX1 U22806 ( .A(reg_file[244]), .Y(n30726) );
  NOR2X1 U22807 ( .A(n25854), .B(n30684), .Y(n24883) );
  INVX1 U22808 ( .A(reg_file[245]), .Y(n30684) );
  NOR2X1 U22809 ( .A(n25854), .B(n30642), .Y(n24882) );
  INVX1 U22810 ( .A(reg_file[246]), .Y(n30642) );
  NOR2X1 U22811 ( .A(n25854), .B(n30600), .Y(n24881) );
  INVX1 U22812 ( .A(reg_file[247]), .Y(n30600) );
  NOR2X1 U22813 ( .A(n25854), .B(n30516), .Y(n24880) );
  INVX1 U22814 ( .A(reg_file[248]), .Y(n30516) );
  NOR2X1 U22815 ( .A(n25854), .B(n30474), .Y(n24879) );
  INVX1 U22816 ( .A(reg_file[249]), .Y(n30474) );
  NOR2X1 U22817 ( .A(n25854), .B(n30432), .Y(n24878) );
  INVX1 U22818 ( .A(reg_file[250]), .Y(n30432) );
  NOR2X1 U22819 ( .A(n25854), .B(n30390), .Y(n24877) );
  INVX1 U22820 ( .A(reg_file[251]), .Y(n30390) );
  NOR2X1 U22821 ( .A(n25854), .B(n30348), .Y(n24876) );
  INVX1 U22822 ( .A(reg_file[252]), .Y(n30348) );
  NOR2X1 U22823 ( .A(n25854), .B(n30306), .Y(n24875) );
  INVX1 U22824 ( .A(reg_file[253]), .Y(n30306) );
  NOR2X1 U22825 ( .A(n25854), .B(n30264), .Y(n24874) );
  INVX1 U22826 ( .A(reg_file[254]), .Y(n30264) );
  NOR2X1 U22827 ( .A(n25854), .B(n30222), .Y(n24873) );
  INVX1 U22828 ( .A(reg_file[255]), .Y(n30222) );
  NOR2X1 U22829 ( .A(n34925), .B(n34923), .Y(n34924) );
  MUX2X1 U22830 ( .B(n31491), .A(n25129), .S(n25855), .Y(n24872) );
  INVX1 U22831 ( .A(reg_file[256]), .Y(n31491) );
  MUX2X1 U22832 ( .B(n29843), .A(n25130), .S(n25855), .Y(n24871) );
  INVX1 U22833 ( .A(reg_file[257]), .Y(n29843) );
  MUX2X1 U22834 ( .B(n29381), .A(n25131), .S(n25855), .Y(n24870) );
  INVX1 U22835 ( .A(reg_file[258]), .Y(n29381) );
  MUX2X1 U22836 ( .B(n28919), .A(n25132), .S(n25855), .Y(n24869) );
  INVX1 U22837 ( .A(reg_file[259]), .Y(n28919) );
  MUX2X1 U22838 ( .B(n28457), .A(n25133), .S(n25855), .Y(n24868) );
  INVX1 U22839 ( .A(reg_file[260]), .Y(n28457) );
  MUX2X1 U22840 ( .B(n27995), .A(n25134), .S(n25855), .Y(n24867) );
  INVX1 U22841 ( .A(reg_file[261]), .Y(n27995) );
  MUX2X1 U22842 ( .B(n27533), .A(n25135), .S(n25855), .Y(n24866) );
  INVX1 U22843 ( .A(reg_file[262]), .Y(n27533) );
  MUX2X1 U22844 ( .B(n27071), .A(n25136), .S(n25855), .Y(n24865) );
  INVX1 U22845 ( .A(reg_file[263]), .Y(n27071) );
  NOR2X1 U22846 ( .A(n25855), .B(n26609), .Y(n24864) );
  INVX1 U22847 ( .A(reg_file[264]), .Y(n26609) );
  NOR2X1 U22848 ( .A(n25855), .B(n26125), .Y(n24863) );
  INVX1 U22849 ( .A(reg_file[265]), .Y(n26125) );
  NOR2X1 U22850 ( .A(n25855), .B(n31019), .Y(n24862) );
  INVX1 U22851 ( .A(reg_file[266]), .Y(n31019) );
  NOR2X1 U22852 ( .A(n25855), .B(n30557), .Y(n24861) );
  INVX1 U22853 ( .A(reg_file[267]), .Y(n30557) );
  NOR2X1 U22854 ( .A(n25855), .B(n30179), .Y(n24860) );
  INVX1 U22855 ( .A(reg_file[268]), .Y(n30179) );
  NOR2X1 U22856 ( .A(n25855), .B(n30137), .Y(n24859) );
  INVX1 U22857 ( .A(reg_file[269]), .Y(n30137) );
  NOR2X1 U22858 ( .A(n25856), .B(n30095), .Y(n24858) );
  INVX1 U22859 ( .A(reg_file[270]), .Y(n30095) );
  NOR2X1 U22860 ( .A(n25856), .B(n30053), .Y(n24857) );
  INVX1 U22861 ( .A(reg_file[271]), .Y(n30053) );
  NOR2X1 U22862 ( .A(n25856), .B(n30011), .Y(n24856) );
  INVX1 U22863 ( .A(reg_file[272]), .Y(n30011) );
  NOR2X1 U22864 ( .A(n25856), .B(n29969), .Y(n24855) );
  INVX1 U22865 ( .A(reg_file[273]), .Y(n29969) );
  NOR2X1 U22866 ( .A(n25856), .B(n29927), .Y(n24854) );
  INVX1 U22867 ( .A(reg_file[274]), .Y(n29927) );
  NOR2X1 U22868 ( .A(n25856), .B(n29885), .Y(n24853) );
  INVX1 U22869 ( .A(reg_file[275]), .Y(n29885) );
  NOR2X1 U22870 ( .A(n25856), .B(n29801), .Y(n24852) );
  INVX1 U22871 ( .A(reg_file[276]), .Y(n29801) );
  NOR2X1 U22872 ( .A(n25856), .B(n29759), .Y(n24851) );
  INVX1 U22873 ( .A(reg_file[277]), .Y(n29759) );
  NOR2X1 U22874 ( .A(n25856), .B(n29717), .Y(n24850) );
  INVX1 U22875 ( .A(reg_file[278]), .Y(n29717) );
  NOR2X1 U22876 ( .A(n25856), .B(n29675), .Y(n24849) );
  INVX1 U22877 ( .A(reg_file[279]), .Y(n29675) );
  NOR2X1 U22878 ( .A(n25856), .B(n29633), .Y(n24848) );
  INVX1 U22879 ( .A(reg_file[280]), .Y(n29633) );
  NOR2X1 U22880 ( .A(n25856), .B(n29591), .Y(n24847) );
  INVX1 U22881 ( .A(reg_file[281]), .Y(n29591) );
  NOR2X1 U22882 ( .A(n25856), .B(n29549), .Y(n24846) );
  INVX1 U22883 ( .A(reg_file[282]), .Y(n29549) );
  NOR2X1 U22884 ( .A(n25856), .B(n29507), .Y(n24845) );
  INVX1 U22885 ( .A(reg_file[283]), .Y(n29507) );
  NOR2X1 U22886 ( .A(n25856), .B(n29465), .Y(n24844) );
  INVX1 U22887 ( .A(reg_file[284]), .Y(n29465) );
  NOR2X1 U22888 ( .A(n25856), .B(n29423), .Y(n24843) );
  INVX1 U22889 ( .A(reg_file[285]), .Y(n29423) );
  NOR2X1 U22890 ( .A(n25856), .B(n29339), .Y(n24842) );
  INVX1 U22891 ( .A(reg_file[286]), .Y(n29339) );
  NOR2X1 U22892 ( .A(n25857), .B(n29297), .Y(n24841) );
  INVX1 U22893 ( .A(reg_file[287]), .Y(n29297) );
  NOR2X1 U22894 ( .A(n25857), .B(n29255), .Y(n24840) );
  INVX1 U22895 ( .A(reg_file[288]), .Y(n29255) );
  NOR2X1 U22896 ( .A(n25857), .B(n29213), .Y(n24839) );
  INVX1 U22897 ( .A(reg_file[289]), .Y(n29213) );
  NOR2X1 U22898 ( .A(n25857), .B(n29171), .Y(n24838) );
  INVX1 U22899 ( .A(reg_file[290]), .Y(n29171) );
  NOR2X1 U22900 ( .A(n25857), .B(n29129), .Y(n24837) );
  INVX1 U22901 ( .A(reg_file[291]), .Y(n29129) );
  NOR2X1 U22902 ( .A(n25857), .B(n29087), .Y(n24836) );
  INVX1 U22903 ( .A(reg_file[292]), .Y(n29087) );
  NOR2X1 U22904 ( .A(n25857), .B(n29045), .Y(n24835) );
  INVX1 U22905 ( .A(reg_file[293]), .Y(n29045) );
  NOR2X1 U22906 ( .A(n25857), .B(n29003), .Y(n24834) );
  INVX1 U22907 ( .A(reg_file[294]), .Y(n29003) );
  NOR2X1 U22908 ( .A(n25857), .B(n28961), .Y(n24833) );
  INVX1 U22909 ( .A(reg_file[295]), .Y(n28961) );
  NOR2X1 U22910 ( .A(n25857), .B(n28877), .Y(n24832) );
  INVX1 U22911 ( .A(reg_file[296]), .Y(n28877) );
  NOR2X1 U22912 ( .A(n25857), .B(n28835), .Y(n24831) );
  INVX1 U22913 ( .A(reg_file[297]), .Y(n28835) );
  NOR2X1 U22914 ( .A(n25857), .B(n28793), .Y(n24830) );
  INVX1 U22915 ( .A(reg_file[298]), .Y(n28793) );
  NOR2X1 U22916 ( .A(n25857), .B(n28751), .Y(n24829) );
  INVX1 U22917 ( .A(reg_file[299]), .Y(n28751) );
  NOR2X1 U22918 ( .A(n25857), .B(n28709), .Y(n24828) );
  INVX1 U22919 ( .A(reg_file[300]), .Y(n28709) );
  NOR2X1 U22920 ( .A(n25857), .B(n28667), .Y(n24827) );
  INVX1 U22921 ( .A(reg_file[301]), .Y(n28667) );
  NOR2X1 U22922 ( .A(n25857), .B(n28625), .Y(n24826) );
  INVX1 U22923 ( .A(reg_file[302]), .Y(n28625) );
  NOR2X1 U22924 ( .A(n25857), .B(n28583), .Y(n24825) );
  INVX1 U22925 ( .A(reg_file[303]), .Y(n28583) );
  NOR2X1 U22926 ( .A(n25858), .B(n28541), .Y(n24824) );
  INVX1 U22927 ( .A(reg_file[304]), .Y(n28541) );
  NOR2X1 U22928 ( .A(n25858), .B(n28499), .Y(n24823) );
  INVX1 U22929 ( .A(reg_file[305]), .Y(n28499) );
  NOR2X1 U22930 ( .A(n25858), .B(n28415), .Y(n24822) );
  INVX1 U22931 ( .A(reg_file[306]), .Y(n28415) );
  NOR2X1 U22932 ( .A(n25858), .B(n28373), .Y(n24821) );
  INVX1 U22933 ( .A(reg_file[307]), .Y(n28373) );
  NOR2X1 U22934 ( .A(n25858), .B(n28331), .Y(n24820) );
  INVX1 U22935 ( .A(reg_file[308]), .Y(n28331) );
  NOR2X1 U22936 ( .A(n25858), .B(n28289), .Y(n24819) );
  INVX1 U22937 ( .A(reg_file[309]), .Y(n28289) );
  NOR2X1 U22938 ( .A(n25858), .B(n28247), .Y(n24818) );
  INVX1 U22939 ( .A(reg_file[310]), .Y(n28247) );
  NOR2X1 U22940 ( .A(n25858), .B(n28205), .Y(n24817) );
  INVX1 U22941 ( .A(reg_file[311]), .Y(n28205) );
  NOR2X1 U22942 ( .A(n25858), .B(n28163), .Y(n24816) );
  INVX1 U22943 ( .A(reg_file[312]), .Y(n28163) );
  NOR2X1 U22944 ( .A(n25858), .B(n28121), .Y(n24815) );
  INVX1 U22945 ( .A(reg_file[313]), .Y(n28121) );
  NOR2X1 U22946 ( .A(n25858), .B(n28079), .Y(n24814) );
  INVX1 U22947 ( .A(reg_file[314]), .Y(n28079) );
  NOR2X1 U22948 ( .A(n25858), .B(n28037), .Y(n24813) );
  INVX1 U22949 ( .A(reg_file[315]), .Y(n28037) );
  NOR2X1 U22950 ( .A(n25858), .B(n27953), .Y(n24812) );
  INVX1 U22951 ( .A(reg_file[316]), .Y(n27953) );
  NOR2X1 U22952 ( .A(n25858), .B(n27911), .Y(n24811) );
  INVX1 U22953 ( .A(reg_file[317]), .Y(n27911) );
  NOR2X1 U22954 ( .A(n25858), .B(n27869), .Y(n24810) );
  INVX1 U22955 ( .A(reg_file[318]), .Y(n27869) );
  NOR2X1 U22956 ( .A(n25858), .B(n27827), .Y(n24809) );
  INVX1 U22957 ( .A(reg_file[319]), .Y(n27827) );
  NOR2X1 U22958 ( .A(n25858), .B(n27785), .Y(n24808) );
  INVX1 U22959 ( .A(reg_file[320]), .Y(n27785) );
  NOR2X1 U22960 ( .A(n25859), .B(n27743), .Y(n24807) );
  INVX1 U22961 ( .A(reg_file[321]), .Y(n27743) );
  NOR2X1 U22962 ( .A(n25859), .B(n27701), .Y(n24806) );
  INVX1 U22963 ( .A(reg_file[322]), .Y(n27701) );
  NOR2X1 U22964 ( .A(n25859), .B(n27659), .Y(n24805) );
  INVX1 U22965 ( .A(reg_file[323]), .Y(n27659) );
  NOR2X1 U22966 ( .A(n25859), .B(n27617), .Y(n24804) );
  INVX1 U22967 ( .A(reg_file[324]), .Y(n27617) );
  NOR2X1 U22968 ( .A(n25859), .B(n27575), .Y(n24803) );
  INVX1 U22969 ( .A(reg_file[325]), .Y(n27575) );
  NOR2X1 U22970 ( .A(n25859), .B(n27491), .Y(n24802) );
  INVX1 U22971 ( .A(reg_file[326]), .Y(n27491) );
  NOR2X1 U22972 ( .A(n25859), .B(n27449), .Y(n24801) );
  INVX1 U22973 ( .A(reg_file[327]), .Y(n27449) );
  NOR2X1 U22974 ( .A(n25859), .B(n27407), .Y(n24800) );
  INVX1 U22975 ( .A(reg_file[328]), .Y(n27407) );
  NOR2X1 U22976 ( .A(n25859), .B(n27365), .Y(n24799) );
  INVX1 U22977 ( .A(reg_file[329]), .Y(n27365) );
  NOR2X1 U22978 ( .A(n25859), .B(n27323), .Y(n24798) );
  INVX1 U22979 ( .A(reg_file[330]), .Y(n27323) );
  NOR2X1 U22980 ( .A(n25859), .B(n27281), .Y(n24797) );
  INVX1 U22981 ( .A(reg_file[331]), .Y(n27281) );
  NOR2X1 U22982 ( .A(n25859), .B(n27239), .Y(n24796) );
  INVX1 U22983 ( .A(reg_file[332]), .Y(n27239) );
  NOR2X1 U22984 ( .A(n25859), .B(n27197), .Y(n24795) );
  INVX1 U22985 ( .A(reg_file[333]), .Y(n27197) );
  NOR2X1 U22986 ( .A(n25859), .B(n27155), .Y(n24794) );
  INVX1 U22987 ( .A(reg_file[334]), .Y(n27155) );
  NOR2X1 U22988 ( .A(n25859), .B(n27113), .Y(n24793) );
  INVX1 U22989 ( .A(reg_file[335]), .Y(n27113) );
  NOR2X1 U22990 ( .A(n25859), .B(n27029), .Y(n24792) );
  INVX1 U22991 ( .A(reg_file[336]), .Y(n27029) );
  NOR2X1 U22992 ( .A(n25859), .B(n26987), .Y(n24791) );
  INVX1 U22993 ( .A(reg_file[337]), .Y(n26987) );
  NOR2X1 U22994 ( .A(n25860), .B(n26945), .Y(n24790) );
  INVX1 U22995 ( .A(reg_file[338]), .Y(n26945) );
  NOR2X1 U22996 ( .A(n25860), .B(n26903), .Y(n24789) );
  INVX1 U22997 ( .A(reg_file[339]), .Y(n26903) );
  NOR2X1 U22998 ( .A(n25860), .B(n26861), .Y(n24788) );
  INVX1 U22999 ( .A(reg_file[340]), .Y(n26861) );
  NOR2X1 U23000 ( .A(n25860), .B(n26819), .Y(n24787) );
  INVX1 U23001 ( .A(reg_file[341]), .Y(n26819) );
  NOR2X1 U23002 ( .A(n25860), .B(n26777), .Y(n24786) );
  INVX1 U23003 ( .A(reg_file[342]), .Y(n26777) );
  NOR2X1 U23004 ( .A(n25860), .B(n26735), .Y(n24785) );
  INVX1 U23005 ( .A(reg_file[343]), .Y(n26735) );
  NOR2X1 U23006 ( .A(n25860), .B(n26693), .Y(n24784) );
  INVX1 U23007 ( .A(reg_file[344]), .Y(n26693) );
  NOR2X1 U23008 ( .A(n25860), .B(n26651), .Y(n24783) );
  INVX1 U23009 ( .A(reg_file[345]), .Y(n26651) );
  NOR2X1 U23010 ( .A(n25860), .B(n26567), .Y(n24782) );
  INVX1 U23011 ( .A(reg_file[346]), .Y(n26567) );
  NOR2X1 U23012 ( .A(n25860), .B(n26525), .Y(n24781) );
  INVX1 U23013 ( .A(reg_file[347]), .Y(n26525) );
  NOR2X1 U23014 ( .A(n25860), .B(n26483), .Y(n24780) );
  INVX1 U23015 ( .A(reg_file[348]), .Y(n26483) );
  NOR2X1 U23016 ( .A(n25860), .B(n26441), .Y(n24779) );
  INVX1 U23017 ( .A(reg_file[349]), .Y(n26441) );
  NOR2X1 U23018 ( .A(n25860), .B(n26399), .Y(n24778) );
  INVX1 U23019 ( .A(reg_file[350]), .Y(n26399) );
  NOR2X1 U23020 ( .A(n25860), .B(n26357), .Y(n24777) );
  INVX1 U23021 ( .A(reg_file[351]), .Y(n26357) );
  NOR2X1 U23022 ( .A(n25860), .B(n26315), .Y(n24776) );
  INVX1 U23023 ( .A(reg_file[352]), .Y(n26315) );
  NOR2X1 U23024 ( .A(n25860), .B(n26273), .Y(n24775) );
  INVX1 U23025 ( .A(reg_file[353]), .Y(n26273) );
  NOR2X1 U23026 ( .A(n25860), .B(n26231), .Y(n24774) );
  INVX1 U23027 ( .A(reg_file[354]), .Y(n26231) );
  NOR2X1 U23028 ( .A(n25861), .B(n26189), .Y(n24773) );
  INVX1 U23029 ( .A(reg_file[355]), .Y(n26189) );
  NOR2X1 U23030 ( .A(n25861), .B(n31439), .Y(n24772) );
  INVX1 U23031 ( .A(reg_file[356]), .Y(n31439) );
  NOR2X1 U23032 ( .A(n25861), .B(n31397), .Y(n24771) );
  INVX1 U23033 ( .A(reg_file[357]), .Y(n31397) );
  NOR2X1 U23034 ( .A(n25861), .B(n31355), .Y(n24770) );
  INVX1 U23035 ( .A(reg_file[358]), .Y(n31355) );
  NOR2X1 U23036 ( .A(n25861), .B(n31313), .Y(n24769) );
  INVX1 U23037 ( .A(reg_file[359]), .Y(n31313) );
  NOR2X1 U23038 ( .A(n25861), .B(n31271), .Y(n24768) );
  INVX1 U23039 ( .A(reg_file[360]), .Y(n31271) );
  NOR2X1 U23040 ( .A(n25861), .B(n31229), .Y(n24767) );
  INVX1 U23041 ( .A(reg_file[361]), .Y(n31229) );
  NOR2X1 U23042 ( .A(n25861), .B(n31187), .Y(n24766) );
  INVX1 U23043 ( .A(reg_file[362]), .Y(n31187) );
  NOR2X1 U23044 ( .A(n25861), .B(n31145), .Y(n24765) );
  INVX1 U23045 ( .A(reg_file[363]), .Y(n31145) );
  NOR2X1 U23046 ( .A(n25861), .B(n31103), .Y(n24764) );
  INVX1 U23047 ( .A(reg_file[364]), .Y(n31103) );
  NOR2X1 U23048 ( .A(n25861), .B(n31061), .Y(n24763) );
  INVX1 U23049 ( .A(reg_file[365]), .Y(n31061) );
  NOR2X1 U23050 ( .A(n25861), .B(n30977), .Y(n24762) );
  INVX1 U23051 ( .A(reg_file[366]), .Y(n30977) );
  NOR2X1 U23052 ( .A(n25861), .B(n30935), .Y(n24761) );
  INVX1 U23053 ( .A(reg_file[367]), .Y(n30935) );
  NOR2X1 U23054 ( .A(n25861), .B(n30893), .Y(n24760) );
  INVX1 U23055 ( .A(reg_file[368]), .Y(n30893) );
  NOR2X1 U23056 ( .A(n25861), .B(n30851), .Y(n24759) );
  INVX1 U23057 ( .A(reg_file[369]), .Y(n30851) );
  NOR2X1 U23058 ( .A(n25861), .B(n30809), .Y(n24758) );
  INVX1 U23059 ( .A(reg_file[370]), .Y(n30809) );
  NOR2X1 U23060 ( .A(n25861), .B(n30767), .Y(n24757) );
  INVX1 U23061 ( .A(reg_file[371]), .Y(n30767) );
  NOR2X1 U23062 ( .A(n25862), .B(n30725), .Y(n24756) );
  INVX1 U23063 ( .A(reg_file[372]), .Y(n30725) );
  NOR2X1 U23064 ( .A(n25862), .B(n30683), .Y(n24755) );
  INVX1 U23065 ( .A(reg_file[373]), .Y(n30683) );
  NOR2X1 U23066 ( .A(n25862), .B(n30641), .Y(n24754) );
  INVX1 U23067 ( .A(reg_file[374]), .Y(n30641) );
  NOR2X1 U23068 ( .A(n25862), .B(n30599), .Y(n24753) );
  INVX1 U23069 ( .A(reg_file[375]), .Y(n30599) );
  NOR2X1 U23070 ( .A(n25862), .B(n30515), .Y(n24752) );
  INVX1 U23071 ( .A(reg_file[376]), .Y(n30515) );
  NOR2X1 U23072 ( .A(n25862), .B(n30473), .Y(n24751) );
  INVX1 U23073 ( .A(reg_file[377]), .Y(n30473) );
  NOR2X1 U23074 ( .A(n25862), .B(n30431), .Y(n24750) );
  INVX1 U23075 ( .A(reg_file[378]), .Y(n30431) );
  NOR2X1 U23076 ( .A(n25862), .B(n30389), .Y(n24749) );
  INVX1 U23077 ( .A(reg_file[379]), .Y(n30389) );
  NOR2X1 U23078 ( .A(n25862), .B(n30347), .Y(n24748) );
  INVX1 U23079 ( .A(reg_file[380]), .Y(n30347) );
  NOR2X1 U23080 ( .A(n25862), .B(n30305), .Y(n24747) );
  INVX1 U23081 ( .A(reg_file[381]), .Y(n30305) );
  NOR2X1 U23082 ( .A(n25862), .B(n30263), .Y(n24746) );
  INVX1 U23083 ( .A(reg_file[382]), .Y(n30263) );
  NOR2X1 U23084 ( .A(n25862), .B(n30221), .Y(n24745) );
  INVX1 U23085 ( .A(reg_file[383]), .Y(n30221) );
  NOR2X1 U23086 ( .A(n34927), .B(n34922), .Y(n34926) );
  MUX2X1 U23087 ( .B(n31490), .A(n25129), .S(n25863), .Y(n24744) );
  INVX1 U23088 ( .A(reg_file[384]), .Y(n31490) );
  MUX2X1 U23089 ( .B(n29842), .A(n25130), .S(n25863), .Y(n24743) );
  INVX1 U23090 ( .A(reg_file[385]), .Y(n29842) );
  MUX2X1 U23091 ( .B(n29380), .A(n25131), .S(n25863), .Y(n24742) );
  INVX1 U23092 ( .A(reg_file[386]), .Y(n29380) );
  MUX2X1 U23093 ( .B(n28918), .A(n25132), .S(n25863), .Y(n24741) );
  INVX1 U23094 ( .A(reg_file[387]), .Y(n28918) );
  MUX2X1 U23095 ( .B(n28456), .A(n25133), .S(n25863), .Y(n24740) );
  INVX1 U23096 ( .A(reg_file[388]), .Y(n28456) );
  MUX2X1 U23097 ( .B(n27994), .A(n25134), .S(n25863), .Y(n24739) );
  INVX1 U23098 ( .A(reg_file[389]), .Y(n27994) );
  MUX2X1 U23099 ( .B(n27532), .A(n25135), .S(n25863), .Y(n24738) );
  INVX1 U23100 ( .A(reg_file[390]), .Y(n27532) );
  MUX2X1 U23101 ( .B(n27070), .A(n25136), .S(n25863), .Y(n24737) );
  INVX1 U23102 ( .A(reg_file[391]), .Y(n27070) );
  NOR2X1 U23103 ( .A(n25863), .B(n26608), .Y(n24736) );
  INVX1 U23104 ( .A(reg_file[392]), .Y(n26608) );
  NOR2X1 U23105 ( .A(n25863), .B(n26123), .Y(n24735) );
  INVX1 U23106 ( .A(reg_file[393]), .Y(n26123) );
  NOR2X1 U23107 ( .A(n25863), .B(n31018), .Y(n24734) );
  INVX1 U23108 ( .A(reg_file[394]), .Y(n31018) );
  NOR2X1 U23109 ( .A(n25863), .B(n30556), .Y(n24733) );
  INVX1 U23110 ( .A(reg_file[395]), .Y(n30556) );
  NOR2X1 U23111 ( .A(n25863), .B(n30178), .Y(n24732) );
  INVX1 U23112 ( .A(reg_file[396]), .Y(n30178) );
  NOR2X1 U23113 ( .A(n25863), .B(n30136), .Y(n24731) );
  INVX1 U23114 ( .A(reg_file[397]), .Y(n30136) );
  NOR2X1 U23115 ( .A(n25864), .B(n30094), .Y(n24730) );
  INVX1 U23116 ( .A(reg_file[398]), .Y(n30094) );
  NOR2X1 U23117 ( .A(n25864), .B(n30052), .Y(n24729) );
  INVX1 U23118 ( .A(reg_file[399]), .Y(n30052) );
  NOR2X1 U23119 ( .A(n25864), .B(n30010), .Y(n24728) );
  INVX1 U23120 ( .A(reg_file[400]), .Y(n30010) );
  NOR2X1 U23121 ( .A(n25864), .B(n29968), .Y(n24727) );
  INVX1 U23122 ( .A(reg_file[401]), .Y(n29968) );
  NOR2X1 U23123 ( .A(n25864), .B(n29926), .Y(n24726) );
  INVX1 U23124 ( .A(reg_file[402]), .Y(n29926) );
  NOR2X1 U23125 ( .A(n25864), .B(n29884), .Y(n24725) );
  INVX1 U23126 ( .A(reg_file[403]), .Y(n29884) );
  NOR2X1 U23127 ( .A(n25864), .B(n29800), .Y(n24724) );
  INVX1 U23128 ( .A(reg_file[404]), .Y(n29800) );
  NOR2X1 U23129 ( .A(n25864), .B(n29758), .Y(n24723) );
  INVX1 U23130 ( .A(reg_file[405]), .Y(n29758) );
  NOR2X1 U23131 ( .A(n25864), .B(n29716), .Y(n24722) );
  INVX1 U23132 ( .A(reg_file[406]), .Y(n29716) );
  NOR2X1 U23133 ( .A(n25864), .B(n29674), .Y(n24721) );
  INVX1 U23134 ( .A(reg_file[407]), .Y(n29674) );
  NOR2X1 U23135 ( .A(n25864), .B(n29632), .Y(n24720) );
  INVX1 U23136 ( .A(reg_file[408]), .Y(n29632) );
  NOR2X1 U23137 ( .A(n25864), .B(n29590), .Y(n24719) );
  INVX1 U23138 ( .A(reg_file[409]), .Y(n29590) );
  NOR2X1 U23139 ( .A(n25864), .B(n29548), .Y(n24718) );
  INVX1 U23140 ( .A(reg_file[410]), .Y(n29548) );
  NOR2X1 U23141 ( .A(n25864), .B(n29506), .Y(n24717) );
  INVX1 U23142 ( .A(reg_file[411]), .Y(n29506) );
  NOR2X1 U23143 ( .A(n25864), .B(n29464), .Y(n24716) );
  INVX1 U23144 ( .A(reg_file[412]), .Y(n29464) );
  NOR2X1 U23145 ( .A(n25864), .B(n29422), .Y(n24715) );
  INVX1 U23146 ( .A(reg_file[413]), .Y(n29422) );
  NOR2X1 U23147 ( .A(n25864), .B(n29338), .Y(n24714) );
  INVX1 U23148 ( .A(reg_file[414]), .Y(n29338) );
  NOR2X1 U23149 ( .A(n25865), .B(n29296), .Y(n24713) );
  INVX1 U23150 ( .A(reg_file[415]), .Y(n29296) );
  NOR2X1 U23151 ( .A(n25865), .B(n29254), .Y(n24712) );
  INVX1 U23152 ( .A(reg_file[416]), .Y(n29254) );
  NOR2X1 U23153 ( .A(n25865), .B(n29212), .Y(n24711) );
  INVX1 U23154 ( .A(reg_file[417]), .Y(n29212) );
  NOR2X1 U23155 ( .A(n25865), .B(n29170), .Y(n24710) );
  INVX1 U23156 ( .A(reg_file[418]), .Y(n29170) );
  NOR2X1 U23157 ( .A(n25865), .B(n29128), .Y(n24709) );
  INVX1 U23158 ( .A(reg_file[419]), .Y(n29128) );
  NOR2X1 U23159 ( .A(n25865), .B(n29086), .Y(n24708) );
  INVX1 U23160 ( .A(reg_file[420]), .Y(n29086) );
  NOR2X1 U23161 ( .A(n25865), .B(n29044), .Y(n24707) );
  INVX1 U23162 ( .A(reg_file[421]), .Y(n29044) );
  NOR2X1 U23163 ( .A(n25865), .B(n29002), .Y(n24706) );
  INVX1 U23164 ( .A(reg_file[422]), .Y(n29002) );
  NOR2X1 U23165 ( .A(n25865), .B(n28960), .Y(n24705) );
  INVX1 U23166 ( .A(reg_file[423]), .Y(n28960) );
  NOR2X1 U23167 ( .A(n25865), .B(n28876), .Y(n24704) );
  INVX1 U23168 ( .A(reg_file[424]), .Y(n28876) );
  NOR2X1 U23169 ( .A(n25865), .B(n28834), .Y(n24703) );
  INVX1 U23170 ( .A(reg_file[425]), .Y(n28834) );
  NOR2X1 U23171 ( .A(n25865), .B(n28792), .Y(n24702) );
  INVX1 U23172 ( .A(reg_file[426]), .Y(n28792) );
  NOR2X1 U23173 ( .A(n25865), .B(n28750), .Y(n24701) );
  INVX1 U23174 ( .A(reg_file[427]), .Y(n28750) );
  NOR2X1 U23175 ( .A(n25865), .B(n28708), .Y(n24700) );
  INVX1 U23176 ( .A(reg_file[428]), .Y(n28708) );
  NOR2X1 U23177 ( .A(n25865), .B(n28666), .Y(n24699) );
  INVX1 U23178 ( .A(reg_file[429]), .Y(n28666) );
  NOR2X1 U23179 ( .A(n25865), .B(n28624), .Y(n24698) );
  INVX1 U23180 ( .A(reg_file[430]), .Y(n28624) );
  NOR2X1 U23181 ( .A(n25865), .B(n28582), .Y(n24697) );
  INVX1 U23182 ( .A(reg_file[431]), .Y(n28582) );
  NOR2X1 U23183 ( .A(n25866), .B(n28540), .Y(n24696) );
  INVX1 U23184 ( .A(reg_file[432]), .Y(n28540) );
  NOR2X1 U23185 ( .A(n25866), .B(n28498), .Y(n24695) );
  INVX1 U23186 ( .A(reg_file[433]), .Y(n28498) );
  NOR2X1 U23187 ( .A(n25866), .B(n28414), .Y(n24694) );
  INVX1 U23188 ( .A(reg_file[434]), .Y(n28414) );
  NOR2X1 U23189 ( .A(n25866), .B(n28372), .Y(n24693) );
  INVX1 U23190 ( .A(reg_file[435]), .Y(n28372) );
  NOR2X1 U23191 ( .A(n25866), .B(n28330), .Y(n24692) );
  INVX1 U23192 ( .A(reg_file[436]), .Y(n28330) );
  NOR2X1 U23193 ( .A(n25866), .B(n28288), .Y(n24691) );
  INVX1 U23194 ( .A(reg_file[437]), .Y(n28288) );
  NOR2X1 U23195 ( .A(n25866), .B(n28246), .Y(n24690) );
  INVX1 U23196 ( .A(reg_file[438]), .Y(n28246) );
  NOR2X1 U23197 ( .A(n25866), .B(n28204), .Y(n24689) );
  INVX1 U23198 ( .A(reg_file[439]), .Y(n28204) );
  NOR2X1 U23199 ( .A(n25866), .B(n28162), .Y(n24688) );
  INVX1 U23200 ( .A(reg_file[440]), .Y(n28162) );
  NOR2X1 U23201 ( .A(n25866), .B(n28120), .Y(n24687) );
  INVX1 U23202 ( .A(reg_file[441]), .Y(n28120) );
  NOR2X1 U23203 ( .A(n25866), .B(n28078), .Y(n24686) );
  INVX1 U23204 ( .A(reg_file[442]), .Y(n28078) );
  NOR2X1 U23205 ( .A(n25866), .B(n28036), .Y(n24685) );
  INVX1 U23206 ( .A(reg_file[443]), .Y(n28036) );
  NOR2X1 U23207 ( .A(n25866), .B(n27952), .Y(n24684) );
  INVX1 U23208 ( .A(reg_file[444]), .Y(n27952) );
  NOR2X1 U23209 ( .A(n25866), .B(n27910), .Y(n24683) );
  INVX1 U23210 ( .A(reg_file[445]), .Y(n27910) );
  NOR2X1 U23211 ( .A(n25866), .B(n27868), .Y(n24682) );
  INVX1 U23212 ( .A(reg_file[446]), .Y(n27868) );
  NOR2X1 U23213 ( .A(n25866), .B(n27826), .Y(n24681) );
  INVX1 U23214 ( .A(reg_file[447]), .Y(n27826) );
  NOR2X1 U23215 ( .A(n25866), .B(n27784), .Y(n24680) );
  INVX1 U23216 ( .A(reg_file[448]), .Y(n27784) );
  NOR2X1 U23217 ( .A(n25867), .B(n27742), .Y(n24679) );
  INVX1 U23218 ( .A(reg_file[449]), .Y(n27742) );
  NOR2X1 U23219 ( .A(n25867), .B(n27700), .Y(n24678) );
  INVX1 U23220 ( .A(reg_file[450]), .Y(n27700) );
  NOR2X1 U23221 ( .A(n25867), .B(n27658), .Y(n24677) );
  INVX1 U23222 ( .A(reg_file[451]), .Y(n27658) );
  NOR2X1 U23223 ( .A(n25867), .B(n27616), .Y(n24676) );
  INVX1 U23224 ( .A(reg_file[452]), .Y(n27616) );
  NOR2X1 U23225 ( .A(n25867), .B(n27574), .Y(n24675) );
  INVX1 U23226 ( .A(reg_file[453]), .Y(n27574) );
  NOR2X1 U23227 ( .A(n25867), .B(n27490), .Y(n24674) );
  INVX1 U23228 ( .A(reg_file[454]), .Y(n27490) );
  NOR2X1 U23229 ( .A(n25867), .B(n27448), .Y(n24673) );
  INVX1 U23230 ( .A(reg_file[455]), .Y(n27448) );
  NOR2X1 U23231 ( .A(n25867), .B(n27406), .Y(n24672) );
  INVX1 U23232 ( .A(reg_file[456]), .Y(n27406) );
  NOR2X1 U23233 ( .A(n25867), .B(n27364), .Y(n24671) );
  INVX1 U23234 ( .A(reg_file[457]), .Y(n27364) );
  NOR2X1 U23235 ( .A(n25867), .B(n27322), .Y(n24670) );
  INVX1 U23236 ( .A(reg_file[458]), .Y(n27322) );
  NOR2X1 U23237 ( .A(n25867), .B(n27280), .Y(n24669) );
  INVX1 U23238 ( .A(reg_file[459]), .Y(n27280) );
  NOR2X1 U23239 ( .A(n25867), .B(n27238), .Y(n24668) );
  INVX1 U23240 ( .A(reg_file[460]), .Y(n27238) );
  NOR2X1 U23241 ( .A(n25867), .B(n27196), .Y(n24667) );
  INVX1 U23242 ( .A(reg_file[461]), .Y(n27196) );
  NOR2X1 U23243 ( .A(n25867), .B(n27154), .Y(n24666) );
  INVX1 U23244 ( .A(reg_file[462]), .Y(n27154) );
  NOR2X1 U23245 ( .A(n25867), .B(n27112), .Y(n24665) );
  INVX1 U23246 ( .A(reg_file[463]), .Y(n27112) );
  NOR2X1 U23247 ( .A(n25867), .B(n27028), .Y(n24664) );
  INVX1 U23248 ( .A(reg_file[464]), .Y(n27028) );
  NOR2X1 U23249 ( .A(n25867), .B(n26986), .Y(n24663) );
  INVX1 U23250 ( .A(reg_file[465]), .Y(n26986) );
  NOR2X1 U23251 ( .A(n25868), .B(n26944), .Y(n24662) );
  INVX1 U23252 ( .A(reg_file[466]), .Y(n26944) );
  NOR2X1 U23253 ( .A(n25868), .B(n26902), .Y(n24661) );
  INVX1 U23254 ( .A(reg_file[467]), .Y(n26902) );
  NOR2X1 U23255 ( .A(n25868), .B(n26860), .Y(n24660) );
  INVX1 U23256 ( .A(reg_file[468]), .Y(n26860) );
  NOR2X1 U23257 ( .A(n25868), .B(n26818), .Y(n24659) );
  INVX1 U23258 ( .A(reg_file[469]), .Y(n26818) );
  NOR2X1 U23259 ( .A(n25868), .B(n26776), .Y(n24658) );
  INVX1 U23260 ( .A(reg_file[470]), .Y(n26776) );
  NOR2X1 U23261 ( .A(n25868), .B(n26734), .Y(n24657) );
  INVX1 U23262 ( .A(reg_file[471]), .Y(n26734) );
  NOR2X1 U23263 ( .A(n25868), .B(n26692), .Y(n24656) );
  INVX1 U23264 ( .A(reg_file[472]), .Y(n26692) );
  NOR2X1 U23265 ( .A(n25868), .B(n26650), .Y(n24655) );
  INVX1 U23266 ( .A(reg_file[473]), .Y(n26650) );
  NOR2X1 U23267 ( .A(n25868), .B(n26566), .Y(n24654) );
  INVX1 U23268 ( .A(reg_file[474]), .Y(n26566) );
  NOR2X1 U23269 ( .A(n25868), .B(n26524), .Y(n24653) );
  INVX1 U23270 ( .A(reg_file[475]), .Y(n26524) );
  NOR2X1 U23271 ( .A(n25868), .B(n26482), .Y(n24652) );
  INVX1 U23272 ( .A(reg_file[476]), .Y(n26482) );
  NOR2X1 U23273 ( .A(n25868), .B(n26440), .Y(n24651) );
  INVX1 U23274 ( .A(reg_file[477]), .Y(n26440) );
  NOR2X1 U23275 ( .A(n25868), .B(n26398), .Y(n24650) );
  INVX1 U23276 ( .A(reg_file[478]), .Y(n26398) );
  NOR2X1 U23277 ( .A(n25868), .B(n26356), .Y(n24649) );
  INVX1 U23278 ( .A(reg_file[479]), .Y(n26356) );
  NOR2X1 U23279 ( .A(n25868), .B(n26314), .Y(n24648) );
  INVX1 U23280 ( .A(reg_file[480]), .Y(n26314) );
  NOR2X1 U23281 ( .A(n25868), .B(n26272), .Y(n24647) );
  INVX1 U23282 ( .A(reg_file[481]), .Y(n26272) );
  NOR2X1 U23283 ( .A(n25868), .B(n26230), .Y(n24646) );
  INVX1 U23284 ( .A(reg_file[482]), .Y(n26230) );
  NOR2X1 U23285 ( .A(n25869), .B(n26188), .Y(n24645) );
  INVX1 U23286 ( .A(reg_file[483]), .Y(n26188) );
  NOR2X1 U23287 ( .A(n25869), .B(n31438), .Y(n24644) );
  INVX1 U23288 ( .A(reg_file[484]), .Y(n31438) );
  NOR2X1 U23289 ( .A(n25869), .B(n31396), .Y(n24643) );
  INVX1 U23290 ( .A(reg_file[485]), .Y(n31396) );
  NOR2X1 U23291 ( .A(n25869), .B(n31354), .Y(n24642) );
  INVX1 U23292 ( .A(reg_file[486]), .Y(n31354) );
  NOR2X1 U23293 ( .A(n25869), .B(n31312), .Y(n24641) );
  INVX1 U23294 ( .A(reg_file[487]), .Y(n31312) );
  NOR2X1 U23295 ( .A(n25869), .B(n31270), .Y(n24640) );
  INVX1 U23296 ( .A(reg_file[488]), .Y(n31270) );
  NOR2X1 U23297 ( .A(n25869), .B(n31228), .Y(n24639) );
  INVX1 U23298 ( .A(reg_file[489]), .Y(n31228) );
  NOR2X1 U23299 ( .A(n25869), .B(n31186), .Y(n24638) );
  INVX1 U23300 ( .A(reg_file[490]), .Y(n31186) );
  NOR2X1 U23301 ( .A(n25869), .B(n31144), .Y(n24637) );
  INVX1 U23302 ( .A(reg_file[491]), .Y(n31144) );
  NOR2X1 U23303 ( .A(n25869), .B(n31102), .Y(n24636) );
  INVX1 U23304 ( .A(reg_file[492]), .Y(n31102) );
  NOR2X1 U23305 ( .A(n25869), .B(n31060), .Y(n24635) );
  INVX1 U23306 ( .A(reg_file[493]), .Y(n31060) );
  NOR2X1 U23307 ( .A(n25869), .B(n30976), .Y(n24634) );
  INVX1 U23308 ( .A(reg_file[494]), .Y(n30976) );
  NOR2X1 U23309 ( .A(n25869), .B(n30934), .Y(n24633) );
  INVX1 U23310 ( .A(reg_file[495]), .Y(n30934) );
  NOR2X1 U23311 ( .A(n25869), .B(n30892), .Y(n24632) );
  INVX1 U23312 ( .A(reg_file[496]), .Y(n30892) );
  NOR2X1 U23313 ( .A(n25869), .B(n30850), .Y(n24631) );
  INVX1 U23314 ( .A(reg_file[497]), .Y(n30850) );
  NOR2X1 U23315 ( .A(n25869), .B(n30808), .Y(n24630) );
  INVX1 U23316 ( .A(reg_file[498]), .Y(n30808) );
  NOR2X1 U23317 ( .A(n25869), .B(n30766), .Y(n24629) );
  INVX1 U23318 ( .A(reg_file[499]), .Y(n30766) );
  NOR2X1 U23319 ( .A(n25870), .B(n30724), .Y(n24628) );
  INVX1 U23320 ( .A(reg_file[500]), .Y(n30724) );
  NOR2X1 U23321 ( .A(n25870), .B(n30682), .Y(n24627) );
  INVX1 U23322 ( .A(reg_file[501]), .Y(n30682) );
  NOR2X1 U23323 ( .A(n25870), .B(n30640), .Y(n24626) );
  INVX1 U23324 ( .A(reg_file[502]), .Y(n30640) );
  NOR2X1 U23325 ( .A(n25870), .B(n30598), .Y(n24625) );
  INVX1 U23326 ( .A(reg_file[503]), .Y(n30598) );
  NOR2X1 U23327 ( .A(n25870), .B(n30514), .Y(n24624) );
  INVX1 U23328 ( .A(reg_file[504]), .Y(n30514) );
  NOR2X1 U23329 ( .A(n25870), .B(n30472), .Y(n24623) );
  INVX1 U23330 ( .A(reg_file[505]), .Y(n30472) );
  NOR2X1 U23331 ( .A(n25870), .B(n30430), .Y(n24622) );
  INVX1 U23332 ( .A(reg_file[506]), .Y(n30430) );
  NOR2X1 U23333 ( .A(n25870), .B(n30388), .Y(n24621) );
  INVX1 U23334 ( .A(reg_file[507]), .Y(n30388) );
  NOR2X1 U23335 ( .A(n25870), .B(n30346), .Y(n24620) );
  INVX1 U23336 ( .A(reg_file[508]), .Y(n30346) );
  NOR2X1 U23337 ( .A(n25870), .B(n30304), .Y(n24619) );
  INVX1 U23338 ( .A(reg_file[509]), .Y(n30304) );
  NOR2X1 U23339 ( .A(n25870), .B(n30262), .Y(n24618) );
  INVX1 U23340 ( .A(reg_file[510]), .Y(n30262) );
  NOR2X1 U23341 ( .A(n25870), .B(n30220), .Y(n24617) );
  INVX1 U23342 ( .A(reg_file[511]), .Y(n30220) );
  NOR2X1 U23343 ( .A(n34927), .B(n34925), .Y(n34928) );
  MUX2X1 U23344 ( .B(n34929), .A(n25129), .S(n25871), .Y(n24616) );
  INVX1 U23345 ( .A(reg_file[512]), .Y(n34929) );
  MUX2X1 U23346 ( .B(n34931), .A(n25130), .S(n25871), .Y(n24615) );
  INVX1 U23347 ( .A(reg_file[513]), .Y(n34931) );
  MUX2X1 U23348 ( .B(n34932), .A(n25131), .S(n25871), .Y(n24614) );
  INVX1 U23349 ( .A(reg_file[514]), .Y(n34932) );
  MUX2X1 U23350 ( .B(n34933), .A(n25132), .S(n25871), .Y(n24613) );
  INVX1 U23351 ( .A(reg_file[515]), .Y(n34933) );
  MUX2X1 U23352 ( .B(n34934), .A(n25133), .S(n25871), .Y(n24612) );
  INVX1 U23353 ( .A(reg_file[516]), .Y(n34934) );
  MUX2X1 U23354 ( .B(n34935), .A(n25134), .S(n25871), .Y(n24611) );
  INVX1 U23355 ( .A(reg_file[517]), .Y(n34935) );
  MUX2X1 U23356 ( .B(n34936), .A(n25135), .S(n25871), .Y(n24610) );
  INVX1 U23357 ( .A(reg_file[518]), .Y(n34936) );
  MUX2X1 U23358 ( .B(n34937), .A(n25136), .S(n25871), .Y(n24609) );
  INVX1 U23359 ( .A(reg_file[519]), .Y(n34937) );
  NOR2X1 U23360 ( .A(n25871), .B(n34938), .Y(n24608) );
  INVX1 U23361 ( .A(reg_file[520]), .Y(n34938) );
  NOR2X1 U23362 ( .A(n25871), .B(n34939), .Y(n24607) );
  INVX1 U23363 ( .A(reg_file[521]), .Y(n34939) );
  NOR2X1 U23364 ( .A(n25871), .B(n34940), .Y(n24606) );
  INVX1 U23365 ( .A(reg_file[522]), .Y(n34940) );
  NOR2X1 U23366 ( .A(n25871), .B(n34941), .Y(n24605) );
  INVX1 U23367 ( .A(reg_file[523]), .Y(n34941) );
  NOR2X1 U23368 ( .A(n25871), .B(n34942), .Y(n24604) );
  INVX1 U23369 ( .A(reg_file[524]), .Y(n34942) );
  NOR2X1 U23370 ( .A(n25871), .B(n34943), .Y(n24603) );
  INVX1 U23371 ( .A(reg_file[525]), .Y(n34943) );
  NOR2X1 U23372 ( .A(n25872), .B(n34944), .Y(n24602) );
  INVX1 U23373 ( .A(reg_file[526]), .Y(n34944) );
  NOR2X1 U23374 ( .A(n25872), .B(n34945), .Y(n24601) );
  INVX1 U23375 ( .A(reg_file[527]), .Y(n34945) );
  NOR2X1 U23376 ( .A(n25872), .B(n34946), .Y(n24600) );
  INVX1 U23377 ( .A(reg_file[528]), .Y(n34946) );
  NOR2X1 U23378 ( .A(n25872), .B(n34947), .Y(n24599) );
  INVX1 U23379 ( .A(reg_file[529]), .Y(n34947) );
  NOR2X1 U23380 ( .A(n25872), .B(n34948), .Y(n24598) );
  INVX1 U23381 ( .A(reg_file[530]), .Y(n34948) );
  NOR2X1 U23382 ( .A(n25872), .B(n34949), .Y(n24597) );
  INVX1 U23383 ( .A(reg_file[531]), .Y(n34949) );
  NOR2X1 U23384 ( .A(n25872), .B(n34950), .Y(n24596) );
  INVX1 U23385 ( .A(reg_file[532]), .Y(n34950) );
  NOR2X1 U23386 ( .A(n25872), .B(n34951), .Y(n24595) );
  INVX1 U23387 ( .A(reg_file[533]), .Y(n34951) );
  NOR2X1 U23388 ( .A(n25872), .B(n34952), .Y(n24594) );
  INVX1 U23389 ( .A(reg_file[534]), .Y(n34952) );
  NOR2X1 U23390 ( .A(n25872), .B(n34953), .Y(n24593) );
  INVX1 U23391 ( .A(reg_file[535]), .Y(n34953) );
  NOR2X1 U23392 ( .A(n25872), .B(n34954), .Y(n24592) );
  INVX1 U23393 ( .A(reg_file[536]), .Y(n34954) );
  NOR2X1 U23394 ( .A(n25872), .B(n34955), .Y(n24591) );
  INVX1 U23395 ( .A(reg_file[537]), .Y(n34955) );
  NOR2X1 U23396 ( .A(n25872), .B(n34956), .Y(n24590) );
  INVX1 U23397 ( .A(reg_file[538]), .Y(n34956) );
  NOR2X1 U23398 ( .A(n25872), .B(n34957), .Y(n24589) );
  INVX1 U23399 ( .A(reg_file[539]), .Y(n34957) );
  NOR2X1 U23400 ( .A(n25872), .B(n34958), .Y(n24588) );
  INVX1 U23401 ( .A(reg_file[540]), .Y(n34958) );
  NOR2X1 U23402 ( .A(n25872), .B(n34959), .Y(n24587) );
  INVX1 U23403 ( .A(reg_file[541]), .Y(n34959) );
  NOR2X1 U23404 ( .A(n25872), .B(n34960), .Y(n24586) );
  INVX1 U23405 ( .A(reg_file[542]), .Y(n34960) );
  NOR2X1 U23406 ( .A(n25873), .B(n34961), .Y(n24585) );
  INVX1 U23407 ( .A(reg_file[543]), .Y(n34961) );
  NOR2X1 U23408 ( .A(n25873), .B(n34962), .Y(n24584) );
  INVX1 U23409 ( .A(reg_file[544]), .Y(n34962) );
  NOR2X1 U23410 ( .A(n25873), .B(n34963), .Y(n24583) );
  INVX1 U23411 ( .A(reg_file[545]), .Y(n34963) );
  NOR2X1 U23412 ( .A(n25873), .B(n34964), .Y(n24582) );
  INVX1 U23413 ( .A(reg_file[546]), .Y(n34964) );
  NOR2X1 U23414 ( .A(n25873), .B(n34965), .Y(n24581) );
  INVX1 U23415 ( .A(reg_file[547]), .Y(n34965) );
  NOR2X1 U23416 ( .A(n25873), .B(n34966), .Y(n24580) );
  INVX1 U23417 ( .A(reg_file[548]), .Y(n34966) );
  NOR2X1 U23418 ( .A(n25873), .B(n34967), .Y(n24579) );
  INVX1 U23419 ( .A(reg_file[549]), .Y(n34967) );
  NOR2X1 U23420 ( .A(n25873), .B(n34968), .Y(n24578) );
  INVX1 U23421 ( .A(reg_file[550]), .Y(n34968) );
  NOR2X1 U23422 ( .A(n25873), .B(n34969), .Y(n24577) );
  INVX1 U23423 ( .A(reg_file[551]), .Y(n34969) );
  NOR2X1 U23424 ( .A(n25873), .B(n34970), .Y(n24576) );
  INVX1 U23425 ( .A(reg_file[552]), .Y(n34970) );
  NOR2X1 U23426 ( .A(n25873), .B(n34971), .Y(n24575) );
  INVX1 U23427 ( .A(reg_file[553]), .Y(n34971) );
  NOR2X1 U23428 ( .A(n25873), .B(n34972), .Y(n24574) );
  INVX1 U23429 ( .A(reg_file[554]), .Y(n34972) );
  NOR2X1 U23430 ( .A(n25873), .B(n34973), .Y(n24573) );
  INVX1 U23431 ( .A(reg_file[555]), .Y(n34973) );
  NOR2X1 U23432 ( .A(n25873), .B(n34974), .Y(n24572) );
  INVX1 U23433 ( .A(reg_file[556]), .Y(n34974) );
  NOR2X1 U23434 ( .A(n25873), .B(n34975), .Y(n24571) );
  INVX1 U23435 ( .A(reg_file[557]), .Y(n34975) );
  NOR2X1 U23436 ( .A(n25873), .B(n34976), .Y(n24570) );
  INVX1 U23437 ( .A(reg_file[558]), .Y(n34976) );
  NOR2X1 U23438 ( .A(n25873), .B(n34977), .Y(n24569) );
  INVX1 U23439 ( .A(reg_file[559]), .Y(n34977) );
  NOR2X1 U23440 ( .A(n25874), .B(n34978), .Y(n24568) );
  INVX1 U23441 ( .A(reg_file[560]), .Y(n34978) );
  NOR2X1 U23442 ( .A(n25874), .B(n34979), .Y(n24567) );
  INVX1 U23443 ( .A(reg_file[561]), .Y(n34979) );
  NOR2X1 U23444 ( .A(n25874), .B(n34980), .Y(n24566) );
  INVX1 U23445 ( .A(reg_file[562]), .Y(n34980) );
  NOR2X1 U23446 ( .A(n25874), .B(n34981), .Y(n24565) );
  INVX1 U23447 ( .A(reg_file[563]), .Y(n34981) );
  NOR2X1 U23448 ( .A(n25874), .B(n34982), .Y(n24564) );
  INVX1 U23449 ( .A(reg_file[564]), .Y(n34982) );
  NOR2X1 U23450 ( .A(n25874), .B(n34983), .Y(n24563) );
  INVX1 U23451 ( .A(reg_file[565]), .Y(n34983) );
  NOR2X1 U23452 ( .A(n25874), .B(n34984), .Y(n24562) );
  INVX1 U23453 ( .A(reg_file[566]), .Y(n34984) );
  NOR2X1 U23454 ( .A(n25874), .B(n34985), .Y(n24561) );
  INVX1 U23455 ( .A(reg_file[567]), .Y(n34985) );
  NOR2X1 U23456 ( .A(n25874), .B(n34986), .Y(n24560) );
  INVX1 U23457 ( .A(reg_file[568]), .Y(n34986) );
  NOR2X1 U23458 ( .A(n25874), .B(n34987), .Y(n24559) );
  INVX1 U23459 ( .A(reg_file[569]), .Y(n34987) );
  NOR2X1 U23460 ( .A(n25874), .B(n34988), .Y(n24558) );
  INVX1 U23461 ( .A(reg_file[570]), .Y(n34988) );
  NOR2X1 U23462 ( .A(n25874), .B(n34989), .Y(n24557) );
  INVX1 U23463 ( .A(reg_file[571]), .Y(n34989) );
  NOR2X1 U23464 ( .A(n25874), .B(n34990), .Y(n24556) );
  INVX1 U23465 ( .A(reg_file[572]), .Y(n34990) );
  NOR2X1 U23466 ( .A(n25874), .B(n34991), .Y(n24555) );
  INVX1 U23467 ( .A(reg_file[573]), .Y(n34991) );
  NOR2X1 U23468 ( .A(n25874), .B(n34992), .Y(n24554) );
  INVX1 U23469 ( .A(reg_file[574]), .Y(n34992) );
  NOR2X1 U23470 ( .A(n25874), .B(n34993), .Y(n24553) );
  INVX1 U23471 ( .A(reg_file[575]), .Y(n34993) );
  NOR2X1 U23472 ( .A(n25874), .B(n34994), .Y(n24552) );
  INVX1 U23473 ( .A(reg_file[576]), .Y(n34994) );
  NOR2X1 U23474 ( .A(n25875), .B(n34995), .Y(n24551) );
  INVX1 U23475 ( .A(reg_file[577]), .Y(n34995) );
  NOR2X1 U23476 ( .A(n25875), .B(n34996), .Y(n24550) );
  INVX1 U23477 ( .A(reg_file[578]), .Y(n34996) );
  NOR2X1 U23478 ( .A(n25875), .B(n34997), .Y(n24549) );
  INVX1 U23479 ( .A(reg_file[579]), .Y(n34997) );
  NOR2X1 U23480 ( .A(n25875), .B(n34998), .Y(n24548) );
  INVX1 U23481 ( .A(reg_file[580]), .Y(n34998) );
  NOR2X1 U23482 ( .A(n25875), .B(n34999), .Y(n24547) );
  INVX1 U23483 ( .A(reg_file[581]), .Y(n34999) );
  NOR2X1 U23484 ( .A(n25875), .B(n35000), .Y(n24546) );
  INVX1 U23485 ( .A(reg_file[582]), .Y(n35000) );
  NOR2X1 U23486 ( .A(n25875), .B(n35001), .Y(n24545) );
  INVX1 U23487 ( .A(reg_file[583]), .Y(n35001) );
  NOR2X1 U23488 ( .A(n25875), .B(n35002), .Y(n24544) );
  INVX1 U23489 ( .A(reg_file[584]), .Y(n35002) );
  NOR2X1 U23490 ( .A(n25875), .B(n35003), .Y(n24543) );
  INVX1 U23491 ( .A(reg_file[585]), .Y(n35003) );
  NOR2X1 U23492 ( .A(n25875), .B(n35004), .Y(n24542) );
  INVX1 U23493 ( .A(reg_file[586]), .Y(n35004) );
  NOR2X1 U23494 ( .A(n25875), .B(n35005), .Y(n24541) );
  INVX1 U23495 ( .A(reg_file[587]), .Y(n35005) );
  NOR2X1 U23496 ( .A(n25875), .B(n35006), .Y(n24540) );
  INVX1 U23497 ( .A(reg_file[588]), .Y(n35006) );
  NOR2X1 U23498 ( .A(n25875), .B(n35007), .Y(n24539) );
  INVX1 U23499 ( .A(reg_file[589]), .Y(n35007) );
  NOR2X1 U23500 ( .A(n25875), .B(n35008), .Y(n24538) );
  INVX1 U23501 ( .A(reg_file[590]), .Y(n35008) );
  NOR2X1 U23502 ( .A(n25875), .B(n35009), .Y(n24537) );
  INVX1 U23503 ( .A(reg_file[591]), .Y(n35009) );
  NOR2X1 U23504 ( .A(n25875), .B(n35010), .Y(n24536) );
  INVX1 U23505 ( .A(reg_file[592]), .Y(n35010) );
  NOR2X1 U23506 ( .A(n25875), .B(n35011), .Y(n24535) );
  INVX1 U23507 ( .A(reg_file[593]), .Y(n35011) );
  NOR2X1 U23508 ( .A(n25876), .B(n35012), .Y(n24534) );
  INVX1 U23509 ( .A(reg_file[594]), .Y(n35012) );
  NOR2X1 U23510 ( .A(n25876), .B(n35013), .Y(n24533) );
  INVX1 U23511 ( .A(reg_file[595]), .Y(n35013) );
  NOR2X1 U23512 ( .A(n25876), .B(n35014), .Y(n24532) );
  INVX1 U23513 ( .A(reg_file[596]), .Y(n35014) );
  NOR2X1 U23514 ( .A(n25876), .B(n35015), .Y(n24531) );
  INVX1 U23515 ( .A(reg_file[597]), .Y(n35015) );
  NOR2X1 U23516 ( .A(n25876), .B(n35016), .Y(n24530) );
  INVX1 U23517 ( .A(reg_file[598]), .Y(n35016) );
  NOR2X1 U23518 ( .A(n25876), .B(n35017), .Y(n24529) );
  INVX1 U23519 ( .A(reg_file[599]), .Y(n35017) );
  NOR2X1 U23520 ( .A(n25876), .B(n35018), .Y(n24528) );
  INVX1 U23521 ( .A(reg_file[600]), .Y(n35018) );
  NOR2X1 U23522 ( .A(n25876), .B(n35019), .Y(n24527) );
  INVX1 U23523 ( .A(reg_file[601]), .Y(n35019) );
  NOR2X1 U23524 ( .A(n25876), .B(n35020), .Y(n24526) );
  INVX1 U23525 ( .A(reg_file[602]), .Y(n35020) );
  NOR2X1 U23526 ( .A(n25876), .B(n35021), .Y(n24525) );
  INVX1 U23527 ( .A(reg_file[603]), .Y(n35021) );
  NOR2X1 U23528 ( .A(n25876), .B(n35022), .Y(n24524) );
  INVX1 U23529 ( .A(reg_file[604]), .Y(n35022) );
  NOR2X1 U23530 ( .A(n25876), .B(n35023), .Y(n24523) );
  INVX1 U23531 ( .A(reg_file[605]), .Y(n35023) );
  NOR2X1 U23532 ( .A(n25876), .B(n35024), .Y(n24522) );
  INVX1 U23533 ( .A(reg_file[606]), .Y(n35024) );
  NOR2X1 U23534 ( .A(n25876), .B(n35025), .Y(n24521) );
  INVX1 U23535 ( .A(reg_file[607]), .Y(n35025) );
  NOR2X1 U23536 ( .A(n25876), .B(n35026), .Y(n24520) );
  INVX1 U23537 ( .A(reg_file[608]), .Y(n35026) );
  NOR2X1 U23538 ( .A(n25876), .B(n35027), .Y(n24519) );
  INVX1 U23539 ( .A(reg_file[609]), .Y(n35027) );
  NOR2X1 U23540 ( .A(n25876), .B(n35028), .Y(n24518) );
  INVX1 U23541 ( .A(reg_file[610]), .Y(n35028) );
  NOR2X1 U23542 ( .A(n25877), .B(n35029), .Y(n24517) );
  INVX1 U23543 ( .A(reg_file[611]), .Y(n35029) );
  NOR2X1 U23544 ( .A(n25877), .B(n35030), .Y(n24516) );
  INVX1 U23545 ( .A(reg_file[612]), .Y(n35030) );
  NOR2X1 U23546 ( .A(n25877), .B(n35031), .Y(n24515) );
  INVX1 U23547 ( .A(reg_file[613]), .Y(n35031) );
  NOR2X1 U23548 ( .A(n25877), .B(n35032), .Y(n24514) );
  INVX1 U23549 ( .A(reg_file[614]), .Y(n35032) );
  NOR2X1 U23550 ( .A(n25877), .B(n35033), .Y(n24513) );
  INVX1 U23551 ( .A(reg_file[615]), .Y(n35033) );
  NOR2X1 U23552 ( .A(n25877), .B(n35034), .Y(n24512) );
  INVX1 U23553 ( .A(reg_file[616]), .Y(n35034) );
  NOR2X1 U23554 ( .A(n25877), .B(n35035), .Y(n24511) );
  INVX1 U23555 ( .A(reg_file[617]), .Y(n35035) );
  NOR2X1 U23556 ( .A(n25877), .B(n35036), .Y(n24510) );
  INVX1 U23557 ( .A(reg_file[618]), .Y(n35036) );
  NOR2X1 U23558 ( .A(n25877), .B(n35037), .Y(n24509) );
  INVX1 U23559 ( .A(reg_file[619]), .Y(n35037) );
  NOR2X1 U23560 ( .A(n25877), .B(n35038), .Y(n24508) );
  INVX1 U23561 ( .A(reg_file[620]), .Y(n35038) );
  NOR2X1 U23562 ( .A(n25877), .B(n35039), .Y(n24507) );
  INVX1 U23563 ( .A(reg_file[621]), .Y(n35039) );
  NOR2X1 U23564 ( .A(n25877), .B(n35040), .Y(n24506) );
  INVX1 U23565 ( .A(reg_file[622]), .Y(n35040) );
  NOR2X1 U23566 ( .A(n25877), .B(n35041), .Y(n24505) );
  INVX1 U23567 ( .A(reg_file[623]), .Y(n35041) );
  NOR2X1 U23568 ( .A(n25877), .B(n35042), .Y(n24504) );
  INVX1 U23569 ( .A(reg_file[624]), .Y(n35042) );
  NOR2X1 U23570 ( .A(n25877), .B(n35043), .Y(n24503) );
  INVX1 U23571 ( .A(reg_file[625]), .Y(n35043) );
  NOR2X1 U23572 ( .A(n25877), .B(n35044), .Y(n24502) );
  INVX1 U23573 ( .A(reg_file[626]), .Y(n35044) );
  NOR2X1 U23574 ( .A(n25877), .B(n35045), .Y(n24501) );
  INVX1 U23575 ( .A(reg_file[627]), .Y(n35045) );
  NOR2X1 U23576 ( .A(n25878), .B(n35046), .Y(n24500) );
  INVX1 U23577 ( .A(reg_file[628]), .Y(n35046) );
  NOR2X1 U23578 ( .A(n25878), .B(n35047), .Y(n24499) );
  INVX1 U23579 ( .A(reg_file[629]), .Y(n35047) );
  NOR2X1 U23580 ( .A(n25878), .B(n35048), .Y(n24498) );
  INVX1 U23581 ( .A(reg_file[630]), .Y(n35048) );
  NOR2X1 U23582 ( .A(n25878), .B(n35049), .Y(n24497) );
  INVX1 U23583 ( .A(reg_file[631]), .Y(n35049) );
  NOR2X1 U23584 ( .A(n25878), .B(n35050), .Y(n24496) );
  INVX1 U23585 ( .A(reg_file[632]), .Y(n35050) );
  NOR2X1 U23586 ( .A(n25878), .B(n35051), .Y(n24495) );
  INVX1 U23587 ( .A(reg_file[633]), .Y(n35051) );
  NOR2X1 U23588 ( .A(n25878), .B(n35052), .Y(n24494) );
  INVX1 U23589 ( .A(reg_file[634]), .Y(n35052) );
  NOR2X1 U23590 ( .A(n25878), .B(n35053), .Y(n24493) );
  INVX1 U23591 ( .A(reg_file[635]), .Y(n35053) );
  NOR2X1 U23592 ( .A(n25878), .B(n35054), .Y(n24492) );
  INVX1 U23593 ( .A(reg_file[636]), .Y(n35054) );
  NOR2X1 U23594 ( .A(n25878), .B(n35055), .Y(n24491) );
  INVX1 U23595 ( .A(reg_file[637]), .Y(n35055) );
  NOR2X1 U23596 ( .A(n25878), .B(n35056), .Y(n24490) );
  INVX1 U23597 ( .A(reg_file[638]), .Y(n35056) );
  NOR2X1 U23598 ( .A(n25878), .B(n35057), .Y(n24489) );
  INVX1 U23599 ( .A(reg_file[639]), .Y(n35057) );
  NOR2X1 U23600 ( .A(n35058), .B(n34922), .Y(n34930) );
  MUX2X1 U23601 ( .B(n35059), .A(n25129), .S(n25879), .Y(n24488) );
  INVX1 U23602 ( .A(reg_file[640]), .Y(n35059) );
  MUX2X1 U23603 ( .B(n35061), .A(n25130), .S(n25879), .Y(n24487) );
  INVX1 U23604 ( .A(reg_file[641]), .Y(n35061) );
  MUX2X1 U23605 ( .B(n35062), .A(n25131), .S(n25879), .Y(n24486) );
  INVX1 U23606 ( .A(reg_file[642]), .Y(n35062) );
  MUX2X1 U23607 ( .B(n35063), .A(n25132), .S(n25879), .Y(n24485) );
  INVX1 U23608 ( .A(reg_file[643]), .Y(n35063) );
  MUX2X1 U23609 ( .B(n35064), .A(n25133), .S(n25879), .Y(n24484) );
  INVX1 U23610 ( .A(reg_file[644]), .Y(n35064) );
  MUX2X1 U23611 ( .B(n35065), .A(n25134), .S(n25879), .Y(n24483) );
  INVX1 U23612 ( .A(reg_file[645]), .Y(n35065) );
  MUX2X1 U23613 ( .B(n35066), .A(n25135), .S(n25879), .Y(n24482) );
  INVX1 U23614 ( .A(reg_file[646]), .Y(n35066) );
  MUX2X1 U23615 ( .B(n35067), .A(n25136), .S(n25879), .Y(n24481) );
  INVX1 U23616 ( .A(reg_file[647]), .Y(n35067) );
  NOR2X1 U23617 ( .A(n25879), .B(n35068), .Y(n24480) );
  INVX1 U23618 ( .A(reg_file[648]), .Y(n35068) );
  NOR2X1 U23619 ( .A(n25879), .B(n35069), .Y(n24479) );
  INVX1 U23620 ( .A(reg_file[649]), .Y(n35069) );
  NOR2X1 U23621 ( .A(n25879), .B(n35070), .Y(n24478) );
  INVX1 U23622 ( .A(reg_file[650]), .Y(n35070) );
  NOR2X1 U23623 ( .A(n25879), .B(n35071), .Y(n24477) );
  INVX1 U23624 ( .A(reg_file[651]), .Y(n35071) );
  NOR2X1 U23625 ( .A(n25879), .B(n35072), .Y(n24476) );
  INVX1 U23626 ( .A(reg_file[652]), .Y(n35072) );
  NOR2X1 U23627 ( .A(n25879), .B(n35073), .Y(n24475) );
  INVX1 U23628 ( .A(reg_file[653]), .Y(n35073) );
  NOR2X1 U23629 ( .A(n25880), .B(n35074), .Y(n24474) );
  INVX1 U23630 ( .A(reg_file[654]), .Y(n35074) );
  NOR2X1 U23631 ( .A(n25880), .B(n35075), .Y(n24473) );
  INVX1 U23632 ( .A(reg_file[655]), .Y(n35075) );
  NOR2X1 U23633 ( .A(n25880), .B(n35076), .Y(n24472) );
  INVX1 U23634 ( .A(reg_file[656]), .Y(n35076) );
  NOR2X1 U23635 ( .A(n25880), .B(n35077), .Y(n24471) );
  INVX1 U23636 ( .A(reg_file[657]), .Y(n35077) );
  NOR2X1 U23637 ( .A(n25880), .B(n35078), .Y(n24470) );
  INVX1 U23638 ( .A(reg_file[658]), .Y(n35078) );
  NOR2X1 U23639 ( .A(n25880), .B(n35079), .Y(n24469) );
  INVX1 U23640 ( .A(reg_file[659]), .Y(n35079) );
  NOR2X1 U23641 ( .A(n25880), .B(n35080), .Y(n24468) );
  INVX1 U23642 ( .A(reg_file[660]), .Y(n35080) );
  NOR2X1 U23643 ( .A(n25880), .B(n35081), .Y(n24467) );
  INVX1 U23644 ( .A(reg_file[661]), .Y(n35081) );
  NOR2X1 U23645 ( .A(n25880), .B(n35082), .Y(n24466) );
  INVX1 U23646 ( .A(reg_file[662]), .Y(n35082) );
  NOR2X1 U23647 ( .A(n25880), .B(n35083), .Y(n24465) );
  INVX1 U23648 ( .A(reg_file[663]), .Y(n35083) );
  NOR2X1 U23649 ( .A(n25880), .B(n35084), .Y(n24464) );
  INVX1 U23650 ( .A(reg_file[664]), .Y(n35084) );
  NOR2X1 U23651 ( .A(n25880), .B(n35085), .Y(n24463) );
  INVX1 U23652 ( .A(reg_file[665]), .Y(n35085) );
  NOR2X1 U23653 ( .A(n25880), .B(n35086), .Y(n24462) );
  INVX1 U23654 ( .A(reg_file[666]), .Y(n35086) );
  NOR2X1 U23655 ( .A(n25880), .B(n35087), .Y(n24461) );
  INVX1 U23656 ( .A(reg_file[667]), .Y(n35087) );
  NOR2X1 U23657 ( .A(n25880), .B(n35088), .Y(n24460) );
  INVX1 U23658 ( .A(reg_file[668]), .Y(n35088) );
  NOR2X1 U23659 ( .A(n25880), .B(n35089), .Y(n24459) );
  INVX1 U23660 ( .A(reg_file[669]), .Y(n35089) );
  NOR2X1 U23661 ( .A(n25880), .B(n35090), .Y(n24458) );
  INVX1 U23662 ( .A(reg_file[670]), .Y(n35090) );
  NOR2X1 U23663 ( .A(n25881), .B(n35091), .Y(n24457) );
  INVX1 U23664 ( .A(reg_file[671]), .Y(n35091) );
  NOR2X1 U23665 ( .A(n25881), .B(n35092), .Y(n24456) );
  INVX1 U23666 ( .A(reg_file[672]), .Y(n35092) );
  NOR2X1 U23667 ( .A(n25881), .B(n35093), .Y(n24455) );
  INVX1 U23668 ( .A(reg_file[673]), .Y(n35093) );
  NOR2X1 U23669 ( .A(n25881), .B(n35094), .Y(n24454) );
  INVX1 U23670 ( .A(reg_file[674]), .Y(n35094) );
  NOR2X1 U23671 ( .A(n25881), .B(n35095), .Y(n24453) );
  INVX1 U23672 ( .A(reg_file[675]), .Y(n35095) );
  NOR2X1 U23673 ( .A(n25881), .B(n35096), .Y(n24452) );
  INVX1 U23674 ( .A(reg_file[676]), .Y(n35096) );
  NOR2X1 U23675 ( .A(n25881), .B(n35097), .Y(n24451) );
  INVX1 U23676 ( .A(reg_file[677]), .Y(n35097) );
  NOR2X1 U23677 ( .A(n25881), .B(n35098), .Y(n24450) );
  INVX1 U23678 ( .A(reg_file[678]), .Y(n35098) );
  NOR2X1 U23679 ( .A(n25881), .B(n35099), .Y(n24449) );
  INVX1 U23680 ( .A(reg_file[679]), .Y(n35099) );
  NOR2X1 U23681 ( .A(n25881), .B(n35100), .Y(n24448) );
  INVX1 U23682 ( .A(reg_file[680]), .Y(n35100) );
  NOR2X1 U23683 ( .A(n25881), .B(n35101), .Y(n24447) );
  INVX1 U23684 ( .A(reg_file[681]), .Y(n35101) );
  NOR2X1 U23685 ( .A(n25881), .B(n35102), .Y(n24446) );
  INVX1 U23686 ( .A(reg_file[682]), .Y(n35102) );
  NOR2X1 U23687 ( .A(n25881), .B(n35103), .Y(n24445) );
  INVX1 U23688 ( .A(reg_file[683]), .Y(n35103) );
  NOR2X1 U23689 ( .A(n25881), .B(n35104), .Y(n24444) );
  INVX1 U23690 ( .A(reg_file[684]), .Y(n35104) );
  NOR2X1 U23691 ( .A(n25881), .B(n35105), .Y(n24443) );
  INVX1 U23692 ( .A(reg_file[685]), .Y(n35105) );
  NOR2X1 U23693 ( .A(n25881), .B(n35106), .Y(n24442) );
  INVX1 U23694 ( .A(reg_file[686]), .Y(n35106) );
  NOR2X1 U23695 ( .A(n25881), .B(n35107), .Y(n24441) );
  INVX1 U23696 ( .A(reg_file[687]), .Y(n35107) );
  NOR2X1 U23697 ( .A(n25882), .B(n35108), .Y(n24440) );
  INVX1 U23698 ( .A(reg_file[688]), .Y(n35108) );
  NOR2X1 U23699 ( .A(n25882), .B(n35109), .Y(n24439) );
  INVX1 U23700 ( .A(reg_file[689]), .Y(n35109) );
  NOR2X1 U23701 ( .A(n25882), .B(n35110), .Y(n24438) );
  INVX1 U23702 ( .A(reg_file[690]), .Y(n35110) );
  NOR2X1 U23703 ( .A(n25882), .B(n35111), .Y(n24437) );
  INVX1 U23704 ( .A(reg_file[691]), .Y(n35111) );
  NOR2X1 U23705 ( .A(n25882), .B(n35112), .Y(n24436) );
  INVX1 U23706 ( .A(reg_file[692]), .Y(n35112) );
  NOR2X1 U23707 ( .A(n25882), .B(n35113), .Y(n24435) );
  INVX1 U23708 ( .A(reg_file[693]), .Y(n35113) );
  NOR2X1 U23709 ( .A(n25882), .B(n35114), .Y(n24434) );
  INVX1 U23710 ( .A(reg_file[694]), .Y(n35114) );
  NOR2X1 U23711 ( .A(n25882), .B(n35115), .Y(n24433) );
  INVX1 U23712 ( .A(reg_file[695]), .Y(n35115) );
  NOR2X1 U23713 ( .A(n25882), .B(n35116), .Y(n24432) );
  INVX1 U23714 ( .A(reg_file[696]), .Y(n35116) );
  NOR2X1 U23715 ( .A(n25882), .B(n35117), .Y(n24431) );
  INVX1 U23716 ( .A(reg_file[697]), .Y(n35117) );
  NOR2X1 U23717 ( .A(n25882), .B(n35118), .Y(n24430) );
  INVX1 U23718 ( .A(reg_file[698]), .Y(n35118) );
  NOR2X1 U23719 ( .A(n25882), .B(n35119), .Y(n24429) );
  INVX1 U23720 ( .A(reg_file[699]), .Y(n35119) );
  NOR2X1 U23721 ( .A(n25882), .B(n35120), .Y(n24428) );
  INVX1 U23722 ( .A(reg_file[700]), .Y(n35120) );
  NOR2X1 U23723 ( .A(n25882), .B(n35121), .Y(n24427) );
  INVX1 U23724 ( .A(reg_file[701]), .Y(n35121) );
  NOR2X1 U23725 ( .A(n25882), .B(n35122), .Y(n24426) );
  INVX1 U23726 ( .A(reg_file[702]), .Y(n35122) );
  NOR2X1 U23727 ( .A(n25882), .B(n35123), .Y(n24425) );
  INVX1 U23728 ( .A(reg_file[703]), .Y(n35123) );
  NOR2X1 U23729 ( .A(n25882), .B(n35124), .Y(n24424) );
  INVX1 U23730 ( .A(reg_file[704]), .Y(n35124) );
  NOR2X1 U23731 ( .A(n25883), .B(n35125), .Y(n24423) );
  INVX1 U23732 ( .A(reg_file[705]), .Y(n35125) );
  NOR2X1 U23733 ( .A(n25883), .B(n35126), .Y(n24422) );
  INVX1 U23734 ( .A(reg_file[706]), .Y(n35126) );
  NOR2X1 U23735 ( .A(n25883), .B(n35127), .Y(n24421) );
  INVX1 U23736 ( .A(reg_file[707]), .Y(n35127) );
  NOR2X1 U23737 ( .A(n25883), .B(n35128), .Y(n24420) );
  INVX1 U23738 ( .A(reg_file[708]), .Y(n35128) );
  NOR2X1 U23739 ( .A(n25883), .B(n35129), .Y(n24419) );
  INVX1 U23740 ( .A(reg_file[709]), .Y(n35129) );
  NOR2X1 U23741 ( .A(n25883), .B(n35130), .Y(n24418) );
  INVX1 U23742 ( .A(reg_file[710]), .Y(n35130) );
  NOR2X1 U23743 ( .A(n25883), .B(n35131), .Y(n24417) );
  INVX1 U23744 ( .A(reg_file[711]), .Y(n35131) );
  NOR2X1 U23745 ( .A(n25883), .B(n35132), .Y(n24416) );
  INVX1 U23746 ( .A(reg_file[712]), .Y(n35132) );
  NOR2X1 U23747 ( .A(n25883), .B(n35133), .Y(n24415) );
  INVX1 U23748 ( .A(reg_file[713]), .Y(n35133) );
  NOR2X1 U23749 ( .A(n25883), .B(n35134), .Y(n24414) );
  INVX1 U23750 ( .A(reg_file[714]), .Y(n35134) );
  NOR2X1 U23751 ( .A(n25883), .B(n35135), .Y(n24413) );
  INVX1 U23752 ( .A(reg_file[715]), .Y(n35135) );
  NOR2X1 U23753 ( .A(n25883), .B(n35136), .Y(n24412) );
  INVX1 U23754 ( .A(reg_file[716]), .Y(n35136) );
  NOR2X1 U23755 ( .A(n25883), .B(n35137), .Y(n24411) );
  INVX1 U23756 ( .A(reg_file[717]), .Y(n35137) );
  NOR2X1 U23757 ( .A(n25883), .B(n35138), .Y(n24410) );
  INVX1 U23758 ( .A(reg_file[718]), .Y(n35138) );
  NOR2X1 U23759 ( .A(n25883), .B(n35139), .Y(n24409) );
  INVX1 U23760 ( .A(reg_file[719]), .Y(n35139) );
  NOR2X1 U23761 ( .A(n25883), .B(n35140), .Y(n24408) );
  INVX1 U23762 ( .A(reg_file[720]), .Y(n35140) );
  NOR2X1 U23763 ( .A(n25883), .B(n35141), .Y(n24407) );
  INVX1 U23764 ( .A(reg_file[721]), .Y(n35141) );
  NOR2X1 U23765 ( .A(n25884), .B(n35142), .Y(n24406) );
  INVX1 U23766 ( .A(reg_file[722]), .Y(n35142) );
  NOR2X1 U23767 ( .A(n25884), .B(n35143), .Y(n24405) );
  INVX1 U23768 ( .A(reg_file[723]), .Y(n35143) );
  NOR2X1 U23769 ( .A(n25884), .B(n35144), .Y(n24404) );
  INVX1 U23770 ( .A(reg_file[724]), .Y(n35144) );
  NOR2X1 U23771 ( .A(n25884), .B(n35145), .Y(n24403) );
  INVX1 U23772 ( .A(reg_file[725]), .Y(n35145) );
  NOR2X1 U23773 ( .A(n25884), .B(n35146), .Y(n24402) );
  INVX1 U23774 ( .A(reg_file[726]), .Y(n35146) );
  NOR2X1 U23775 ( .A(n25884), .B(n35147), .Y(n24401) );
  INVX1 U23776 ( .A(reg_file[727]), .Y(n35147) );
  NOR2X1 U23777 ( .A(n25884), .B(n35148), .Y(n24400) );
  INVX1 U23778 ( .A(reg_file[728]), .Y(n35148) );
  NOR2X1 U23779 ( .A(n25884), .B(n35149), .Y(n24399) );
  INVX1 U23780 ( .A(reg_file[729]), .Y(n35149) );
  NOR2X1 U23781 ( .A(n25884), .B(n35150), .Y(n24398) );
  INVX1 U23782 ( .A(reg_file[730]), .Y(n35150) );
  NOR2X1 U23783 ( .A(n25884), .B(n35151), .Y(n24397) );
  INVX1 U23784 ( .A(reg_file[731]), .Y(n35151) );
  NOR2X1 U23785 ( .A(n25884), .B(n35152), .Y(n24396) );
  INVX1 U23786 ( .A(reg_file[732]), .Y(n35152) );
  NOR2X1 U23787 ( .A(n25884), .B(n35153), .Y(n24395) );
  INVX1 U23788 ( .A(reg_file[733]), .Y(n35153) );
  NOR2X1 U23789 ( .A(n25884), .B(n35154), .Y(n24394) );
  INVX1 U23790 ( .A(reg_file[734]), .Y(n35154) );
  NOR2X1 U23791 ( .A(n25884), .B(n35155), .Y(n24393) );
  INVX1 U23792 ( .A(reg_file[735]), .Y(n35155) );
  NOR2X1 U23793 ( .A(n25884), .B(n35156), .Y(n24392) );
  INVX1 U23794 ( .A(reg_file[736]), .Y(n35156) );
  NOR2X1 U23795 ( .A(n25884), .B(n35157), .Y(n24391) );
  INVX1 U23796 ( .A(reg_file[737]), .Y(n35157) );
  NOR2X1 U23797 ( .A(n25884), .B(n35158), .Y(n24390) );
  INVX1 U23798 ( .A(reg_file[738]), .Y(n35158) );
  NOR2X1 U23799 ( .A(n25885), .B(n35159), .Y(n24389) );
  INVX1 U23800 ( .A(reg_file[739]), .Y(n35159) );
  NOR2X1 U23801 ( .A(n25885), .B(n35160), .Y(n24388) );
  INVX1 U23802 ( .A(reg_file[740]), .Y(n35160) );
  NOR2X1 U23803 ( .A(n25885), .B(n35161), .Y(n24387) );
  INVX1 U23804 ( .A(reg_file[741]), .Y(n35161) );
  NOR2X1 U23805 ( .A(n25885), .B(n35162), .Y(n24386) );
  INVX1 U23806 ( .A(reg_file[742]), .Y(n35162) );
  NOR2X1 U23807 ( .A(n25885), .B(n35163), .Y(n24385) );
  INVX1 U23808 ( .A(reg_file[743]), .Y(n35163) );
  NOR2X1 U23809 ( .A(n25885), .B(n35164), .Y(n24384) );
  INVX1 U23810 ( .A(reg_file[744]), .Y(n35164) );
  NOR2X1 U23811 ( .A(n25885), .B(n35165), .Y(n24383) );
  INVX1 U23812 ( .A(reg_file[745]), .Y(n35165) );
  NOR2X1 U23813 ( .A(n25885), .B(n35166), .Y(n24382) );
  INVX1 U23814 ( .A(reg_file[746]), .Y(n35166) );
  NOR2X1 U23815 ( .A(n25885), .B(n35167), .Y(n24381) );
  INVX1 U23816 ( .A(reg_file[747]), .Y(n35167) );
  NOR2X1 U23817 ( .A(n25885), .B(n35168), .Y(n24380) );
  INVX1 U23818 ( .A(reg_file[748]), .Y(n35168) );
  NOR2X1 U23819 ( .A(n25885), .B(n35169), .Y(n24379) );
  INVX1 U23820 ( .A(reg_file[749]), .Y(n35169) );
  NOR2X1 U23821 ( .A(n25885), .B(n35170), .Y(n24378) );
  INVX1 U23822 ( .A(reg_file[750]), .Y(n35170) );
  NOR2X1 U23823 ( .A(n25885), .B(n35171), .Y(n24377) );
  INVX1 U23824 ( .A(reg_file[751]), .Y(n35171) );
  NOR2X1 U23825 ( .A(n25885), .B(n35172), .Y(n24376) );
  INVX1 U23826 ( .A(reg_file[752]), .Y(n35172) );
  NOR2X1 U23827 ( .A(n25885), .B(n35173), .Y(n24375) );
  INVX1 U23828 ( .A(reg_file[753]), .Y(n35173) );
  NOR2X1 U23829 ( .A(n25885), .B(n35174), .Y(n24374) );
  INVX1 U23830 ( .A(reg_file[754]), .Y(n35174) );
  NOR2X1 U23831 ( .A(n25885), .B(n35175), .Y(n24373) );
  INVX1 U23832 ( .A(reg_file[755]), .Y(n35175) );
  NOR2X1 U23833 ( .A(n25886), .B(n35176), .Y(n24372) );
  INVX1 U23834 ( .A(reg_file[756]), .Y(n35176) );
  NOR2X1 U23835 ( .A(n25886), .B(n35177), .Y(n24371) );
  INVX1 U23836 ( .A(reg_file[757]), .Y(n35177) );
  NOR2X1 U23837 ( .A(n25886), .B(n35178), .Y(n24370) );
  INVX1 U23838 ( .A(reg_file[758]), .Y(n35178) );
  NOR2X1 U23839 ( .A(n25886), .B(n35179), .Y(n24369) );
  INVX1 U23840 ( .A(reg_file[759]), .Y(n35179) );
  NOR2X1 U23841 ( .A(n25886), .B(n35180), .Y(n24368) );
  INVX1 U23842 ( .A(reg_file[760]), .Y(n35180) );
  NOR2X1 U23843 ( .A(n25886), .B(n35181), .Y(n24367) );
  INVX1 U23844 ( .A(reg_file[761]), .Y(n35181) );
  NOR2X1 U23845 ( .A(n25886), .B(n35182), .Y(n24366) );
  INVX1 U23846 ( .A(reg_file[762]), .Y(n35182) );
  NOR2X1 U23847 ( .A(n25886), .B(n35183), .Y(n24365) );
  INVX1 U23848 ( .A(reg_file[763]), .Y(n35183) );
  NOR2X1 U23849 ( .A(n25886), .B(n35184), .Y(n24364) );
  INVX1 U23850 ( .A(reg_file[764]), .Y(n35184) );
  NOR2X1 U23851 ( .A(n25886), .B(n35185), .Y(n24363) );
  INVX1 U23852 ( .A(reg_file[765]), .Y(n35185) );
  NOR2X1 U23853 ( .A(n25886), .B(n35186), .Y(n24362) );
  INVX1 U23854 ( .A(reg_file[766]), .Y(n35186) );
  NOR2X1 U23855 ( .A(n25886), .B(n35187), .Y(n24361) );
  INVX1 U23856 ( .A(reg_file[767]), .Y(n35187) );
  NOR2X1 U23857 ( .A(n35058), .B(n34925), .Y(n35060) );
  MUX2X1 U23858 ( .B(n35188), .A(n25129), .S(n25887), .Y(n24360) );
  INVX1 U23859 ( .A(reg_file[768]), .Y(n35188) );
  MUX2X1 U23860 ( .B(n35190), .A(n25130), .S(n25887), .Y(n24359) );
  INVX1 U23861 ( .A(reg_file[769]), .Y(n35190) );
  MUX2X1 U23862 ( .B(n35191), .A(n25131), .S(n25887), .Y(n24358) );
  INVX1 U23863 ( .A(reg_file[770]), .Y(n35191) );
  MUX2X1 U23864 ( .B(n35192), .A(n25132), .S(n25887), .Y(n24357) );
  INVX1 U23865 ( .A(reg_file[771]), .Y(n35192) );
  MUX2X1 U23866 ( .B(n35193), .A(n25133), .S(n25887), .Y(n24356) );
  INVX1 U23867 ( .A(reg_file[772]), .Y(n35193) );
  MUX2X1 U23868 ( .B(n35194), .A(n25134), .S(n25887), .Y(n24355) );
  INVX1 U23869 ( .A(reg_file[773]), .Y(n35194) );
  MUX2X1 U23870 ( .B(n35195), .A(n25135), .S(n25887), .Y(n24354) );
  INVX1 U23871 ( .A(reg_file[774]), .Y(n35195) );
  MUX2X1 U23872 ( .B(n35196), .A(n25136), .S(n25887), .Y(n24353) );
  INVX1 U23873 ( .A(reg_file[775]), .Y(n35196) );
  NOR2X1 U23874 ( .A(n25887), .B(n35197), .Y(n24352) );
  INVX1 U23875 ( .A(reg_file[776]), .Y(n35197) );
  NOR2X1 U23876 ( .A(n25887), .B(n35198), .Y(n24351) );
  INVX1 U23877 ( .A(reg_file[777]), .Y(n35198) );
  NOR2X1 U23878 ( .A(n25887), .B(n35199), .Y(n24350) );
  INVX1 U23879 ( .A(reg_file[778]), .Y(n35199) );
  NOR2X1 U23880 ( .A(n25887), .B(n35200), .Y(n24349) );
  INVX1 U23881 ( .A(reg_file[779]), .Y(n35200) );
  NOR2X1 U23882 ( .A(n25887), .B(n35201), .Y(n24348) );
  INVX1 U23883 ( .A(reg_file[780]), .Y(n35201) );
  NOR2X1 U23884 ( .A(n25887), .B(n35202), .Y(n24347) );
  INVX1 U23885 ( .A(reg_file[781]), .Y(n35202) );
  NOR2X1 U23886 ( .A(n25888), .B(n35203), .Y(n24346) );
  INVX1 U23887 ( .A(reg_file[782]), .Y(n35203) );
  NOR2X1 U23888 ( .A(n25888), .B(n35204), .Y(n24345) );
  INVX1 U23889 ( .A(reg_file[783]), .Y(n35204) );
  NOR2X1 U23890 ( .A(n25888), .B(n35205), .Y(n24344) );
  INVX1 U23891 ( .A(reg_file[784]), .Y(n35205) );
  NOR2X1 U23892 ( .A(n25888), .B(n35206), .Y(n24343) );
  INVX1 U23893 ( .A(reg_file[785]), .Y(n35206) );
  NOR2X1 U23894 ( .A(n25888), .B(n35207), .Y(n24342) );
  INVX1 U23895 ( .A(reg_file[786]), .Y(n35207) );
  NOR2X1 U23896 ( .A(n25888), .B(n35208), .Y(n24341) );
  INVX1 U23897 ( .A(reg_file[787]), .Y(n35208) );
  NOR2X1 U23898 ( .A(n25888), .B(n35209), .Y(n24340) );
  INVX1 U23899 ( .A(reg_file[788]), .Y(n35209) );
  NOR2X1 U23900 ( .A(n25888), .B(n35210), .Y(n24339) );
  INVX1 U23901 ( .A(reg_file[789]), .Y(n35210) );
  NOR2X1 U23902 ( .A(n25888), .B(n35211), .Y(n24338) );
  INVX1 U23903 ( .A(reg_file[790]), .Y(n35211) );
  NOR2X1 U23904 ( .A(n25888), .B(n35212), .Y(n24337) );
  INVX1 U23905 ( .A(reg_file[791]), .Y(n35212) );
  NOR2X1 U23906 ( .A(n25888), .B(n35213), .Y(n24336) );
  INVX1 U23907 ( .A(reg_file[792]), .Y(n35213) );
  NOR2X1 U23908 ( .A(n25888), .B(n35214), .Y(n24335) );
  INVX1 U23909 ( .A(reg_file[793]), .Y(n35214) );
  NOR2X1 U23910 ( .A(n25888), .B(n35215), .Y(n24334) );
  INVX1 U23911 ( .A(reg_file[794]), .Y(n35215) );
  NOR2X1 U23912 ( .A(n25888), .B(n35216), .Y(n24333) );
  INVX1 U23913 ( .A(reg_file[795]), .Y(n35216) );
  NOR2X1 U23914 ( .A(n25888), .B(n35217), .Y(n24332) );
  INVX1 U23915 ( .A(reg_file[796]), .Y(n35217) );
  NOR2X1 U23916 ( .A(n25888), .B(n35218), .Y(n24331) );
  INVX1 U23917 ( .A(reg_file[797]), .Y(n35218) );
  NOR2X1 U23918 ( .A(n25888), .B(n35219), .Y(n24330) );
  INVX1 U23919 ( .A(reg_file[798]), .Y(n35219) );
  NOR2X1 U23920 ( .A(n25889), .B(n35220), .Y(n24329) );
  INVX1 U23921 ( .A(reg_file[799]), .Y(n35220) );
  NOR2X1 U23922 ( .A(n25889), .B(n35221), .Y(n24328) );
  INVX1 U23923 ( .A(reg_file[800]), .Y(n35221) );
  NOR2X1 U23924 ( .A(n25889), .B(n35222), .Y(n24327) );
  INVX1 U23925 ( .A(reg_file[801]), .Y(n35222) );
  NOR2X1 U23926 ( .A(n25889), .B(n35223), .Y(n24326) );
  INVX1 U23927 ( .A(reg_file[802]), .Y(n35223) );
  NOR2X1 U23928 ( .A(n25889), .B(n35224), .Y(n24325) );
  INVX1 U23929 ( .A(reg_file[803]), .Y(n35224) );
  NOR2X1 U23930 ( .A(n25889), .B(n35225), .Y(n24324) );
  INVX1 U23931 ( .A(reg_file[804]), .Y(n35225) );
  NOR2X1 U23932 ( .A(n25889), .B(n35226), .Y(n24323) );
  INVX1 U23933 ( .A(reg_file[805]), .Y(n35226) );
  NOR2X1 U23934 ( .A(n25889), .B(n35227), .Y(n24322) );
  INVX1 U23935 ( .A(reg_file[806]), .Y(n35227) );
  NOR2X1 U23936 ( .A(n25889), .B(n35228), .Y(n24321) );
  INVX1 U23937 ( .A(reg_file[807]), .Y(n35228) );
  NOR2X1 U23938 ( .A(n25889), .B(n35229), .Y(n24320) );
  INVX1 U23939 ( .A(reg_file[808]), .Y(n35229) );
  NOR2X1 U23940 ( .A(n25889), .B(n35230), .Y(n24319) );
  INVX1 U23941 ( .A(reg_file[809]), .Y(n35230) );
  NOR2X1 U23942 ( .A(n25889), .B(n35231), .Y(n24318) );
  INVX1 U23943 ( .A(reg_file[810]), .Y(n35231) );
  NOR2X1 U23944 ( .A(n25889), .B(n35232), .Y(n24317) );
  INVX1 U23945 ( .A(reg_file[811]), .Y(n35232) );
  NOR2X1 U23946 ( .A(n25889), .B(n35233), .Y(n24316) );
  INVX1 U23947 ( .A(reg_file[812]), .Y(n35233) );
  NOR2X1 U23948 ( .A(n25889), .B(n35234), .Y(n24315) );
  INVX1 U23949 ( .A(reg_file[813]), .Y(n35234) );
  NOR2X1 U23950 ( .A(n25889), .B(n35235), .Y(n24314) );
  INVX1 U23951 ( .A(reg_file[814]), .Y(n35235) );
  NOR2X1 U23952 ( .A(n25889), .B(n35236), .Y(n24313) );
  INVX1 U23953 ( .A(reg_file[815]), .Y(n35236) );
  NOR2X1 U23954 ( .A(n25890), .B(n35237), .Y(n24312) );
  INVX1 U23955 ( .A(reg_file[816]), .Y(n35237) );
  NOR2X1 U23956 ( .A(n25890), .B(n35238), .Y(n24311) );
  INVX1 U23957 ( .A(reg_file[817]), .Y(n35238) );
  NOR2X1 U23958 ( .A(n25890), .B(n35239), .Y(n24310) );
  INVX1 U23959 ( .A(reg_file[818]), .Y(n35239) );
  NOR2X1 U23960 ( .A(n25890), .B(n35240), .Y(n24309) );
  INVX1 U23961 ( .A(reg_file[819]), .Y(n35240) );
  NOR2X1 U23962 ( .A(n25890), .B(n35241), .Y(n24308) );
  INVX1 U23963 ( .A(reg_file[820]), .Y(n35241) );
  NOR2X1 U23964 ( .A(n25890), .B(n35242), .Y(n24307) );
  INVX1 U23965 ( .A(reg_file[821]), .Y(n35242) );
  NOR2X1 U23966 ( .A(n25890), .B(n35243), .Y(n24306) );
  INVX1 U23967 ( .A(reg_file[822]), .Y(n35243) );
  NOR2X1 U23968 ( .A(n25890), .B(n35244), .Y(n24305) );
  INVX1 U23969 ( .A(reg_file[823]), .Y(n35244) );
  NOR2X1 U23970 ( .A(n25890), .B(n35245), .Y(n24304) );
  INVX1 U23971 ( .A(reg_file[824]), .Y(n35245) );
  NOR2X1 U23972 ( .A(n25890), .B(n35246), .Y(n24303) );
  INVX1 U23973 ( .A(reg_file[825]), .Y(n35246) );
  NOR2X1 U23974 ( .A(n25890), .B(n35247), .Y(n24302) );
  INVX1 U23975 ( .A(reg_file[826]), .Y(n35247) );
  NOR2X1 U23976 ( .A(n25890), .B(n35248), .Y(n24301) );
  INVX1 U23977 ( .A(reg_file[827]), .Y(n35248) );
  NOR2X1 U23978 ( .A(n25890), .B(n35249), .Y(n24300) );
  INVX1 U23979 ( .A(reg_file[828]), .Y(n35249) );
  NOR2X1 U23980 ( .A(n25890), .B(n35250), .Y(n24299) );
  INVX1 U23981 ( .A(reg_file[829]), .Y(n35250) );
  NOR2X1 U23982 ( .A(n25890), .B(n35251), .Y(n24298) );
  INVX1 U23983 ( .A(reg_file[830]), .Y(n35251) );
  NOR2X1 U23984 ( .A(n25890), .B(n35252), .Y(n24297) );
  INVX1 U23985 ( .A(reg_file[831]), .Y(n35252) );
  NOR2X1 U23986 ( .A(n25890), .B(n35253), .Y(n24296) );
  INVX1 U23987 ( .A(reg_file[832]), .Y(n35253) );
  NOR2X1 U23988 ( .A(n25891), .B(n35254), .Y(n24295) );
  INVX1 U23989 ( .A(reg_file[833]), .Y(n35254) );
  NOR2X1 U23990 ( .A(n25891), .B(n35255), .Y(n24294) );
  INVX1 U23991 ( .A(reg_file[834]), .Y(n35255) );
  NOR2X1 U23992 ( .A(n25891), .B(n35256), .Y(n24293) );
  INVX1 U23993 ( .A(reg_file[835]), .Y(n35256) );
  NOR2X1 U23994 ( .A(n25891), .B(n35257), .Y(n24292) );
  INVX1 U23995 ( .A(reg_file[836]), .Y(n35257) );
  NOR2X1 U23996 ( .A(n25891), .B(n35258), .Y(n24291) );
  INVX1 U23997 ( .A(reg_file[837]), .Y(n35258) );
  NOR2X1 U23998 ( .A(n25891), .B(n35259), .Y(n24290) );
  INVX1 U23999 ( .A(reg_file[838]), .Y(n35259) );
  NOR2X1 U24000 ( .A(n25891), .B(n35260), .Y(n24289) );
  INVX1 U24001 ( .A(reg_file[839]), .Y(n35260) );
  NOR2X1 U24002 ( .A(n25891), .B(n35261), .Y(n24288) );
  INVX1 U24003 ( .A(reg_file[840]), .Y(n35261) );
  NOR2X1 U24004 ( .A(n25891), .B(n35262), .Y(n24287) );
  INVX1 U24005 ( .A(reg_file[841]), .Y(n35262) );
  NOR2X1 U24006 ( .A(n25891), .B(n35263), .Y(n24286) );
  INVX1 U24007 ( .A(reg_file[842]), .Y(n35263) );
  NOR2X1 U24008 ( .A(n25891), .B(n35264), .Y(n24285) );
  INVX1 U24009 ( .A(reg_file[843]), .Y(n35264) );
  NOR2X1 U24010 ( .A(n25891), .B(n35265), .Y(n24284) );
  INVX1 U24011 ( .A(reg_file[844]), .Y(n35265) );
  NOR2X1 U24012 ( .A(n25891), .B(n35266), .Y(n24283) );
  INVX1 U24013 ( .A(reg_file[845]), .Y(n35266) );
  NOR2X1 U24014 ( .A(n25891), .B(n35267), .Y(n24282) );
  INVX1 U24015 ( .A(reg_file[846]), .Y(n35267) );
  NOR2X1 U24016 ( .A(n25891), .B(n35268), .Y(n24281) );
  INVX1 U24017 ( .A(reg_file[847]), .Y(n35268) );
  NOR2X1 U24018 ( .A(n25891), .B(n35269), .Y(n24280) );
  INVX1 U24019 ( .A(reg_file[848]), .Y(n35269) );
  NOR2X1 U24020 ( .A(n25891), .B(n35270), .Y(n24279) );
  INVX1 U24021 ( .A(reg_file[849]), .Y(n35270) );
  NOR2X1 U24022 ( .A(n25892), .B(n35271), .Y(n24278) );
  INVX1 U24023 ( .A(reg_file[850]), .Y(n35271) );
  NOR2X1 U24024 ( .A(n25892), .B(n35272), .Y(n24277) );
  INVX1 U24025 ( .A(reg_file[851]), .Y(n35272) );
  NOR2X1 U24026 ( .A(n25892), .B(n35273), .Y(n24276) );
  INVX1 U24027 ( .A(reg_file[852]), .Y(n35273) );
  NOR2X1 U24028 ( .A(n25892), .B(n35274), .Y(n24275) );
  INVX1 U24029 ( .A(reg_file[853]), .Y(n35274) );
  NOR2X1 U24030 ( .A(n25892), .B(n35275), .Y(n24274) );
  INVX1 U24031 ( .A(reg_file[854]), .Y(n35275) );
  NOR2X1 U24032 ( .A(n25892), .B(n35276), .Y(n24273) );
  INVX1 U24033 ( .A(reg_file[855]), .Y(n35276) );
  NOR2X1 U24034 ( .A(n25892), .B(n35277), .Y(n24272) );
  INVX1 U24035 ( .A(reg_file[856]), .Y(n35277) );
  NOR2X1 U24036 ( .A(n25892), .B(n35278), .Y(n24271) );
  INVX1 U24037 ( .A(reg_file[857]), .Y(n35278) );
  NOR2X1 U24038 ( .A(n25892), .B(n35279), .Y(n24270) );
  INVX1 U24039 ( .A(reg_file[858]), .Y(n35279) );
  NOR2X1 U24040 ( .A(n25892), .B(n35280), .Y(n24269) );
  INVX1 U24041 ( .A(reg_file[859]), .Y(n35280) );
  NOR2X1 U24042 ( .A(n25892), .B(n35281), .Y(n24268) );
  INVX1 U24043 ( .A(reg_file[860]), .Y(n35281) );
  NOR2X1 U24044 ( .A(n25892), .B(n35282), .Y(n24267) );
  INVX1 U24045 ( .A(reg_file[861]), .Y(n35282) );
  NOR2X1 U24046 ( .A(n25892), .B(n35283), .Y(n24266) );
  INVX1 U24047 ( .A(reg_file[862]), .Y(n35283) );
  NOR2X1 U24048 ( .A(n25892), .B(n35284), .Y(n24265) );
  INVX1 U24049 ( .A(reg_file[863]), .Y(n35284) );
  NOR2X1 U24050 ( .A(n25892), .B(n35285), .Y(n24264) );
  INVX1 U24051 ( .A(reg_file[864]), .Y(n35285) );
  NOR2X1 U24052 ( .A(n25892), .B(n35286), .Y(n24263) );
  INVX1 U24053 ( .A(reg_file[865]), .Y(n35286) );
  NOR2X1 U24054 ( .A(n25892), .B(n35287), .Y(n24262) );
  INVX1 U24055 ( .A(reg_file[866]), .Y(n35287) );
  NOR2X1 U24056 ( .A(n25893), .B(n35288), .Y(n24261) );
  INVX1 U24057 ( .A(reg_file[867]), .Y(n35288) );
  NOR2X1 U24058 ( .A(n25893), .B(n35289), .Y(n24260) );
  INVX1 U24059 ( .A(reg_file[868]), .Y(n35289) );
  NOR2X1 U24060 ( .A(n25893), .B(n35290), .Y(n24259) );
  INVX1 U24061 ( .A(reg_file[869]), .Y(n35290) );
  NOR2X1 U24062 ( .A(n25893), .B(n35291), .Y(n24258) );
  INVX1 U24063 ( .A(reg_file[870]), .Y(n35291) );
  NOR2X1 U24064 ( .A(n25893), .B(n35292), .Y(n24257) );
  INVX1 U24065 ( .A(reg_file[871]), .Y(n35292) );
  NOR2X1 U24066 ( .A(n25893), .B(n35293), .Y(n24256) );
  INVX1 U24067 ( .A(reg_file[872]), .Y(n35293) );
  NOR2X1 U24068 ( .A(n25893), .B(n35294), .Y(n24255) );
  INVX1 U24069 ( .A(reg_file[873]), .Y(n35294) );
  NOR2X1 U24070 ( .A(n25893), .B(n35295), .Y(n24254) );
  INVX1 U24071 ( .A(reg_file[874]), .Y(n35295) );
  NOR2X1 U24072 ( .A(n25893), .B(n35296), .Y(n24253) );
  INVX1 U24073 ( .A(reg_file[875]), .Y(n35296) );
  NOR2X1 U24074 ( .A(n25893), .B(n35297), .Y(n24252) );
  INVX1 U24075 ( .A(reg_file[876]), .Y(n35297) );
  NOR2X1 U24076 ( .A(n25893), .B(n35298), .Y(n24251) );
  INVX1 U24077 ( .A(reg_file[877]), .Y(n35298) );
  NOR2X1 U24078 ( .A(n25893), .B(n35299), .Y(n24250) );
  INVX1 U24079 ( .A(reg_file[878]), .Y(n35299) );
  NOR2X1 U24080 ( .A(n25893), .B(n35300), .Y(n24249) );
  INVX1 U24081 ( .A(reg_file[879]), .Y(n35300) );
  NOR2X1 U24082 ( .A(n25893), .B(n35301), .Y(n24248) );
  INVX1 U24083 ( .A(reg_file[880]), .Y(n35301) );
  NOR2X1 U24084 ( .A(n25893), .B(n35302), .Y(n24247) );
  INVX1 U24085 ( .A(reg_file[881]), .Y(n35302) );
  NOR2X1 U24086 ( .A(n25893), .B(n35303), .Y(n24246) );
  INVX1 U24087 ( .A(reg_file[882]), .Y(n35303) );
  NOR2X1 U24088 ( .A(n25893), .B(n35304), .Y(n24245) );
  INVX1 U24089 ( .A(reg_file[883]), .Y(n35304) );
  NOR2X1 U24090 ( .A(n25894), .B(n35305), .Y(n24244) );
  INVX1 U24091 ( .A(reg_file[884]), .Y(n35305) );
  NOR2X1 U24092 ( .A(n25894), .B(n35306), .Y(n24243) );
  INVX1 U24093 ( .A(reg_file[885]), .Y(n35306) );
  NOR2X1 U24094 ( .A(n25894), .B(n35307), .Y(n24242) );
  INVX1 U24095 ( .A(reg_file[886]), .Y(n35307) );
  NOR2X1 U24096 ( .A(n25894), .B(n35308), .Y(n24241) );
  INVX1 U24097 ( .A(reg_file[887]), .Y(n35308) );
  NOR2X1 U24098 ( .A(n25894), .B(n35309), .Y(n24240) );
  INVX1 U24099 ( .A(reg_file[888]), .Y(n35309) );
  NOR2X1 U24100 ( .A(n25894), .B(n35310), .Y(n24239) );
  INVX1 U24101 ( .A(reg_file[889]), .Y(n35310) );
  NOR2X1 U24102 ( .A(n25894), .B(n35311), .Y(n24238) );
  INVX1 U24103 ( .A(reg_file[890]), .Y(n35311) );
  NOR2X1 U24104 ( .A(n25894), .B(n35312), .Y(n24237) );
  INVX1 U24105 ( .A(reg_file[891]), .Y(n35312) );
  NOR2X1 U24106 ( .A(n25894), .B(n35313), .Y(n24236) );
  INVX1 U24107 ( .A(reg_file[892]), .Y(n35313) );
  NOR2X1 U24108 ( .A(n25894), .B(n35314), .Y(n24235) );
  INVX1 U24109 ( .A(reg_file[893]), .Y(n35314) );
  NOR2X1 U24110 ( .A(n25894), .B(n35315), .Y(n24234) );
  INVX1 U24111 ( .A(reg_file[894]), .Y(n35315) );
  NOR2X1 U24112 ( .A(n25894), .B(n35316), .Y(n24233) );
  INVX1 U24113 ( .A(reg_file[895]), .Y(n35316) );
  NOR2X1 U24114 ( .A(n35317), .B(n34922), .Y(n35189) );
  NAND3X1 U24115 ( .A(n35318), .B(n35319), .C(n35320), .Y(n34922) );
  MUX2X1 U24116 ( .B(n35321), .A(n25129), .S(n25895), .Y(n24232) );
  INVX1 U24117 ( .A(reg_file[896]), .Y(n35321) );
  MUX2X1 U24118 ( .B(n35323), .A(n25130), .S(n25895), .Y(n24231) );
  INVX1 U24119 ( .A(reg_file[897]), .Y(n35323) );
  MUX2X1 U24120 ( .B(n35324), .A(n25131), .S(n25895), .Y(n24230) );
  INVX1 U24121 ( .A(reg_file[898]), .Y(n35324) );
  MUX2X1 U24122 ( .B(n35325), .A(n25132), .S(n25895), .Y(n24229) );
  INVX1 U24123 ( .A(reg_file[899]), .Y(n35325) );
  MUX2X1 U24124 ( .B(n35326), .A(n25133), .S(n25895), .Y(n24228) );
  INVX1 U24125 ( .A(reg_file[900]), .Y(n35326) );
  MUX2X1 U24126 ( .B(n35327), .A(n25134), .S(n25895), .Y(n24227) );
  INVX1 U24127 ( .A(reg_file[901]), .Y(n35327) );
  MUX2X1 U24128 ( .B(n35328), .A(n25135), .S(n25895), .Y(n24226) );
  INVX1 U24129 ( .A(reg_file[902]), .Y(n35328) );
  MUX2X1 U24130 ( .B(n35329), .A(n25136), .S(n25895), .Y(n24225) );
  INVX1 U24131 ( .A(reg_file[903]), .Y(n35329) );
  NOR2X1 U24132 ( .A(n25895), .B(n35330), .Y(n24224) );
  INVX1 U24133 ( .A(reg_file[904]), .Y(n35330) );
  NOR2X1 U24134 ( .A(n25895), .B(n35331), .Y(n24223) );
  INVX1 U24135 ( .A(reg_file[905]), .Y(n35331) );
  NOR2X1 U24136 ( .A(n25895), .B(n35332), .Y(n24222) );
  INVX1 U24137 ( .A(reg_file[906]), .Y(n35332) );
  NOR2X1 U24138 ( .A(n25895), .B(n35333), .Y(n24221) );
  INVX1 U24139 ( .A(reg_file[907]), .Y(n35333) );
  NOR2X1 U24140 ( .A(n25895), .B(n35334), .Y(n24220) );
  INVX1 U24141 ( .A(reg_file[908]), .Y(n35334) );
  NOR2X1 U24142 ( .A(n25895), .B(n35335), .Y(n24219) );
  INVX1 U24143 ( .A(reg_file[909]), .Y(n35335) );
  NOR2X1 U24144 ( .A(n25896), .B(n35336), .Y(n24218) );
  INVX1 U24145 ( .A(reg_file[910]), .Y(n35336) );
  NOR2X1 U24146 ( .A(n25896), .B(n35337), .Y(n24217) );
  INVX1 U24147 ( .A(reg_file[911]), .Y(n35337) );
  NOR2X1 U24148 ( .A(n25896), .B(n35338), .Y(n24216) );
  INVX1 U24149 ( .A(reg_file[912]), .Y(n35338) );
  NOR2X1 U24150 ( .A(n25896), .B(n35339), .Y(n24215) );
  INVX1 U24151 ( .A(reg_file[913]), .Y(n35339) );
  NOR2X1 U24152 ( .A(n25896), .B(n35340), .Y(n24214) );
  INVX1 U24153 ( .A(reg_file[914]), .Y(n35340) );
  NOR2X1 U24154 ( .A(n25896), .B(n35341), .Y(n24213) );
  INVX1 U24155 ( .A(reg_file[915]), .Y(n35341) );
  NOR2X1 U24156 ( .A(n25896), .B(n35342), .Y(n24212) );
  INVX1 U24157 ( .A(reg_file[916]), .Y(n35342) );
  NOR2X1 U24158 ( .A(n25896), .B(n35343), .Y(n24211) );
  INVX1 U24159 ( .A(reg_file[917]), .Y(n35343) );
  NOR2X1 U24160 ( .A(n25896), .B(n35344), .Y(n24210) );
  INVX1 U24161 ( .A(reg_file[918]), .Y(n35344) );
  NOR2X1 U24162 ( .A(n25896), .B(n35345), .Y(n24209) );
  INVX1 U24163 ( .A(reg_file[919]), .Y(n35345) );
  NOR2X1 U24164 ( .A(n25896), .B(n35346), .Y(n24208) );
  INVX1 U24165 ( .A(reg_file[920]), .Y(n35346) );
  NOR2X1 U24166 ( .A(n25896), .B(n35347), .Y(n24207) );
  INVX1 U24167 ( .A(reg_file[921]), .Y(n35347) );
  NOR2X1 U24168 ( .A(n25896), .B(n35348), .Y(n24206) );
  INVX1 U24169 ( .A(reg_file[922]), .Y(n35348) );
  NOR2X1 U24170 ( .A(n25896), .B(n35349), .Y(n24205) );
  INVX1 U24171 ( .A(reg_file[923]), .Y(n35349) );
  NOR2X1 U24172 ( .A(n25896), .B(n35350), .Y(n24204) );
  INVX1 U24173 ( .A(reg_file[924]), .Y(n35350) );
  NOR2X1 U24174 ( .A(n25896), .B(n35351), .Y(n24203) );
  INVX1 U24175 ( .A(reg_file[925]), .Y(n35351) );
  NOR2X1 U24176 ( .A(n25896), .B(n35352), .Y(n24202) );
  INVX1 U24177 ( .A(reg_file[926]), .Y(n35352) );
  NOR2X1 U24178 ( .A(n25897), .B(n35353), .Y(n24201) );
  INVX1 U24179 ( .A(reg_file[927]), .Y(n35353) );
  NOR2X1 U24180 ( .A(n25897), .B(n35354), .Y(n24200) );
  INVX1 U24181 ( .A(reg_file[928]), .Y(n35354) );
  NOR2X1 U24182 ( .A(n25897), .B(n35355), .Y(n24199) );
  INVX1 U24183 ( .A(reg_file[929]), .Y(n35355) );
  NOR2X1 U24184 ( .A(n25897), .B(n35356), .Y(n24198) );
  INVX1 U24185 ( .A(reg_file[930]), .Y(n35356) );
  NOR2X1 U24186 ( .A(n25897), .B(n35357), .Y(n24197) );
  INVX1 U24187 ( .A(reg_file[931]), .Y(n35357) );
  NOR2X1 U24188 ( .A(n25897), .B(n35358), .Y(n24196) );
  INVX1 U24189 ( .A(reg_file[932]), .Y(n35358) );
  NOR2X1 U24190 ( .A(n25897), .B(n35359), .Y(n24195) );
  INVX1 U24191 ( .A(reg_file[933]), .Y(n35359) );
  NOR2X1 U24192 ( .A(n25897), .B(n35360), .Y(n24194) );
  INVX1 U24193 ( .A(reg_file[934]), .Y(n35360) );
  NOR2X1 U24194 ( .A(n25897), .B(n35361), .Y(n24193) );
  INVX1 U24195 ( .A(reg_file[935]), .Y(n35361) );
  NOR2X1 U24196 ( .A(n25897), .B(n35362), .Y(n24192) );
  INVX1 U24197 ( .A(reg_file[936]), .Y(n35362) );
  NOR2X1 U24198 ( .A(n25897), .B(n35363), .Y(n24191) );
  INVX1 U24199 ( .A(reg_file[937]), .Y(n35363) );
  NOR2X1 U24200 ( .A(n25897), .B(n35364), .Y(n24190) );
  INVX1 U24201 ( .A(reg_file[938]), .Y(n35364) );
  NOR2X1 U24202 ( .A(n25897), .B(n35365), .Y(n24189) );
  INVX1 U24203 ( .A(reg_file[939]), .Y(n35365) );
  NOR2X1 U24204 ( .A(n25897), .B(n35366), .Y(n24188) );
  INVX1 U24205 ( .A(reg_file[940]), .Y(n35366) );
  NOR2X1 U24206 ( .A(n25897), .B(n35367), .Y(n24187) );
  INVX1 U24207 ( .A(reg_file[941]), .Y(n35367) );
  NOR2X1 U24208 ( .A(n25897), .B(n35368), .Y(n24186) );
  INVX1 U24209 ( .A(reg_file[942]), .Y(n35368) );
  NOR2X1 U24210 ( .A(n25897), .B(n35369), .Y(n24185) );
  INVX1 U24211 ( .A(reg_file[943]), .Y(n35369) );
  NOR2X1 U24212 ( .A(n25898), .B(n35370), .Y(n24184) );
  INVX1 U24213 ( .A(reg_file[944]), .Y(n35370) );
  NOR2X1 U24214 ( .A(n25898), .B(n35371), .Y(n24183) );
  INVX1 U24215 ( .A(reg_file[945]), .Y(n35371) );
  NOR2X1 U24216 ( .A(n25898), .B(n35372), .Y(n24182) );
  INVX1 U24217 ( .A(reg_file[946]), .Y(n35372) );
  NOR2X1 U24218 ( .A(n25898), .B(n35373), .Y(n24181) );
  INVX1 U24219 ( .A(reg_file[947]), .Y(n35373) );
  NOR2X1 U24220 ( .A(n25898), .B(n35374), .Y(n24180) );
  INVX1 U24221 ( .A(reg_file[948]), .Y(n35374) );
  NOR2X1 U24222 ( .A(n25898), .B(n35375), .Y(n24179) );
  INVX1 U24223 ( .A(reg_file[949]), .Y(n35375) );
  NOR2X1 U24224 ( .A(n25898), .B(n35376), .Y(n24178) );
  INVX1 U24225 ( .A(reg_file[950]), .Y(n35376) );
  NOR2X1 U24226 ( .A(n25898), .B(n35377), .Y(n24177) );
  INVX1 U24227 ( .A(reg_file[951]), .Y(n35377) );
  NOR2X1 U24228 ( .A(n25898), .B(n35378), .Y(n24176) );
  INVX1 U24229 ( .A(reg_file[952]), .Y(n35378) );
  NOR2X1 U24230 ( .A(n25898), .B(n35379), .Y(n24175) );
  INVX1 U24231 ( .A(reg_file[953]), .Y(n35379) );
  NOR2X1 U24232 ( .A(n25898), .B(n35380), .Y(n24174) );
  INVX1 U24233 ( .A(reg_file[954]), .Y(n35380) );
  NOR2X1 U24234 ( .A(n25898), .B(n35381), .Y(n24173) );
  INVX1 U24235 ( .A(reg_file[955]), .Y(n35381) );
  NOR2X1 U24236 ( .A(n25898), .B(n35382), .Y(n24172) );
  INVX1 U24237 ( .A(reg_file[956]), .Y(n35382) );
  NOR2X1 U24238 ( .A(n25898), .B(n35383), .Y(n24171) );
  INVX1 U24239 ( .A(reg_file[957]), .Y(n35383) );
  NOR2X1 U24240 ( .A(n25898), .B(n35384), .Y(n24170) );
  INVX1 U24241 ( .A(reg_file[958]), .Y(n35384) );
  NOR2X1 U24242 ( .A(n25898), .B(n35385), .Y(n24169) );
  INVX1 U24243 ( .A(reg_file[959]), .Y(n35385) );
  NOR2X1 U24244 ( .A(n25898), .B(n35386), .Y(n24168) );
  INVX1 U24245 ( .A(reg_file[960]), .Y(n35386) );
  NOR2X1 U24246 ( .A(n25899), .B(n35387), .Y(n24167) );
  INVX1 U24247 ( .A(reg_file[961]), .Y(n35387) );
  NOR2X1 U24248 ( .A(n25899), .B(n35388), .Y(n24166) );
  INVX1 U24249 ( .A(reg_file[962]), .Y(n35388) );
  NOR2X1 U24250 ( .A(n25899), .B(n35389), .Y(n24165) );
  INVX1 U24251 ( .A(reg_file[963]), .Y(n35389) );
  NOR2X1 U24252 ( .A(n25899), .B(n35390), .Y(n24164) );
  INVX1 U24253 ( .A(reg_file[964]), .Y(n35390) );
  NOR2X1 U24254 ( .A(n25899), .B(n35391), .Y(n24163) );
  INVX1 U24255 ( .A(reg_file[965]), .Y(n35391) );
  NOR2X1 U24256 ( .A(n25899), .B(n35392), .Y(n24162) );
  INVX1 U24257 ( .A(reg_file[966]), .Y(n35392) );
  NOR2X1 U24258 ( .A(n25899), .B(n35393), .Y(n24161) );
  INVX1 U24259 ( .A(reg_file[967]), .Y(n35393) );
  NOR2X1 U24260 ( .A(n25899), .B(n35394), .Y(n24160) );
  INVX1 U24261 ( .A(reg_file[968]), .Y(n35394) );
  NOR2X1 U24262 ( .A(n25899), .B(n35395), .Y(n24159) );
  INVX1 U24263 ( .A(reg_file[969]), .Y(n35395) );
  NOR2X1 U24264 ( .A(n25899), .B(n35396), .Y(n24158) );
  INVX1 U24265 ( .A(reg_file[970]), .Y(n35396) );
  NOR2X1 U24266 ( .A(n25899), .B(n35397), .Y(n24157) );
  INVX1 U24267 ( .A(reg_file[971]), .Y(n35397) );
  NOR2X1 U24268 ( .A(n25899), .B(n35398), .Y(n24156) );
  INVX1 U24269 ( .A(reg_file[972]), .Y(n35398) );
  NOR2X1 U24270 ( .A(n25899), .B(n35399), .Y(n24155) );
  INVX1 U24271 ( .A(reg_file[973]), .Y(n35399) );
  NOR2X1 U24272 ( .A(n25899), .B(n35400), .Y(n24154) );
  INVX1 U24273 ( .A(reg_file[974]), .Y(n35400) );
  NOR2X1 U24274 ( .A(n25899), .B(n35401), .Y(n24153) );
  INVX1 U24275 ( .A(reg_file[975]), .Y(n35401) );
  NOR2X1 U24276 ( .A(n25899), .B(n35402), .Y(n24152) );
  INVX1 U24277 ( .A(reg_file[976]), .Y(n35402) );
  NOR2X1 U24278 ( .A(n25899), .B(n35403), .Y(n24151) );
  INVX1 U24279 ( .A(reg_file[977]), .Y(n35403) );
  NOR2X1 U24280 ( .A(n25900), .B(n35404), .Y(n24150) );
  INVX1 U24281 ( .A(reg_file[978]), .Y(n35404) );
  NOR2X1 U24282 ( .A(n25900), .B(n35405), .Y(n24149) );
  INVX1 U24283 ( .A(reg_file[979]), .Y(n35405) );
  NOR2X1 U24284 ( .A(n25900), .B(n35406), .Y(n24148) );
  INVX1 U24285 ( .A(reg_file[980]), .Y(n35406) );
  NOR2X1 U24286 ( .A(n25900), .B(n35407), .Y(n24147) );
  INVX1 U24287 ( .A(reg_file[981]), .Y(n35407) );
  NOR2X1 U24288 ( .A(n25900), .B(n35408), .Y(n24146) );
  INVX1 U24289 ( .A(reg_file[982]), .Y(n35408) );
  NOR2X1 U24290 ( .A(n25900), .B(n35409), .Y(n24145) );
  INVX1 U24291 ( .A(reg_file[983]), .Y(n35409) );
  NOR2X1 U24292 ( .A(n25900), .B(n35410), .Y(n24144) );
  INVX1 U24293 ( .A(reg_file[984]), .Y(n35410) );
  NOR2X1 U24294 ( .A(n25900), .B(n35411), .Y(n24143) );
  INVX1 U24295 ( .A(reg_file[985]), .Y(n35411) );
  NOR2X1 U24296 ( .A(n25900), .B(n35412), .Y(n24142) );
  INVX1 U24297 ( .A(reg_file[986]), .Y(n35412) );
  NOR2X1 U24298 ( .A(n25900), .B(n35413), .Y(n24141) );
  INVX1 U24299 ( .A(reg_file[987]), .Y(n35413) );
  NOR2X1 U24300 ( .A(n25900), .B(n35414), .Y(n24140) );
  INVX1 U24301 ( .A(reg_file[988]), .Y(n35414) );
  NOR2X1 U24302 ( .A(n25900), .B(n35415), .Y(n24139) );
  INVX1 U24303 ( .A(reg_file[989]), .Y(n35415) );
  NOR2X1 U24304 ( .A(n25900), .B(n35416), .Y(n24138) );
  INVX1 U24305 ( .A(reg_file[990]), .Y(n35416) );
  NOR2X1 U24306 ( .A(n25900), .B(n35417), .Y(n24137) );
  INVX1 U24307 ( .A(reg_file[991]), .Y(n35417) );
  NOR2X1 U24308 ( .A(n25900), .B(n35418), .Y(n24136) );
  INVX1 U24309 ( .A(reg_file[992]), .Y(n35418) );
  NOR2X1 U24310 ( .A(n25900), .B(n35419), .Y(n24135) );
  INVX1 U24311 ( .A(reg_file[993]), .Y(n35419) );
  NOR2X1 U24312 ( .A(n25900), .B(n35420), .Y(n24134) );
  INVX1 U24313 ( .A(reg_file[994]), .Y(n35420) );
  NOR2X1 U24314 ( .A(n25901), .B(n35421), .Y(n24133) );
  INVX1 U24315 ( .A(reg_file[995]), .Y(n35421) );
  NOR2X1 U24316 ( .A(n25901), .B(n35422), .Y(n24132) );
  INVX1 U24317 ( .A(reg_file[996]), .Y(n35422) );
  NOR2X1 U24318 ( .A(n25901), .B(n35423), .Y(n24131) );
  INVX1 U24319 ( .A(reg_file[997]), .Y(n35423) );
  NOR2X1 U24320 ( .A(n25901), .B(n35424), .Y(n24130) );
  INVX1 U24321 ( .A(reg_file[998]), .Y(n35424) );
  NOR2X1 U24322 ( .A(n25901), .B(n35425), .Y(n24129) );
  INVX1 U24323 ( .A(reg_file[999]), .Y(n35425) );
  NOR2X1 U24324 ( .A(n25901), .B(n35426), .Y(n24128) );
  INVX1 U24325 ( .A(reg_file[1000]), .Y(n35426) );
  NOR2X1 U24326 ( .A(n25901), .B(n35427), .Y(n24127) );
  INVX1 U24327 ( .A(reg_file[1001]), .Y(n35427) );
  NOR2X1 U24328 ( .A(n25901), .B(n35428), .Y(n24126) );
  INVX1 U24329 ( .A(reg_file[1002]), .Y(n35428) );
  NOR2X1 U24330 ( .A(n25901), .B(n35429), .Y(n24125) );
  INVX1 U24331 ( .A(reg_file[1003]), .Y(n35429) );
  NOR2X1 U24332 ( .A(n25901), .B(n35430), .Y(n24124) );
  INVX1 U24333 ( .A(reg_file[1004]), .Y(n35430) );
  NOR2X1 U24334 ( .A(n25901), .B(n35431), .Y(n24123) );
  INVX1 U24335 ( .A(reg_file[1005]), .Y(n35431) );
  NOR2X1 U24336 ( .A(n25901), .B(n35432), .Y(n24122) );
  INVX1 U24337 ( .A(reg_file[1006]), .Y(n35432) );
  NOR2X1 U24338 ( .A(n25901), .B(n35433), .Y(n24121) );
  INVX1 U24339 ( .A(reg_file[1007]), .Y(n35433) );
  NOR2X1 U24340 ( .A(n25901), .B(n35434), .Y(n24120) );
  INVX1 U24341 ( .A(reg_file[1008]), .Y(n35434) );
  NOR2X1 U24342 ( .A(n25901), .B(n35435), .Y(n24119) );
  INVX1 U24343 ( .A(reg_file[1009]), .Y(n35435) );
  NOR2X1 U24344 ( .A(n25901), .B(n35436), .Y(n24118) );
  INVX1 U24345 ( .A(reg_file[1010]), .Y(n35436) );
  NOR2X1 U24346 ( .A(n25901), .B(n35437), .Y(n24117) );
  INVX1 U24347 ( .A(reg_file[1011]), .Y(n35437) );
  NOR2X1 U24348 ( .A(n25902), .B(n35438), .Y(n24116) );
  INVX1 U24349 ( .A(reg_file[1012]), .Y(n35438) );
  NOR2X1 U24350 ( .A(n25902), .B(n35439), .Y(n24115) );
  INVX1 U24351 ( .A(reg_file[1013]), .Y(n35439) );
  NOR2X1 U24352 ( .A(n25902), .B(n35440), .Y(n24114) );
  INVX1 U24353 ( .A(reg_file[1014]), .Y(n35440) );
  NOR2X1 U24354 ( .A(n25902), .B(n35441), .Y(n24113) );
  INVX1 U24355 ( .A(reg_file[1015]), .Y(n35441) );
  NOR2X1 U24356 ( .A(n25902), .B(n35442), .Y(n24112) );
  INVX1 U24357 ( .A(reg_file[1016]), .Y(n35442) );
  NOR2X1 U24358 ( .A(n25902), .B(n35443), .Y(n24111) );
  INVX1 U24359 ( .A(reg_file[1017]), .Y(n35443) );
  NOR2X1 U24360 ( .A(n25902), .B(n35444), .Y(n24110) );
  INVX1 U24361 ( .A(reg_file[1018]), .Y(n35444) );
  NOR2X1 U24362 ( .A(n25902), .B(n35445), .Y(n24109) );
  INVX1 U24363 ( .A(reg_file[1019]), .Y(n35445) );
  NOR2X1 U24364 ( .A(n25902), .B(n35446), .Y(n24108) );
  INVX1 U24365 ( .A(reg_file[1020]), .Y(n35446) );
  NOR2X1 U24366 ( .A(n25902), .B(n35447), .Y(n24107) );
  INVX1 U24367 ( .A(reg_file[1021]), .Y(n35447) );
  NOR2X1 U24368 ( .A(n25902), .B(n35448), .Y(n24106) );
  INVX1 U24369 ( .A(reg_file[1022]), .Y(n35448) );
  NOR2X1 U24370 ( .A(n25902), .B(n35449), .Y(n24105) );
  INVX1 U24371 ( .A(reg_file[1023]), .Y(n35449) );
  NOR2X1 U24372 ( .A(n35317), .B(n34925), .Y(n35322) );
  NAND3X1 U24373 ( .A(n35318), .B(n35319), .C(wraddr[0]), .Y(n34925) );
  MUX2X1 U24374 ( .B(n35450), .A(n25129), .S(n25903), .Y(n24104) );
  INVX1 U24375 ( .A(reg_file[1024]), .Y(n35450) );
  MUX2X1 U24376 ( .B(n35452), .A(n25130), .S(n25903), .Y(n24103) );
  INVX1 U24377 ( .A(reg_file[1025]), .Y(n35452) );
  MUX2X1 U24378 ( .B(n35453), .A(n25131), .S(n25903), .Y(n24102) );
  INVX1 U24379 ( .A(reg_file[1026]), .Y(n35453) );
  MUX2X1 U24380 ( .B(n35454), .A(n25132), .S(n25903), .Y(n24101) );
  INVX1 U24381 ( .A(reg_file[1027]), .Y(n35454) );
  MUX2X1 U24382 ( .B(n35455), .A(n25133), .S(n25903), .Y(n24100) );
  INVX1 U24383 ( .A(reg_file[1028]), .Y(n35455) );
  MUX2X1 U24384 ( .B(n35456), .A(n25134), .S(n25903), .Y(n24099) );
  INVX1 U24385 ( .A(reg_file[1029]), .Y(n35456) );
  MUX2X1 U24386 ( .B(n35457), .A(n25135), .S(n25903), .Y(n24098) );
  INVX1 U24387 ( .A(reg_file[1030]), .Y(n35457) );
  MUX2X1 U24388 ( .B(n35458), .A(n25136), .S(n25903), .Y(n24097) );
  INVX1 U24389 ( .A(reg_file[1031]), .Y(n35458) );
  NOR2X1 U24390 ( .A(n25903), .B(n35459), .Y(n24096) );
  INVX1 U24391 ( .A(reg_file[1032]), .Y(n35459) );
  NOR2X1 U24392 ( .A(n25903), .B(n35460), .Y(n24095) );
  INVX1 U24393 ( .A(reg_file[1033]), .Y(n35460) );
  NOR2X1 U24394 ( .A(n25903), .B(n35461), .Y(n24094) );
  INVX1 U24395 ( .A(reg_file[1034]), .Y(n35461) );
  NOR2X1 U24396 ( .A(n25903), .B(n35462), .Y(n24093) );
  INVX1 U24397 ( .A(reg_file[1035]), .Y(n35462) );
  NOR2X1 U24398 ( .A(n25903), .B(n35463), .Y(n24092) );
  INVX1 U24399 ( .A(reg_file[1036]), .Y(n35463) );
  NOR2X1 U24400 ( .A(n25903), .B(n35464), .Y(n24091) );
  INVX1 U24401 ( .A(reg_file[1037]), .Y(n35464) );
  NOR2X1 U24402 ( .A(n25904), .B(n35465), .Y(n24090) );
  INVX1 U24403 ( .A(reg_file[1038]), .Y(n35465) );
  NOR2X1 U24404 ( .A(n25904), .B(n35466), .Y(n24089) );
  INVX1 U24405 ( .A(reg_file[1039]), .Y(n35466) );
  NOR2X1 U24406 ( .A(n25904), .B(n35467), .Y(n24088) );
  INVX1 U24407 ( .A(reg_file[1040]), .Y(n35467) );
  NOR2X1 U24408 ( .A(n25904), .B(n35468), .Y(n24087) );
  INVX1 U24409 ( .A(reg_file[1041]), .Y(n35468) );
  NOR2X1 U24410 ( .A(n25904), .B(n35469), .Y(n24086) );
  INVX1 U24411 ( .A(reg_file[1042]), .Y(n35469) );
  NOR2X1 U24412 ( .A(n25904), .B(n35470), .Y(n24085) );
  INVX1 U24413 ( .A(reg_file[1043]), .Y(n35470) );
  NOR2X1 U24414 ( .A(n25904), .B(n35471), .Y(n24084) );
  INVX1 U24415 ( .A(reg_file[1044]), .Y(n35471) );
  NOR2X1 U24416 ( .A(n25904), .B(n35472), .Y(n24083) );
  INVX1 U24417 ( .A(reg_file[1045]), .Y(n35472) );
  NOR2X1 U24418 ( .A(n25904), .B(n35473), .Y(n24082) );
  INVX1 U24419 ( .A(reg_file[1046]), .Y(n35473) );
  NOR2X1 U24420 ( .A(n25904), .B(n35474), .Y(n24081) );
  INVX1 U24421 ( .A(reg_file[1047]), .Y(n35474) );
  NOR2X1 U24422 ( .A(n25904), .B(n35475), .Y(n24080) );
  INVX1 U24423 ( .A(reg_file[1048]), .Y(n35475) );
  NOR2X1 U24424 ( .A(n25904), .B(n35476), .Y(n24079) );
  INVX1 U24425 ( .A(reg_file[1049]), .Y(n35476) );
  NOR2X1 U24426 ( .A(n25904), .B(n35477), .Y(n24078) );
  INVX1 U24427 ( .A(reg_file[1050]), .Y(n35477) );
  NOR2X1 U24428 ( .A(n25904), .B(n35478), .Y(n24077) );
  INVX1 U24429 ( .A(reg_file[1051]), .Y(n35478) );
  NOR2X1 U24430 ( .A(n25904), .B(n35479), .Y(n24076) );
  INVX1 U24431 ( .A(reg_file[1052]), .Y(n35479) );
  NOR2X1 U24432 ( .A(n25904), .B(n35480), .Y(n24075) );
  INVX1 U24433 ( .A(reg_file[1053]), .Y(n35480) );
  NOR2X1 U24434 ( .A(n25904), .B(n35481), .Y(n24074) );
  INVX1 U24435 ( .A(reg_file[1054]), .Y(n35481) );
  NOR2X1 U24436 ( .A(n25905), .B(n35482), .Y(n24073) );
  INVX1 U24437 ( .A(reg_file[1055]), .Y(n35482) );
  NOR2X1 U24438 ( .A(n25905), .B(n35483), .Y(n24072) );
  INVX1 U24439 ( .A(reg_file[1056]), .Y(n35483) );
  NOR2X1 U24440 ( .A(n25905), .B(n35484), .Y(n24071) );
  INVX1 U24441 ( .A(reg_file[1057]), .Y(n35484) );
  NOR2X1 U24442 ( .A(n25905), .B(n35485), .Y(n24070) );
  INVX1 U24443 ( .A(reg_file[1058]), .Y(n35485) );
  NOR2X1 U24444 ( .A(n25905), .B(n35486), .Y(n24069) );
  INVX1 U24445 ( .A(reg_file[1059]), .Y(n35486) );
  NOR2X1 U24446 ( .A(n25905), .B(n35487), .Y(n24068) );
  INVX1 U24447 ( .A(reg_file[1060]), .Y(n35487) );
  NOR2X1 U24448 ( .A(n25905), .B(n35488), .Y(n24067) );
  INVX1 U24449 ( .A(reg_file[1061]), .Y(n35488) );
  NOR2X1 U24450 ( .A(n25905), .B(n35489), .Y(n24066) );
  INVX1 U24451 ( .A(reg_file[1062]), .Y(n35489) );
  NOR2X1 U24452 ( .A(n25905), .B(n35490), .Y(n24065) );
  INVX1 U24453 ( .A(reg_file[1063]), .Y(n35490) );
  NOR2X1 U24454 ( .A(n25905), .B(n35491), .Y(n24064) );
  INVX1 U24455 ( .A(reg_file[1064]), .Y(n35491) );
  NOR2X1 U24456 ( .A(n25905), .B(n35492), .Y(n24063) );
  INVX1 U24457 ( .A(reg_file[1065]), .Y(n35492) );
  NOR2X1 U24458 ( .A(n25905), .B(n35493), .Y(n24062) );
  INVX1 U24459 ( .A(reg_file[1066]), .Y(n35493) );
  NOR2X1 U24460 ( .A(n25905), .B(n35494), .Y(n24061) );
  INVX1 U24461 ( .A(reg_file[1067]), .Y(n35494) );
  NOR2X1 U24462 ( .A(n25905), .B(n35495), .Y(n24060) );
  INVX1 U24463 ( .A(reg_file[1068]), .Y(n35495) );
  NOR2X1 U24464 ( .A(n25905), .B(n35496), .Y(n24059) );
  INVX1 U24465 ( .A(reg_file[1069]), .Y(n35496) );
  NOR2X1 U24466 ( .A(n25905), .B(n35497), .Y(n24058) );
  INVX1 U24467 ( .A(reg_file[1070]), .Y(n35497) );
  NOR2X1 U24468 ( .A(n25905), .B(n35498), .Y(n24057) );
  INVX1 U24469 ( .A(reg_file[1071]), .Y(n35498) );
  NOR2X1 U24470 ( .A(n25906), .B(n35499), .Y(n24056) );
  INVX1 U24471 ( .A(reg_file[1072]), .Y(n35499) );
  NOR2X1 U24472 ( .A(n25906), .B(n35500), .Y(n24055) );
  INVX1 U24473 ( .A(reg_file[1073]), .Y(n35500) );
  NOR2X1 U24474 ( .A(n25906), .B(n35501), .Y(n24054) );
  INVX1 U24475 ( .A(reg_file[1074]), .Y(n35501) );
  NOR2X1 U24476 ( .A(n25906), .B(n35502), .Y(n24053) );
  INVX1 U24477 ( .A(reg_file[1075]), .Y(n35502) );
  NOR2X1 U24478 ( .A(n25906), .B(n35503), .Y(n24052) );
  INVX1 U24479 ( .A(reg_file[1076]), .Y(n35503) );
  NOR2X1 U24480 ( .A(n25906), .B(n35504), .Y(n24051) );
  INVX1 U24481 ( .A(reg_file[1077]), .Y(n35504) );
  NOR2X1 U24482 ( .A(n25906), .B(n35505), .Y(n24050) );
  INVX1 U24483 ( .A(reg_file[1078]), .Y(n35505) );
  NOR2X1 U24484 ( .A(n25906), .B(n35506), .Y(n24049) );
  INVX1 U24485 ( .A(reg_file[1079]), .Y(n35506) );
  NOR2X1 U24486 ( .A(n25906), .B(n35507), .Y(n24048) );
  INVX1 U24487 ( .A(reg_file[1080]), .Y(n35507) );
  NOR2X1 U24488 ( .A(n25906), .B(n35508), .Y(n24047) );
  INVX1 U24489 ( .A(reg_file[1081]), .Y(n35508) );
  NOR2X1 U24490 ( .A(n25906), .B(n35509), .Y(n24046) );
  INVX1 U24491 ( .A(reg_file[1082]), .Y(n35509) );
  NOR2X1 U24492 ( .A(n25906), .B(n35510), .Y(n24045) );
  INVX1 U24493 ( .A(reg_file[1083]), .Y(n35510) );
  NOR2X1 U24494 ( .A(n25906), .B(n35511), .Y(n24044) );
  INVX1 U24495 ( .A(reg_file[1084]), .Y(n35511) );
  NOR2X1 U24496 ( .A(n25906), .B(n35512), .Y(n24043) );
  INVX1 U24497 ( .A(reg_file[1085]), .Y(n35512) );
  NOR2X1 U24498 ( .A(n25906), .B(n35513), .Y(n24042) );
  INVX1 U24499 ( .A(reg_file[1086]), .Y(n35513) );
  NOR2X1 U24500 ( .A(n25906), .B(n35514), .Y(n24041) );
  INVX1 U24501 ( .A(reg_file[1087]), .Y(n35514) );
  NOR2X1 U24502 ( .A(n25906), .B(n35515), .Y(n24040) );
  INVX1 U24503 ( .A(reg_file[1088]), .Y(n35515) );
  NOR2X1 U24504 ( .A(n25907), .B(n35516), .Y(n24039) );
  INVX1 U24505 ( .A(reg_file[1089]), .Y(n35516) );
  NOR2X1 U24506 ( .A(n25907), .B(n35517), .Y(n24038) );
  INVX1 U24507 ( .A(reg_file[1090]), .Y(n35517) );
  NOR2X1 U24508 ( .A(n25907), .B(n35518), .Y(n24037) );
  INVX1 U24509 ( .A(reg_file[1091]), .Y(n35518) );
  NOR2X1 U24510 ( .A(n25907), .B(n35519), .Y(n24036) );
  INVX1 U24511 ( .A(reg_file[1092]), .Y(n35519) );
  NOR2X1 U24512 ( .A(n25907), .B(n35520), .Y(n24035) );
  INVX1 U24513 ( .A(reg_file[1093]), .Y(n35520) );
  NOR2X1 U24514 ( .A(n25907), .B(n35521), .Y(n24034) );
  INVX1 U24515 ( .A(reg_file[1094]), .Y(n35521) );
  NOR2X1 U24516 ( .A(n25907), .B(n35522), .Y(n24033) );
  INVX1 U24517 ( .A(reg_file[1095]), .Y(n35522) );
  NOR2X1 U24518 ( .A(n25907), .B(n35523), .Y(n24032) );
  INVX1 U24519 ( .A(reg_file[1096]), .Y(n35523) );
  NOR2X1 U24520 ( .A(n25907), .B(n35524), .Y(n24031) );
  INVX1 U24521 ( .A(reg_file[1097]), .Y(n35524) );
  NOR2X1 U24522 ( .A(n25907), .B(n35525), .Y(n24030) );
  INVX1 U24523 ( .A(reg_file[1098]), .Y(n35525) );
  NOR2X1 U24524 ( .A(n25907), .B(n35526), .Y(n24029) );
  INVX1 U24525 ( .A(reg_file[1099]), .Y(n35526) );
  NOR2X1 U24526 ( .A(n25907), .B(n35527), .Y(n24028) );
  INVX1 U24527 ( .A(reg_file[1100]), .Y(n35527) );
  NOR2X1 U24528 ( .A(n25907), .B(n35528), .Y(n24027) );
  INVX1 U24529 ( .A(reg_file[1101]), .Y(n35528) );
  NOR2X1 U24530 ( .A(n25907), .B(n35529), .Y(n24026) );
  INVX1 U24531 ( .A(reg_file[1102]), .Y(n35529) );
  NOR2X1 U24532 ( .A(n25907), .B(n35530), .Y(n24025) );
  INVX1 U24533 ( .A(reg_file[1103]), .Y(n35530) );
  NOR2X1 U24534 ( .A(n25907), .B(n35531), .Y(n24024) );
  INVX1 U24535 ( .A(reg_file[1104]), .Y(n35531) );
  NOR2X1 U24536 ( .A(n25907), .B(n35532), .Y(n24023) );
  INVX1 U24537 ( .A(reg_file[1105]), .Y(n35532) );
  NOR2X1 U24538 ( .A(n25908), .B(n35533), .Y(n24022) );
  INVX1 U24539 ( .A(reg_file[1106]), .Y(n35533) );
  NOR2X1 U24540 ( .A(n25908), .B(n35534), .Y(n24021) );
  INVX1 U24541 ( .A(reg_file[1107]), .Y(n35534) );
  NOR2X1 U24542 ( .A(n25908), .B(n35535), .Y(n24020) );
  INVX1 U24543 ( .A(reg_file[1108]), .Y(n35535) );
  NOR2X1 U24544 ( .A(n25908), .B(n35536), .Y(n24019) );
  INVX1 U24545 ( .A(reg_file[1109]), .Y(n35536) );
  NOR2X1 U24546 ( .A(n25908), .B(n35537), .Y(n24018) );
  INVX1 U24547 ( .A(reg_file[1110]), .Y(n35537) );
  NOR2X1 U24548 ( .A(n25908), .B(n35538), .Y(n24017) );
  INVX1 U24549 ( .A(reg_file[1111]), .Y(n35538) );
  NOR2X1 U24550 ( .A(n25908), .B(n35539), .Y(n24016) );
  INVX1 U24551 ( .A(reg_file[1112]), .Y(n35539) );
  NOR2X1 U24552 ( .A(n25908), .B(n35540), .Y(n24015) );
  INVX1 U24553 ( .A(reg_file[1113]), .Y(n35540) );
  NOR2X1 U24554 ( .A(n25908), .B(n35541), .Y(n24014) );
  INVX1 U24555 ( .A(reg_file[1114]), .Y(n35541) );
  NOR2X1 U24556 ( .A(n25908), .B(n35542), .Y(n24013) );
  INVX1 U24557 ( .A(reg_file[1115]), .Y(n35542) );
  NOR2X1 U24558 ( .A(n25908), .B(n35543), .Y(n24012) );
  INVX1 U24559 ( .A(reg_file[1116]), .Y(n35543) );
  NOR2X1 U24560 ( .A(n25908), .B(n35544), .Y(n24011) );
  INVX1 U24561 ( .A(reg_file[1117]), .Y(n35544) );
  NOR2X1 U24562 ( .A(n25908), .B(n35545), .Y(n24010) );
  INVX1 U24563 ( .A(reg_file[1118]), .Y(n35545) );
  NOR2X1 U24564 ( .A(n25908), .B(n35546), .Y(n24009) );
  INVX1 U24565 ( .A(reg_file[1119]), .Y(n35546) );
  NOR2X1 U24566 ( .A(n25908), .B(n35547), .Y(n24008) );
  INVX1 U24567 ( .A(reg_file[1120]), .Y(n35547) );
  NOR2X1 U24568 ( .A(n25908), .B(n35548), .Y(n24007) );
  INVX1 U24569 ( .A(reg_file[1121]), .Y(n35548) );
  NOR2X1 U24570 ( .A(n25908), .B(n35549), .Y(n24006) );
  INVX1 U24571 ( .A(reg_file[1122]), .Y(n35549) );
  NOR2X1 U24572 ( .A(n25909), .B(n35550), .Y(n24005) );
  INVX1 U24573 ( .A(reg_file[1123]), .Y(n35550) );
  NOR2X1 U24574 ( .A(n25909), .B(n35551), .Y(n24004) );
  INVX1 U24575 ( .A(reg_file[1124]), .Y(n35551) );
  NOR2X1 U24576 ( .A(n25909), .B(n35552), .Y(n24003) );
  INVX1 U24577 ( .A(reg_file[1125]), .Y(n35552) );
  NOR2X1 U24578 ( .A(n25909), .B(n35553), .Y(n24002) );
  INVX1 U24579 ( .A(reg_file[1126]), .Y(n35553) );
  NOR2X1 U24580 ( .A(n25909), .B(n35554), .Y(n24001) );
  INVX1 U24581 ( .A(reg_file[1127]), .Y(n35554) );
  NOR2X1 U24582 ( .A(n25909), .B(n35555), .Y(n24000) );
  INVX1 U24583 ( .A(reg_file[1128]), .Y(n35555) );
  NOR2X1 U24584 ( .A(n25909), .B(n35556), .Y(n23999) );
  INVX1 U24585 ( .A(reg_file[1129]), .Y(n35556) );
  NOR2X1 U24586 ( .A(n25909), .B(n35557), .Y(n23998) );
  INVX1 U24587 ( .A(reg_file[1130]), .Y(n35557) );
  NOR2X1 U24588 ( .A(n25909), .B(n35558), .Y(n23997) );
  INVX1 U24589 ( .A(reg_file[1131]), .Y(n35558) );
  NOR2X1 U24590 ( .A(n25909), .B(n35559), .Y(n23996) );
  INVX1 U24591 ( .A(reg_file[1132]), .Y(n35559) );
  NOR2X1 U24592 ( .A(n25909), .B(n35560), .Y(n23995) );
  INVX1 U24593 ( .A(reg_file[1133]), .Y(n35560) );
  NOR2X1 U24594 ( .A(n25909), .B(n35561), .Y(n23994) );
  INVX1 U24595 ( .A(reg_file[1134]), .Y(n35561) );
  NOR2X1 U24596 ( .A(n25909), .B(n35562), .Y(n23993) );
  INVX1 U24597 ( .A(reg_file[1135]), .Y(n35562) );
  NOR2X1 U24598 ( .A(n25909), .B(n35563), .Y(n23992) );
  INVX1 U24599 ( .A(reg_file[1136]), .Y(n35563) );
  NOR2X1 U24600 ( .A(n25909), .B(n35564), .Y(n23991) );
  INVX1 U24601 ( .A(reg_file[1137]), .Y(n35564) );
  NOR2X1 U24602 ( .A(n25909), .B(n35565), .Y(n23990) );
  INVX1 U24603 ( .A(reg_file[1138]), .Y(n35565) );
  NOR2X1 U24604 ( .A(n25909), .B(n35566), .Y(n23989) );
  INVX1 U24605 ( .A(reg_file[1139]), .Y(n35566) );
  NOR2X1 U24606 ( .A(n25910), .B(n35567), .Y(n23988) );
  INVX1 U24607 ( .A(reg_file[1140]), .Y(n35567) );
  NOR2X1 U24608 ( .A(n25910), .B(n35568), .Y(n23987) );
  INVX1 U24609 ( .A(reg_file[1141]), .Y(n35568) );
  NOR2X1 U24610 ( .A(n25910), .B(n35569), .Y(n23986) );
  INVX1 U24611 ( .A(reg_file[1142]), .Y(n35569) );
  NOR2X1 U24612 ( .A(n25910), .B(n35570), .Y(n23985) );
  INVX1 U24613 ( .A(reg_file[1143]), .Y(n35570) );
  NOR2X1 U24614 ( .A(n25910), .B(n35571), .Y(n23984) );
  INVX1 U24615 ( .A(reg_file[1144]), .Y(n35571) );
  NOR2X1 U24616 ( .A(n25910), .B(n35572), .Y(n23983) );
  INVX1 U24617 ( .A(reg_file[1145]), .Y(n35572) );
  NOR2X1 U24618 ( .A(n25910), .B(n35573), .Y(n23982) );
  INVX1 U24619 ( .A(reg_file[1146]), .Y(n35573) );
  NOR2X1 U24620 ( .A(n25910), .B(n35574), .Y(n23981) );
  INVX1 U24621 ( .A(reg_file[1147]), .Y(n35574) );
  NOR2X1 U24622 ( .A(n25910), .B(n35575), .Y(n23980) );
  INVX1 U24623 ( .A(reg_file[1148]), .Y(n35575) );
  NOR2X1 U24624 ( .A(n25910), .B(n35576), .Y(n23979) );
  INVX1 U24625 ( .A(reg_file[1149]), .Y(n35576) );
  NOR2X1 U24626 ( .A(n25910), .B(n35577), .Y(n23978) );
  INVX1 U24627 ( .A(reg_file[1150]), .Y(n35577) );
  NOR2X1 U24628 ( .A(n25910), .B(n35578), .Y(n23977) );
  INVX1 U24629 ( .A(reg_file[1151]), .Y(n35578) );
  NOR2X1 U24630 ( .A(n35579), .B(n34923), .Y(n35451) );
  MUX2X1 U24631 ( .B(n35580), .A(n25129), .S(n25911), .Y(n23976) );
  INVX1 U24632 ( .A(reg_file[1152]), .Y(n35580) );
  MUX2X1 U24633 ( .B(n35582), .A(n25130), .S(n25911), .Y(n23975) );
  INVX1 U24634 ( .A(reg_file[1153]), .Y(n35582) );
  MUX2X1 U24635 ( .B(n35583), .A(n25131), .S(n25911), .Y(n23974) );
  INVX1 U24636 ( .A(reg_file[1154]), .Y(n35583) );
  MUX2X1 U24637 ( .B(n35584), .A(n25132), .S(n25911), .Y(n23973) );
  INVX1 U24638 ( .A(reg_file[1155]), .Y(n35584) );
  MUX2X1 U24639 ( .B(n35585), .A(n25133), .S(n25911), .Y(n23972) );
  INVX1 U24640 ( .A(reg_file[1156]), .Y(n35585) );
  MUX2X1 U24641 ( .B(n35586), .A(n25134), .S(n25911), .Y(n23971) );
  INVX1 U24642 ( .A(reg_file[1157]), .Y(n35586) );
  MUX2X1 U24643 ( .B(n35587), .A(n25135), .S(n25911), .Y(n23970) );
  INVX1 U24644 ( .A(reg_file[1158]), .Y(n35587) );
  MUX2X1 U24645 ( .B(n35588), .A(n25136), .S(n25911), .Y(n23969) );
  INVX1 U24646 ( .A(reg_file[1159]), .Y(n35588) );
  NOR2X1 U24647 ( .A(n25911), .B(n35589), .Y(n23968) );
  INVX1 U24648 ( .A(reg_file[1160]), .Y(n35589) );
  NOR2X1 U24649 ( .A(n25911), .B(n35590), .Y(n23967) );
  INVX1 U24650 ( .A(reg_file[1161]), .Y(n35590) );
  NOR2X1 U24651 ( .A(n25911), .B(n35591), .Y(n23966) );
  INVX1 U24652 ( .A(reg_file[1162]), .Y(n35591) );
  NOR2X1 U24653 ( .A(n25911), .B(n35592), .Y(n23965) );
  INVX1 U24654 ( .A(reg_file[1163]), .Y(n35592) );
  NOR2X1 U24655 ( .A(n25911), .B(n35593), .Y(n23964) );
  INVX1 U24656 ( .A(reg_file[1164]), .Y(n35593) );
  NOR2X1 U24657 ( .A(n25911), .B(n35594), .Y(n23963) );
  INVX1 U24658 ( .A(reg_file[1165]), .Y(n35594) );
  NOR2X1 U24659 ( .A(n25912), .B(n35595), .Y(n23962) );
  INVX1 U24660 ( .A(reg_file[1166]), .Y(n35595) );
  NOR2X1 U24661 ( .A(n25912), .B(n35596), .Y(n23961) );
  INVX1 U24662 ( .A(reg_file[1167]), .Y(n35596) );
  NOR2X1 U24663 ( .A(n25912), .B(n35597), .Y(n23960) );
  INVX1 U24664 ( .A(reg_file[1168]), .Y(n35597) );
  NOR2X1 U24665 ( .A(n25912), .B(n35598), .Y(n23959) );
  INVX1 U24666 ( .A(reg_file[1169]), .Y(n35598) );
  NOR2X1 U24667 ( .A(n25912), .B(n35599), .Y(n23958) );
  INVX1 U24668 ( .A(reg_file[1170]), .Y(n35599) );
  NOR2X1 U24669 ( .A(n25912), .B(n35600), .Y(n23957) );
  INVX1 U24670 ( .A(reg_file[1171]), .Y(n35600) );
  NOR2X1 U24671 ( .A(n25912), .B(n35601), .Y(n23956) );
  INVX1 U24672 ( .A(reg_file[1172]), .Y(n35601) );
  NOR2X1 U24673 ( .A(n25912), .B(n35602), .Y(n23955) );
  INVX1 U24674 ( .A(reg_file[1173]), .Y(n35602) );
  NOR2X1 U24675 ( .A(n25912), .B(n35603), .Y(n23954) );
  INVX1 U24676 ( .A(reg_file[1174]), .Y(n35603) );
  NOR2X1 U24677 ( .A(n25912), .B(n35604), .Y(n23953) );
  INVX1 U24678 ( .A(reg_file[1175]), .Y(n35604) );
  NOR2X1 U24679 ( .A(n25912), .B(n35605), .Y(n23952) );
  INVX1 U24680 ( .A(reg_file[1176]), .Y(n35605) );
  NOR2X1 U24681 ( .A(n25912), .B(n35606), .Y(n23951) );
  INVX1 U24682 ( .A(reg_file[1177]), .Y(n35606) );
  NOR2X1 U24683 ( .A(n25912), .B(n35607), .Y(n23950) );
  INVX1 U24684 ( .A(reg_file[1178]), .Y(n35607) );
  NOR2X1 U24685 ( .A(n25912), .B(n35608), .Y(n23949) );
  INVX1 U24686 ( .A(reg_file[1179]), .Y(n35608) );
  NOR2X1 U24687 ( .A(n25912), .B(n35609), .Y(n23948) );
  INVX1 U24688 ( .A(reg_file[1180]), .Y(n35609) );
  NOR2X1 U24689 ( .A(n25912), .B(n35610), .Y(n23947) );
  INVX1 U24690 ( .A(reg_file[1181]), .Y(n35610) );
  NOR2X1 U24691 ( .A(n25912), .B(n35611), .Y(n23946) );
  INVX1 U24692 ( .A(reg_file[1182]), .Y(n35611) );
  NOR2X1 U24693 ( .A(n25913), .B(n35612), .Y(n23945) );
  INVX1 U24694 ( .A(reg_file[1183]), .Y(n35612) );
  NOR2X1 U24695 ( .A(n25913), .B(n35613), .Y(n23944) );
  INVX1 U24696 ( .A(reg_file[1184]), .Y(n35613) );
  NOR2X1 U24697 ( .A(n25913), .B(n35614), .Y(n23943) );
  INVX1 U24698 ( .A(reg_file[1185]), .Y(n35614) );
  NOR2X1 U24699 ( .A(n25913), .B(n35615), .Y(n23942) );
  INVX1 U24700 ( .A(reg_file[1186]), .Y(n35615) );
  NOR2X1 U24701 ( .A(n25913), .B(n35616), .Y(n23941) );
  INVX1 U24702 ( .A(reg_file[1187]), .Y(n35616) );
  NOR2X1 U24703 ( .A(n25913), .B(n35617), .Y(n23940) );
  INVX1 U24704 ( .A(reg_file[1188]), .Y(n35617) );
  NOR2X1 U24705 ( .A(n25913), .B(n35618), .Y(n23939) );
  INVX1 U24706 ( .A(reg_file[1189]), .Y(n35618) );
  NOR2X1 U24707 ( .A(n25913), .B(n35619), .Y(n23938) );
  INVX1 U24708 ( .A(reg_file[1190]), .Y(n35619) );
  NOR2X1 U24709 ( .A(n25913), .B(n35620), .Y(n23937) );
  INVX1 U24710 ( .A(reg_file[1191]), .Y(n35620) );
  NOR2X1 U24711 ( .A(n25913), .B(n35621), .Y(n23936) );
  INVX1 U24712 ( .A(reg_file[1192]), .Y(n35621) );
  NOR2X1 U24713 ( .A(n25913), .B(n35622), .Y(n23935) );
  INVX1 U24714 ( .A(reg_file[1193]), .Y(n35622) );
  NOR2X1 U24715 ( .A(n25913), .B(n35623), .Y(n23934) );
  INVX1 U24716 ( .A(reg_file[1194]), .Y(n35623) );
  NOR2X1 U24717 ( .A(n25913), .B(n35624), .Y(n23933) );
  INVX1 U24718 ( .A(reg_file[1195]), .Y(n35624) );
  NOR2X1 U24719 ( .A(n25913), .B(n35625), .Y(n23932) );
  INVX1 U24720 ( .A(reg_file[1196]), .Y(n35625) );
  NOR2X1 U24721 ( .A(n25913), .B(n35626), .Y(n23931) );
  INVX1 U24722 ( .A(reg_file[1197]), .Y(n35626) );
  NOR2X1 U24723 ( .A(n25913), .B(n35627), .Y(n23930) );
  INVX1 U24724 ( .A(reg_file[1198]), .Y(n35627) );
  NOR2X1 U24725 ( .A(n25913), .B(n35628), .Y(n23929) );
  INVX1 U24726 ( .A(reg_file[1199]), .Y(n35628) );
  NOR2X1 U24727 ( .A(n25914), .B(n35629), .Y(n23928) );
  INVX1 U24728 ( .A(reg_file[1200]), .Y(n35629) );
  NOR2X1 U24729 ( .A(n25914), .B(n35630), .Y(n23927) );
  INVX1 U24730 ( .A(reg_file[1201]), .Y(n35630) );
  NOR2X1 U24731 ( .A(n25914), .B(n35631), .Y(n23926) );
  INVX1 U24732 ( .A(reg_file[1202]), .Y(n35631) );
  NOR2X1 U24733 ( .A(n25914), .B(n35632), .Y(n23925) );
  INVX1 U24734 ( .A(reg_file[1203]), .Y(n35632) );
  NOR2X1 U24735 ( .A(n25914), .B(n35633), .Y(n23924) );
  INVX1 U24736 ( .A(reg_file[1204]), .Y(n35633) );
  NOR2X1 U24737 ( .A(n25914), .B(n35634), .Y(n23923) );
  INVX1 U24738 ( .A(reg_file[1205]), .Y(n35634) );
  NOR2X1 U24739 ( .A(n25914), .B(n35635), .Y(n23922) );
  INVX1 U24740 ( .A(reg_file[1206]), .Y(n35635) );
  NOR2X1 U24741 ( .A(n25914), .B(n35636), .Y(n23921) );
  INVX1 U24742 ( .A(reg_file[1207]), .Y(n35636) );
  NOR2X1 U24743 ( .A(n25914), .B(n35637), .Y(n23920) );
  INVX1 U24744 ( .A(reg_file[1208]), .Y(n35637) );
  NOR2X1 U24745 ( .A(n25914), .B(n35638), .Y(n23919) );
  INVX1 U24746 ( .A(reg_file[1209]), .Y(n35638) );
  NOR2X1 U24747 ( .A(n25914), .B(n35639), .Y(n23918) );
  INVX1 U24748 ( .A(reg_file[1210]), .Y(n35639) );
  NOR2X1 U24749 ( .A(n25914), .B(n35640), .Y(n23917) );
  INVX1 U24750 ( .A(reg_file[1211]), .Y(n35640) );
  NOR2X1 U24751 ( .A(n25914), .B(n35641), .Y(n23916) );
  INVX1 U24752 ( .A(reg_file[1212]), .Y(n35641) );
  NOR2X1 U24753 ( .A(n25914), .B(n35642), .Y(n23915) );
  INVX1 U24754 ( .A(reg_file[1213]), .Y(n35642) );
  NOR2X1 U24755 ( .A(n25914), .B(n35643), .Y(n23914) );
  INVX1 U24756 ( .A(reg_file[1214]), .Y(n35643) );
  NOR2X1 U24757 ( .A(n25914), .B(n35644), .Y(n23913) );
  INVX1 U24758 ( .A(reg_file[1215]), .Y(n35644) );
  NOR2X1 U24759 ( .A(n25914), .B(n35645), .Y(n23912) );
  INVX1 U24760 ( .A(reg_file[1216]), .Y(n35645) );
  NOR2X1 U24761 ( .A(n25915), .B(n35646), .Y(n23911) );
  INVX1 U24762 ( .A(reg_file[1217]), .Y(n35646) );
  NOR2X1 U24763 ( .A(n25915), .B(n35647), .Y(n23910) );
  INVX1 U24764 ( .A(reg_file[1218]), .Y(n35647) );
  NOR2X1 U24765 ( .A(n25915), .B(n35648), .Y(n23909) );
  INVX1 U24766 ( .A(reg_file[1219]), .Y(n35648) );
  NOR2X1 U24767 ( .A(n25915), .B(n35649), .Y(n23908) );
  INVX1 U24768 ( .A(reg_file[1220]), .Y(n35649) );
  NOR2X1 U24769 ( .A(n25915), .B(n35650), .Y(n23907) );
  INVX1 U24770 ( .A(reg_file[1221]), .Y(n35650) );
  NOR2X1 U24771 ( .A(n25915), .B(n35651), .Y(n23906) );
  INVX1 U24772 ( .A(reg_file[1222]), .Y(n35651) );
  NOR2X1 U24773 ( .A(n25915), .B(n35652), .Y(n23905) );
  INVX1 U24774 ( .A(reg_file[1223]), .Y(n35652) );
  NOR2X1 U24775 ( .A(n25915), .B(n35653), .Y(n23904) );
  INVX1 U24776 ( .A(reg_file[1224]), .Y(n35653) );
  NOR2X1 U24777 ( .A(n25915), .B(n35654), .Y(n23903) );
  INVX1 U24778 ( .A(reg_file[1225]), .Y(n35654) );
  NOR2X1 U24779 ( .A(n25915), .B(n35655), .Y(n23902) );
  INVX1 U24780 ( .A(reg_file[1226]), .Y(n35655) );
  NOR2X1 U24781 ( .A(n25915), .B(n35656), .Y(n23901) );
  INVX1 U24782 ( .A(reg_file[1227]), .Y(n35656) );
  NOR2X1 U24783 ( .A(n25915), .B(n35657), .Y(n23900) );
  INVX1 U24784 ( .A(reg_file[1228]), .Y(n35657) );
  NOR2X1 U24785 ( .A(n25915), .B(n35658), .Y(n23899) );
  INVX1 U24786 ( .A(reg_file[1229]), .Y(n35658) );
  NOR2X1 U24787 ( .A(n25915), .B(n35659), .Y(n23898) );
  INVX1 U24788 ( .A(reg_file[1230]), .Y(n35659) );
  NOR2X1 U24789 ( .A(n25915), .B(n35660), .Y(n23897) );
  INVX1 U24790 ( .A(reg_file[1231]), .Y(n35660) );
  NOR2X1 U24791 ( .A(n25915), .B(n35661), .Y(n23896) );
  INVX1 U24792 ( .A(reg_file[1232]), .Y(n35661) );
  NOR2X1 U24793 ( .A(n25915), .B(n35662), .Y(n23895) );
  INVX1 U24794 ( .A(reg_file[1233]), .Y(n35662) );
  NOR2X1 U24795 ( .A(n25916), .B(n35663), .Y(n23894) );
  INVX1 U24796 ( .A(reg_file[1234]), .Y(n35663) );
  NOR2X1 U24797 ( .A(n25916), .B(n35664), .Y(n23893) );
  INVX1 U24798 ( .A(reg_file[1235]), .Y(n35664) );
  NOR2X1 U24799 ( .A(n25916), .B(n35665), .Y(n23892) );
  INVX1 U24800 ( .A(reg_file[1236]), .Y(n35665) );
  NOR2X1 U24801 ( .A(n25916), .B(n35666), .Y(n23891) );
  INVX1 U24802 ( .A(reg_file[1237]), .Y(n35666) );
  NOR2X1 U24803 ( .A(n25916), .B(n35667), .Y(n23890) );
  INVX1 U24804 ( .A(reg_file[1238]), .Y(n35667) );
  NOR2X1 U24805 ( .A(n25916), .B(n35668), .Y(n23889) );
  INVX1 U24806 ( .A(reg_file[1239]), .Y(n35668) );
  NOR2X1 U24807 ( .A(n25916), .B(n35669), .Y(n23888) );
  INVX1 U24808 ( .A(reg_file[1240]), .Y(n35669) );
  NOR2X1 U24809 ( .A(n25916), .B(n35670), .Y(n23887) );
  INVX1 U24810 ( .A(reg_file[1241]), .Y(n35670) );
  NOR2X1 U24811 ( .A(n25916), .B(n35671), .Y(n23886) );
  INVX1 U24812 ( .A(reg_file[1242]), .Y(n35671) );
  NOR2X1 U24813 ( .A(n25916), .B(n35672), .Y(n23885) );
  INVX1 U24814 ( .A(reg_file[1243]), .Y(n35672) );
  NOR2X1 U24815 ( .A(n25916), .B(n35673), .Y(n23884) );
  INVX1 U24816 ( .A(reg_file[1244]), .Y(n35673) );
  NOR2X1 U24817 ( .A(n25916), .B(n35674), .Y(n23883) );
  INVX1 U24818 ( .A(reg_file[1245]), .Y(n35674) );
  NOR2X1 U24819 ( .A(n25916), .B(n35675), .Y(n23882) );
  INVX1 U24820 ( .A(reg_file[1246]), .Y(n35675) );
  NOR2X1 U24821 ( .A(n25916), .B(n35676), .Y(n23881) );
  INVX1 U24822 ( .A(reg_file[1247]), .Y(n35676) );
  NOR2X1 U24823 ( .A(n25916), .B(n35677), .Y(n23880) );
  INVX1 U24824 ( .A(reg_file[1248]), .Y(n35677) );
  NOR2X1 U24825 ( .A(n25916), .B(n35678), .Y(n23879) );
  INVX1 U24826 ( .A(reg_file[1249]), .Y(n35678) );
  NOR2X1 U24827 ( .A(n25916), .B(n35679), .Y(n23878) );
  INVX1 U24828 ( .A(reg_file[1250]), .Y(n35679) );
  NOR2X1 U24829 ( .A(n25917), .B(n35680), .Y(n23877) );
  INVX1 U24830 ( .A(reg_file[1251]), .Y(n35680) );
  NOR2X1 U24831 ( .A(n25917), .B(n35681), .Y(n23876) );
  INVX1 U24832 ( .A(reg_file[1252]), .Y(n35681) );
  NOR2X1 U24833 ( .A(n25917), .B(n35682), .Y(n23875) );
  INVX1 U24834 ( .A(reg_file[1253]), .Y(n35682) );
  NOR2X1 U24835 ( .A(n25917), .B(n35683), .Y(n23874) );
  INVX1 U24836 ( .A(reg_file[1254]), .Y(n35683) );
  NOR2X1 U24837 ( .A(n25917), .B(n35684), .Y(n23873) );
  INVX1 U24838 ( .A(reg_file[1255]), .Y(n35684) );
  NOR2X1 U24839 ( .A(n25917), .B(n35685), .Y(n23872) );
  INVX1 U24840 ( .A(reg_file[1256]), .Y(n35685) );
  NOR2X1 U24841 ( .A(n25917), .B(n35686), .Y(n23871) );
  INVX1 U24842 ( .A(reg_file[1257]), .Y(n35686) );
  NOR2X1 U24843 ( .A(n25917), .B(n35687), .Y(n23870) );
  INVX1 U24844 ( .A(reg_file[1258]), .Y(n35687) );
  NOR2X1 U24845 ( .A(n25917), .B(n35688), .Y(n23869) );
  INVX1 U24846 ( .A(reg_file[1259]), .Y(n35688) );
  NOR2X1 U24847 ( .A(n25917), .B(n35689), .Y(n23868) );
  INVX1 U24848 ( .A(reg_file[1260]), .Y(n35689) );
  NOR2X1 U24849 ( .A(n25917), .B(n35690), .Y(n23867) );
  INVX1 U24850 ( .A(reg_file[1261]), .Y(n35690) );
  NOR2X1 U24851 ( .A(n25917), .B(n35691), .Y(n23866) );
  INVX1 U24852 ( .A(reg_file[1262]), .Y(n35691) );
  NOR2X1 U24853 ( .A(n25917), .B(n35692), .Y(n23865) );
  INVX1 U24854 ( .A(reg_file[1263]), .Y(n35692) );
  NOR2X1 U24855 ( .A(n25917), .B(n35693), .Y(n23864) );
  INVX1 U24856 ( .A(reg_file[1264]), .Y(n35693) );
  NOR2X1 U24857 ( .A(n25917), .B(n35694), .Y(n23863) );
  INVX1 U24858 ( .A(reg_file[1265]), .Y(n35694) );
  NOR2X1 U24859 ( .A(n25917), .B(n35695), .Y(n23862) );
  INVX1 U24860 ( .A(reg_file[1266]), .Y(n35695) );
  NOR2X1 U24861 ( .A(n25917), .B(n35696), .Y(n23861) );
  INVX1 U24862 ( .A(reg_file[1267]), .Y(n35696) );
  NOR2X1 U24863 ( .A(n25918), .B(n35697), .Y(n23860) );
  INVX1 U24864 ( .A(reg_file[1268]), .Y(n35697) );
  NOR2X1 U24865 ( .A(n25918), .B(n35698), .Y(n23859) );
  INVX1 U24866 ( .A(reg_file[1269]), .Y(n35698) );
  NOR2X1 U24867 ( .A(n25918), .B(n35699), .Y(n23858) );
  INVX1 U24868 ( .A(reg_file[1270]), .Y(n35699) );
  NOR2X1 U24869 ( .A(n25918), .B(n35700), .Y(n23857) );
  INVX1 U24870 ( .A(reg_file[1271]), .Y(n35700) );
  NOR2X1 U24871 ( .A(n25918), .B(n35701), .Y(n23856) );
  INVX1 U24872 ( .A(reg_file[1272]), .Y(n35701) );
  NOR2X1 U24873 ( .A(n25918), .B(n35702), .Y(n23855) );
  INVX1 U24874 ( .A(reg_file[1273]), .Y(n35702) );
  NOR2X1 U24875 ( .A(n25918), .B(n35703), .Y(n23854) );
  INVX1 U24876 ( .A(reg_file[1274]), .Y(n35703) );
  NOR2X1 U24877 ( .A(n25918), .B(n35704), .Y(n23853) );
  INVX1 U24878 ( .A(reg_file[1275]), .Y(n35704) );
  NOR2X1 U24879 ( .A(n25918), .B(n35705), .Y(n23852) );
  INVX1 U24880 ( .A(reg_file[1276]), .Y(n35705) );
  NOR2X1 U24881 ( .A(n25918), .B(n35706), .Y(n23851) );
  INVX1 U24882 ( .A(reg_file[1277]), .Y(n35706) );
  NOR2X1 U24883 ( .A(n25918), .B(n35707), .Y(n23850) );
  INVX1 U24884 ( .A(reg_file[1278]), .Y(n35707) );
  NOR2X1 U24885 ( .A(n25918), .B(n35708), .Y(n23849) );
  INVX1 U24886 ( .A(reg_file[1279]), .Y(n35708) );
  NOR2X1 U24887 ( .A(n35709), .B(n34923), .Y(n35581) );
  MUX2X1 U24888 ( .B(n35710), .A(n25129), .S(n25919), .Y(n23848) );
  INVX1 U24889 ( .A(reg_file[1280]), .Y(n35710) );
  MUX2X1 U24890 ( .B(n35712), .A(n25130), .S(n25919), .Y(n23847) );
  INVX1 U24891 ( .A(reg_file[1281]), .Y(n35712) );
  MUX2X1 U24892 ( .B(n35713), .A(n25131), .S(n25919), .Y(n23846) );
  INVX1 U24893 ( .A(reg_file[1282]), .Y(n35713) );
  MUX2X1 U24894 ( .B(n35714), .A(n25132), .S(n25919), .Y(n23845) );
  INVX1 U24895 ( .A(reg_file[1283]), .Y(n35714) );
  MUX2X1 U24896 ( .B(n35715), .A(n25133), .S(n25919), .Y(n23844) );
  INVX1 U24897 ( .A(reg_file[1284]), .Y(n35715) );
  MUX2X1 U24898 ( .B(n35716), .A(n25134), .S(n25919), .Y(n23843) );
  INVX1 U24899 ( .A(reg_file[1285]), .Y(n35716) );
  MUX2X1 U24900 ( .B(n35717), .A(n25135), .S(n25919), .Y(n23842) );
  INVX1 U24901 ( .A(reg_file[1286]), .Y(n35717) );
  MUX2X1 U24902 ( .B(n35718), .A(n25136), .S(n25919), .Y(n23841) );
  INVX1 U24903 ( .A(reg_file[1287]), .Y(n35718) );
  NOR2X1 U24904 ( .A(n25919), .B(n35719), .Y(n23840) );
  INVX1 U24905 ( .A(reg_file[1288]), .Y(n35719) );
  NOR2X1 U24906 ( .A(n25919), .B(n35720), .Y(n23839) );
  INVX1 U24907 ( .A(reg_file[1289]), .Y(n35720) );
  NOR2X1 U24908 ( .A(n25919), .B(n35721), .Y(n23838) );
  INVX1 U24909 ( .A(reg_file[1290]), .Y(n35721) );
  NOR2X1 U24910 ( .A(n25919), .B(n35722), .Y(n23837) );
  INVX1 U24911 ( .A(reg_file[1291]), .Y(n35722) );
  NOR2X1 U24912 ( .A(n25919), .B(n35723), .Y(n23836) );
  INVX1 U24913 ( .A(reg_file[1292]), .Y(n35723) );
  NOR2X1 U24914 ( .A(n25919), .B(n35724), .Y(n23835) );
  INVX1 U24915 ( .A(reg_file[1293]), .Y(n35724) );
  NOR2X1 U24916 ( .A(n25920), .B(n35725), .Y(n23834) );
  INVX1 U24917 ( .A(reg_file[1294]), .Y(n35725) );
  NOR2X1 U24918 ( .A(n25920), .B(n35726), .Y(n23833) );
  INVX1 U24919 ( .A(reg_file[1295]), .Y(n35726) );
  NOR2X1 U24920 ( .A(n25920), .B(n35727), .Y(n23832) );
  INVX1 U24921 ( .A(reg_file[1296]), .Y(n35727) );
  NOR2X1 U24922 ( .A(n25920), .B(n35728), .Y(n23831) );
  INVX1 U24923 ( .A(reg_file[1297]), .Y(n35728) );
  NOR2X1 U24924 ( .A(n25920), .B(n35729), .Y(n23830) );
  INVX1 U24925 ( .A(reg_file[1298]), .Y(n35729) );
  NOR2X1 U24926 ( .A(n25920), .B(n35730), .Y(n23829) );
  INVX1 U24927 ( .A(reg_file[1299]), .Y(n35730) );
  NOR2X1 U24928 ( .A(n25920), .B(n35731), .Y(n23828) );
  INVX1 U24929 ( .A(reg_file[1300]), .Y(n35731) );
  NOR2X1 U24930 ( .A(n25920), .B(n35732), .Y(n23827) );
  INVX1 U24931 ( .A(reg_file[1301]), .Y(n35732) );
  NOR2X1 U24932 ( .A(n25920), .B(n35733), .Y(n23826) );
  INVX1 U24933 ( .A(reg_file[1302]), .Y(n35733) );
  NOR2X1 U24934 ( .A(n25920), .B(n35734), .Y(n23825) );
  INVX1 U24935 ( .A(reg_file[1303]), .Y(n35734) );
  NOR2X1 U24936 ( .A(n25920), .B(n35735), .Y(n23824) );
  INVX1 U24937 ( .A(reg_file[1304]), .Y(n35735) );
  NOR2X1 U24938 ( .A(n25920), .B(n35736), .Y(n23823) );
  INVX1 U24939 ( .A(reg_file[1305]), .Y(n35736) );
  NOR2X1 U24940 ( .A(n25920), .B(n35737), .Y(n23822) );
  INVX1 U24941 ( .A(reg_file[1306]), .Y(n35737) );
  NOR2X1 U24942 ( .A(n25920), .B(n35738), .Y(n23821) );
  INVX1 U24943 ( .A(reg_file[1307]), .Y(n35738) );
  NOR2X1 U24944 ( .A(n25920), .B(n35739), .Y(n23820) );
  INVX1 U24945 ( .A(reg_file[1308]), .Y(n35739) );
  NOR2X1 U24946 ( .A(n25920), .B(n35740), .Y(n23819) );
  INVX1 U24947 ( .A(reg_file[1309]), .Y(n35740) );
  NOR2X1 U24948 ( .A(n25920), .B(n35741), .Y(n23818) );
  INVX1 U24949 ( .A(reg_file[1310]), .Y(n35741) );
  NOR2X1 U24950 ( .A(n25921), .B(n35742), .Y(n23817) );
  INVX1 U24951 ( .A(reg_file[1311]), .Y(n35742) );
  NOR2X1 U24952 ( .A(n25921), .B(n35743), .Y(n23816) );
  INVX1 U24953 ( .A(reg_file[1312]), .Y(n35743) );
  NOR2X1 U24954 ( .A(n25921), .B(n35744), .Y(n23815) );
  INVX1 U24955 ( .A(reg_file[1313]), .Y(n35744) );
  NOR2X1 U24956 ( .A(n25921), .B(n35745), .Y(n23814) );
  INVX1 U24957 ( .A(reg_file[1314]), .Y(n35745) );
  NOR2X1 U24958 ( .A(n25921), .B(n35746), .Y(n23813) );
  INVX1 U24959 ( .A(reg_file[1315]), .Y(n35746) );
  NOR2X1 U24960 ( .A(n25921), .B(n35747), .Y(n23812) );
  INVX1 U24961 ( .A(reg_file[1316]), .Y(n35747) );
  NOR2X1 U24962 ( .A(n25921), .B(n35748), .Y(n23811) );
  INVX1 U24963 ( .A(reg_file[1317]), .Y(n35748) );
  NOR2X1 U24964 ( .A(n25921), .B(n35749), .Y(n23810) );
  INVX1 U24965 ( .A(reg_file[1318]), .Y(n35749) );
  NOR2X1 U24966 ( .A(n25921), .B(n35750), .Y(n23809) );
  INVX1 U24967 ( .A(reg_file[1319]), .Y(n35750) );
  NOR2X1 U24968 ( .A(n25921), .B(n35751), .Y(n23808) );
  INVX1 U24969 ( .A(reg_file[1320]), .Y(n35751) );
  NOR2X1 U24970 ( .A(n25921), .B(n35752), .Y(n23807) );
  INVX1 U24971 ( .A(reg_file[1321]), .Y(n35752) );
  NOR2X1 U24972 ( .A(n25921), .B(n35753), .Y(n23806) );
  INVX1 U24973 ( .A(reg_file[1322]), .Y(n35753) );
  NOR2X1 U24974 ( .A(n25921), .B(n35754), .Y(n23805) );
  INVX1 U24975 ( .A(reg_file[1323]), .Y(n35754) );
  NOR2X1 U24976 ( .A(n25921), .B(n35755), .Y(n23804) );
  INVX1 U24977 ( .A(reg_file[1324]), .Y(n35755) );
  NOR2X1 U24978 ( .A(n25921), .B(n35756), .Y(n23803) );
  INVX1 U24979 ( .A(reg_file[1325]), .Y(n35756) );
  NOR2X1 U24980 ( .A(n25921), .B(n35757), .Y(n23802) );
  INVX1 U24981 ( .A(reg_file[1326]), .Y(n35757) );
  NOR2X1 U24982 ( .A(n25921), .B(n35758), .Y(n23801) );
  INVX1 U24983 ( .A(reg_file[1327]), .Y(n35758) );
  NOR2X1 U24984 ( .A(n25922), .B(n35759), .Y(n23800) );
  INVX1 U24985 ( .A(reg_file[1328]), .Y(n35759) );
  NOR2X1 U24986 ( .A(n25922), .B(n35760), .Y(n23799) );
  INVX1 U24987 ( .A(reg_file[1329]), .Y(n35760) );
  NOR2X1 U24988 ( .A(n25922), .B(n35761), .Y(n23798) );
  INVX1 U24989 ( .A(reg_file[1330]), .Y(n35761) );
  NOR2X1 U24990 ( .A(n25922), .B(n35762), .Y(n23797) );
  INVX1 U24991 ( .A(reg_file[1331]), .Y(n35762) );
  NOR2X1 U24992 ( .A(n25922), .B(n35763), .Y(n23796) );
  INVX1 U24993 ( .A(reg_file[1332]), .Y(n35763) );
  NOR2X1 U24994 ( .A(n25922), .B(n35764), .Y(n23795) );
  INVX1 U24995 ( .A(reg_file[1333]), .Y(n35764) );
  NOR2X1 U24996 ( .A(n25922), .B(n35765), .Y(n23794) );
  INVX1 U24997 ( .A(reg_file[1334]), .Y(n35765) );
  NOR2X1 U24998 ( .A(n25922), .B(n35766), .Y(n23793) );
  INVX1 U24999 ( .A(reg_file[1335]), .Y(n35766) );
  NOR2X1 U25000 ( .A(n25922), .B(n35767), .Y(n23792) );
  INVX1 U25001 ( .A(reg_file[1336]), .Y(n35767) );
  NOR2X1 U25002 ( .A(n25922), .B(n35768), .Y(n23791) );
  INVX1 U25003 ( .A(reg_file[1337]), .Y(n35768) );
  NOR2X1 U25004 ( .A(n25922), .B(n35769), .Y(n23790) );
  INVX1 U25005 ( .A(reg_file[1338]), .Y(n35769) );
  NOR2X1 U25006 ( .A(n25922), .B(n35770), .Y(n23789) );
  INVX1 U25007 ( .A(reg_file[1339]), .Y(n35770) );
  NOR2X1 U25008 ( .A(n25922), .B(n35771), .Y(n23788) );
  INVX1 U25009 ( .A(reg_file[1340]), .Y(n35771) );
  NOR2X1 U25010 ( .A(n25922), .B(n35772), .Y(n23787) );
  INVX1 U25011 ( .A(reg_file[1341]), .Y(n35772) );
  NOR2X1 U25012 ( .A(n25922), .B(n35773), .Y(n23786) );
  INVX1 U25013 ( .A(reg_file[1342]), .Y(n35773) );
  NOR2X1 U25014 ( .A(n25922), .B(n35774), .Y(n23785) );
  INVX1 U25015 ( .A(reg_file[1343]), .Y(n35774) );
  NOR2X1 U25016 ( .A(n25922), .B(n35775), .Y(n23784) );
  INVX1 U25017 ( .A(reg_file[1344]), .Y(n35775) );
  NOR2X1 U25018 ( .A(n25923), .B(n35776), .Y(n23783) );
  INVX1 U25019 ( .A(reg_file[1345]), .Y(n35776) );
  NOR2X1 U25020 ( .A(n25923), .B(n35777), .Y(n23782) );
  INVX1 U25021 ( .A(reg_file[1346]), .Y(n35777) );
  NOR2X1 U25022 ( .A(n25923), .B(n35778), .Y(n23781) );
  INVX1 U25023 ( .A(reg_file[1347]), .Y(n35778) );
  NOR2X1 U25024 ( .A(n25923), .B(n35779), .Y(n23780) );
  INVX1 U25025 ( .A(reg_file[1348]), .Y(n35779) );
  NOR2X1 U25026 ( .A(n25923), .B(n35780), .Y(n23779) );
  INVX1 U25027 ( .A(reg_file[1349]), .Y(n35780) );
  NOR2X1 U25028 ( .A(n25923), .B(n35781), .Y(n23778) );
  INVX1 U25029 ( .A(reg_file[1350]), .Y(n35781) );
  NOR2X1 U25030 ( .A(n25923), .B(n35782), .Y(n23777) );
  INVX1 U25031 ( .A(reg_file[1351]), .Y(n35782) );
  NOR2X1 U25032 ( .A(n25923), .B(n35783), .Y(n23776) );
  INVX1 U25033 ( .A(reg_file[1352]), .Y(n35783) );
  NOR2X1 U25034 ( .A(n25923), .B(n35784), .Y(n23775) );
  INVX1 U25035 ( .A(reg_file[1353]), .Y(n35784) );
  NOR2X1 U25036 ( .A(n25923), .B(n35785), .Y(n23774) );
  INVX1 U25037 ( .A(reg_file[1354]), .Y(n35785) );
  NOR2X1 U25038 ( .A(n25923), .B(n35786), .Y(n23773) );
  INVX1 U25039 ( .A(reg_file[1355]), .Y(n35786) );
  NOR2X1 U25040 ( .A(n25923), .B(n35787), .Y(n23772) );
  INVX1 U25041 ( .A(reg_file[1356]), .Y(n35787) );
  NOR2X1 U25042 ( .A(n25923), .B(n35788), .Y(n23771) );
  INVX1 U25043 ( .A(reg_file[1357]), .Y(n35788) );
  NOR2X1 U25044 ( .A(n25923), .B(n35789), .Y(n23770) );
  INVX1 U25045 ( .A(reg_file[1358]), .Y(n35789) );
  NOR2X1 U25046 ( .A(n25923), .B(n35790), .Y(n23769) );
  INVX1 U25047 ( .A(reg_file[1359]), .Y(n35790) );
  NOR2X1 U25048 ( .A(n25923), .B(n35791), .Y(n23768) );
  INVX1 U25049 ( .A(reg_file[1360]), .Y(n35791) );
  NOR2X1 U25050 ( .A(n25923), .B(n35792), .Y(n23767) );
  INVX1 U25051 ( .A(reg_file[1361]), .Y(n35792) );
  NOR2X1 U25052 ( .A(n25924), .B(n35793), .Y(n23766) );
  INVX1 U25053 ( .A(reg_file[1362]), .Y(n35793) );
  NOR2X1 U25054 ( .A(n25924), .B(n35794), .Y(n23765) );
  INVX1 U25055 ( .A(reg_file[1363]), .Y(n35794) );
  NOR2X1 U25056 ( .A(n25924), .B(n35795), .Y(n23764) );
  INVX1 U25057 ( .A(reg_file[1364]), .Y(n35795) );
  NOR2X1 U25058 ( .A(n25924), .B(n35796), .Y(n23763) );
  INVX1 U25059 ( .A(reg_file[1365]), .Y(n35796) );
  NOR2X1 U25060 ( .A(n25924), .B(n35797), .Y(n23762) );
  INVX1 U25061 ( .A(reg_file[1366]), .Y(n35797) );
  NOR2X1 U25062 ( .A(n25924), .B(n35798), .Y(n23761) );
  INVX1 U25063 ( .A(reg_file[1367]), .Y(n35798) );
  NOR2X1 U25064 ( .A(n25924), .B(n35799), .Y(n23760) );
  INVX1 U25065 ( .A(reg_file[1368]), .Y(n35799) );
  NOR2X1 U25066 ( .A(n25924), .B(n35800), .Y(n23759) );
  INVX1 U25067 ( .A(reg_file[1369]), .Y(n35800) );
  NOR2X1 U25068 ( .A(n25924), .B(n35801), .Y(n23758) );
  INVX1 U25069 ( .A(reg_file[1370]), .Y(n35801) );
  NOR2X1 U25070 ( .A(n25924), .B(n35802), .Y(n23757) );
  INVX1 U25071 ( .A(reg_file[1371]), .Y(n35802) );
  NOR2X1 U25072 ( .A(n25924), .B(n35803), .Y(n23756) );
  INVX1 U25073 ( .A(reg_file[1372]), .Y(n35803) );
  NOR2X1 U25074 ( .A(n25924), .B(n35804), .Y(n23755) );
  INVX1 U25075 ( .A(reg_file[1373]), .Y(n35804) );
  NOR2X1 U25076 ( .A(n25924), .B(n35805), .Y(n23754) );
  INVX1 U25077 ( .A(reg_file[1374]), .Y(n35805) );
  NOR2X1 U25078 ( .A(n25924), .B(n35806), .Y(n23753) );
  INVX1 U25079 ( .A(reg_file[1375]), .Y(n35806) );
  NOR2X1 U25080 ( .A(n25924), .B(n35807), .Y(n23752) );
  INVX1 U25081 ( .A(reg_file[1376]), .Y(n35807) );
  NOR2X1 U25082 ( .A(n25924), .B(n35808), .Y(n23751) );
  INVX1 U25083 ( .A(reg_file[1377]), .Y(n35808) );
  NOR2X1 U25084 ( .A(n25924), .B(n35809), .Y(n23750) );
  INVX1 U25085 ( .A(reg_file[1378]), .Y(n35809) );
  NOR2X1 U25086 ( .A(n25925), .B(n35810), .Y(n23749) );
  INVX1 U25087 ( .A(reg_file[1379]), .Y(n35810) );
  NOR2X1 U25088 ( .A(n25925), .B(n35811), .Y(n23748) );
  INVX1 U25089 ( .A(reg_file[1380]), .Y(n35811) );
  NOR2X1 U25090 ( .A(n25925), .B(n35812), .Y(n23747) );
  INVX1 U25091 ( .A(reg_file[1381]), .Y(n35812) );
  NOR2X1 U25092 ( .A(n25925), .B(n35813), .Y(n23746) );
  INVX1 U25093 ( .A(reg_file[1382]), .Y(n35813) );
  NOR2X1 U25094 ( .A(n25925), .B(n35814), .Y(n23745) );
  INVX1 U25095 ( .A(reg_file[1383]), .Y(n35814) );
  NOR2X1 U25096 ( .A(n25925), .B(n35815), .Y(n23744) );
  INVX1 U25097 ( .A(reg_file[1384]), .Y(n35815) );
  NOR2X1 U25098 ( .A(n25925), .B(n35816), .Y(n23743) );
  INVX1 U25099 ( .A(reg_file[1385]), .Y(n35816) );
  NOR2X1 U25100 ( .A(n25925), .B(n35817), .Y(n23742) );
  INVX1 U25101 ( .A(reg_file[1386]), .Y(n35817) );
  NOR2X1 U25102 ( .A(n25925), .B(n35818), .Y(n23741) );
  INVX1 U25103 ( .A(reg_file[1387]), .Y(n35818) );
  NOR2X1 U25104 ( .A(n25925), .B(n35819), .Y(n23740) );
  INVX1 U25105 ( .A(reg_file[1388]), .Y(n35819) );
  NOR2X1 U25106 ( .A(n25925), .B(n35820), .Y(n23739) );
  INVX1 U25107 ( .A(reg_file[1389]), .Y(n35820) );
  NOR2X1 U25108 ( .A(n25925), .B(n35821), .Y(n23738) );
  INVX1 U25109 ( .A(reg_file[1390]), .Y(n35821) );
  NOR2X1 U25110 ( .A(n25925), .B(n35822), .Y(n23737) );
  INVX1 U25111 ( .A(reg_file[1391]), .Y(n35822) );
  NOR2X1 U25112 ( .A(n25925), .B(n35823), .Y(n23736) );
  INVX1 U25113 ( .A(reg_file[1392]), .Y(n35823) );
  NOR2X1 U25114 ( .A(n25925), .B(n35824), .Y(n23735) );
  INVX1 U25115 ( .A(reg_file[1393]), .Y(n35824) );
  NOR2X1 U25116 ( .A(n25925), .B(n35825), .Y(n23734) );
  INVX1 U25117 ( .A(reg_file[1394]), .Y(n35825) );
  NOR2X1 U25118 ( .A(n25925), .B(n35826), .Y(n23733) );
  INVX1 U25119 ( .A(reg_file[1395]), .Y(n35826) );
  NOR2X1 U25120 ( .A(n25926), .B(n35827), .Y(n23732) );
  INVX1 U25121 ( .A(reg_file[1396]), .Y(n35827) );
  NOR2X1 U25122 ( .A(n25926), .B(n35828), .Y(n23731) );
  INVX1 U25123 ( .A(reg_file[1397]), .Y(n35828) );
  NOR2X1 U25124 ( .A(n25926), .B(n35829), .Y(n23730) );
  INVX1 U25125 ( .A(reg_file[1398]), .Y(n35829) );
  NOR2X1 U25126 ( .A(n25926), .B(n35830), .Y(n23729) );
  INVX1 U25127 ( .A(reg_file[1399]), .Y(n35830) );
  NOR2X1 U25128 ( .A(n25926), .B(n35831), .Y(n23728) );
  INVX1 U25129 ( .A(reg_file[1400]), .Y(n35831) );
  NOR2X1 U25130 ( .A(n25926), .B(n35832), .Y(n23727) );
  INVX1 U25131 ( .A(reg_file[1401]), .Y(n35832) );
  NOR2X1 U25132 ( .A(n25926), .B(n35833), .Y(n23726) );
  INVX1 U25133 ( .A(reg_file[1402]), .Y(n35833) );
  NOR2X1 U25134 ( .A(n25926), .B(n35834), .Y(n23725) );
  INVX1 U25135 ( .A(reg_file[1403]), .Y(n35834) );
  NOR2X1 U25136 ( .A(n25926), .B(n35835), .Y(n23724) );
  INVX1 U25137 ( .A(reg_file[1404]), .Y(n35835) );
  NOR2X1 U25138 ( .A(n25926), .B(n35836), .Y(n23723) );
  INVX1 U25139 ( .A(reg_file[1405]), .Y(n35836) );
  NOR2X1 U25140 ( .A(n25926), .B(n35837), .Y(n23722) );
  INVX1 U25141 ( .A(reg_file[1406]), .Y(n35837) );
  NOR2X1 U25142 ( .A(n25926), .B(n35838), .Y(n23721) );
  INVX1 U25143 ( .A(reg_file[1407]), .Y(n35838) );
  NOR2X1 U25144 ( .A(n35579), .B(n34927), .Y(n35711) );
  MUX2X1 U25145 ( .B(n35839), .A(n25129), .S(n25927), .Y(n23720) );
  INVX1 U25146 ( .A(reg_file[1408]), .Y(n35839) );
  MUX2X1 U25147 ( .B(n35841), .A(n25130), .S(n25927), .Y(n23719) );
  INVX1 U25148 ( .A(reg_file[1409]), .Y(n35841) );
  MUX2X1 U25149 ( .B(n35842), .A(n25131), .S(n25927), .Y(n23718) );
  INVX1 U25150 ( .A(reg_file[1410]), .Y(n35842) );
  MUX2X1 U25151 ( .B(n35843), .A(n25132), .S(n25927), .Y(n23717) );
  INVX1 U25152 ( .A(reg_file[1411]), .Y(n35843) );
  MUX2X1 U25153 ( .B(n35844), .A(n25133), .S(n25927), .Y(n23716) );
  INVX1 U25154 ( .A(reg_file[1412]), .Y(n35844) );
  MUX2X1 U25155 ( .B(n35845), .A(n25134), .S(n25927), .Y(n23715) );
  INVX1 U25156 ( .A(reg_file[1413]), .Y(n35845) );
  MUX2X1 U25157 ( .B(n35846), .A(n25135), .S(n25927), .Y(n23714) );
  INVX1 U25158 ( .A(reg_file[1414]), .Y(n35846) );
  MUX2X1 U25159 ( .B(n35847), .A(n25136), .S(n25927), .Y(n23713) );
  INVX1 U25160 ( .A(reg_file[1415]), .Y(n35847) );
  NOR2X1 U25161 ( .A(n25927), .B(n35848), .Y(n23712) );
  INVX1 U25162 ( .A(reg_file[1416]), .Y(n35848) );
  NOR2X1 U25163 ( .A(n25927), .B(n35849), .Y(n23711) );
  INVX1 U25164 ( .A(reg_file[1417]), .Y(n35849) );
  NOR2X1 U25165 ( .A(n25927), .B(n35850), .Y(n23710) );
  INVX1 U25166 ( .A(reg_file[1418]), .Y(n35850) );
  NOR2X1 U25167 ( .A(n25927), .B(n35851), .Y(n23709) );
  INVX1 U25168 ( .A(reg_file[1419]), .Y(n35851) );
  NOR2X1 U25169 ( .A(n25927), .B(n35852), .Y(n23708) );
  INVX1 U25170 ( .A(reg_file[1420]), .Y(n35852) );
  NOR2X1 U25171 ( .A(n25927), .B(n35853), .Y(n23707) );
  INVX1 U25172 ( .A(reg_file[1421]), .Y(n35853) );
  NOR2X1 U25173 ( .A(n25928), .B(n35854), .Y(n23706) );
  INVX1 U25174 ( .A(reg_file[1422]), .Y(n35854) );
  NOR2X1 U25175 ( .A(n25928), .B(n35855), .Y(n23705) );
  INVX1 U25176 ( .A(reg_file[1423]), .Y(n35855) );
  NOR2X1 U25177 ( .A(n25928), .B(n35856), .Y(n23704) );
  INVX1 U25178 ( .A(reg_file[1424]), .Y(n35856) );
  NOR2X1 U25179 ( .A(n25928), .B(n35857), .Y(n23703) );
  INVX1 U25180 ( .A(reg_file[1425]), .Y(n35857) );
  NOR2X1 U25181 ( .A(n25928), .B(n35858), .Y(n23702) );
  INVX1 U25182 ( .A(reg_file[1426]), .Y(n35858) );
  NOR2X1 U25183 ( .A(n25928), .B(n35859), .Y(n23701) );
  INVX1 U25184 ( .A(reg_file[1427]), .Y(n35859) );
  NOR2X1 U25185 ( .A(n25928), .B(n35860), .Y(n23700) );
  INVX1 U25186 ( .A(reg_file[1428]), .Y(n35860) );
  NOR2X1 U25187 ( .A(n25928), .B(n35861), .Y(n23699) );
  INVX1 U25188 ( .A(reg_file[1429]), .Y(n35861) );
  NOR2X1 U25189 ( .A(n25928), .B(n35862), .Y(n23698) );
  INVX1 U25190 ( .A(reg_file[1430]), .Y(n35862) );
  NOR2X1 U25191 ( .A(n25928), .B(n35863), .Y(n23697) );
  INVX1 U25192 ( .A(reg_file[1431]), .Y(n35863) );
  NOR2X1 U25193 ( .A(n25928), .B(n35864), .Y(n23696) );
  INVX1 U25194 ( .A(reg_file[1432]), .Y(n35864) );
  NOR2X1 U25195 ( .A(n25928), .B(n35865), .Y(n23695) );
  INVX1 U25196 ( .A(reg_file[1433]), .Y(n35865) );
  NOR2X1 U25197 ( .A(n25928), .B(n35866), .Y(n23694) );
  INVX1 U25198 ( .A(reg_file[1434]), .Y(n35866) );
  NOR2X1 U25199 ( .A(n25928), .B(n35867), .Y(n23693) );
  INVX1 U25200 ( .A(reg_file[1435]), .Y(n35867) );
  NOR2X1 U25201 ( .A(n25928), .B(n35868), .Y(n23692) );
  INVX1 U25202 ( .A(reg_file[1436]), .Y(n35868) );
  NOR2X1 U25203 ( .A(n25928), .B(n35869), .Y(n23691) );
  INVX1 U25204 ( .A(reg_file[1437]), .Y(n35869) );
  NOR2X1 U25205 ( .A(n25928), .B(n35870), .Y(n23690) );
  INVX1 U25206 ( .A(reg_file[1438]), .Y(n35870) );
  NOR2X1 U25207 ( .A(n25929), .B(n35871), .Y(n23689) );
  INVX1 U25208 ( .A(reg_file[1439]), .Y(n35871) );
  NOR2X1 U25209 ( .A(n25929), .B(n35872), .Y(n23688) );
  INVX1 U25210 ( .A(reg_file[1440]), .Y(n35872) );
  NOR2X1 U25211 ( .A(n25929), .B(n35873), .Y(n23687) );
  INVX1 U25212 ( .A(reg_file[1441]), .Y(n35873) );
  NOR2X1 U25213 ( .A(n25929), .B(n35874), .Y(n23686) );
  INVX1 U25214 ( .A(reg_file[1442]), .Y(n35874) );
  NOR2X1 U25215 ( .A(n25929), .B(n35875), .Y(n23685) );
  INVX1 U25216 ( .A(reg_file[1443]), .Y(n35875) );
  NOR2X1 U25217 ( .A(n25929), .B(n35876), .Y(n23684) );
  INVX1 U25218 ( .A(reg_file[1444]), .Y(n35876) );
  NOR2X1 U25219 ( .A(n25929), .B(n35877), .Y(n23683) );
  INVX1 U25220 ( .A(reg_file[1445]), .Y(n35877) );
  NOR2X1 U25221 ( .A(n25929), .B(n35878), .Y(n23682) );
  INVX1 U25222 ( .A(reg_file[1446]), .Y(n35878) );
  NOR2X1 U25223 ( .A(n25929), .B(n35879), .Y(n23681) );
  INVX1 U25224 ( .A(reg_file[1447]), .Y(n35879) );
  NOR2X1 U25225 ( .A(n25929), .B(n35880), .Y(n23680) );
  INVX1 U25226 ( .A(reg_file[1448]), .Y(n35880) );
  NOR2X1 U25227 ( .A(n25929), .B(n35881), .Y(n23679) );
  INVX1 U25228 ( .A(reg_file[1449]), .Y(n35881) );
  NOR2X1 U25229 ( .A(n25929), .B(n35882), .Y(n23678) );
  INVX1 U25230 ( .A(reg_file[1450]), .Y(n35882) );
  NOR2X1 U25231 ( .A(n25929), .B(n35883), .Y(n23677) );
  INVX1 U25232 ( .A(reg_file[1451]), .Y(n35883) );
  NOR2X1 U25233 ( .A(n25929), .B(n35884), .Y(n23676) );
  INVX1 U25234 ( .A(reg_file[1452]), .Y(n35884) );
  NOR2X1 U25235 ( .A(n25929), .B(n35885), .Y(n23675) );
  INVX1 U25236 ( .A(reg_file[1453]), .Y(n35885) );
  NOR2X1 U25237 ( .A(n25929), .B(n35886), .Y(n23674) );
  INVX1 U25238 ( .A(reg_file[1454]), .Y(n35886) );
  NOR2X1 U25239 ( .A(n25929), .B(n35887), .Y(n23673) );
  INVX1 U25240 ( .A(reg_file[1455]), .Y(n35887) );
  NOR2X1 U25241 ( .A(n25930), .B(n35888), .Y(n23672) );
  INVX1 U25242 ( .A(reg_file[1456]), .Y(n35888) );
  NOR2X1 U25243 ( .A(n25930), .B(n35889), .Y(n23671) );
  INVX1 U25244 ( .A(reg_file[1457]), .Y(n35889) );
  NOR2X1 U25245 ( .A(n25930), .B(n35890), .Y(n23670) );
  INVX1 U25246 ( .A(reg_file[1458]), .Y(n35890) );
  NOR2X1 U25247 ( .A(n25930), .B(n35891), .Y(n23669) );
  INVX1 U25248 ( .A(reg_file[1459]), .Y(n35891) );
  NOR2X1 U25249 ( .A(n25930), .B(n35892), .Y(n23668) );
  INVX1 U25250 ( .A(reg_file[1460]), .Y(n35892) );
  NOR2X1 U25251 ( .A(n25930), .B(n35893), .Y(n23667) );
  INVX1 U25252 ( .A(reg_file[1461]), .Y(n35893) );
  NOR2X1 U25253 ( .A(n25930), .B(n35894), .Y(n23666) );
  INVX1 U25254 ( .A(reg_file[1462]), .Y(n35894) );
  NOR2X1 U25255 ( .A(n25930), .B(n35895), .Y(n23665) );
  INVX1 U25256 ( .A(reg_file[1463]), .Y(n35895) );
  NOR2X1 U25257 ( .A(n25930), .B(n35896), .Y(n23664) );
  INVX1 U25258 ( .A(reg_file[1464]), .Y(n35896) );
  NOR2X1 U25259 ( .A(n25930), .B(n35897), .Y(n23663) );
  INVX1 U25260 ( .A(reg_file[1465]), .Y(n35897) );
  NOR2X1 U25261 ( .A(n25930), .B(n35898), .Y(n23662) );
  INVX1 U25262 ( .A(reg_file[1466]), .Y(n35898) );
  NOR2X1 U25263 ( .A(n25930), .B(n35899), .Y(n23661) );
  INVX1 U25264 ( .A(reg_file[1467]), .Y(n35899) );
  NOR2X1 U25265 ( .A(n25930), .B(n35900), .Y(n23660) );
  INVX1 U25266 ( .A(reg_file[1468]), .Y(n35900) );
  NOR2X1 U25267 ( .A(n25930), .B(n35901), .Y(n23659) );
  INVX1 U25268 ( .A(reg_file[1469]), .Y(n35901) );
  NOR2X1 U25269 ( .A(n25930), .B(n35902), .Y(n23658) );
  INVX1 U25270 ( .A(reg_file[1470]), .Y(n35902) );
  NOR2X1 U25271 ( .A(n25930), .B(n35903), .Y(n23657) );
  INVX1 U25272 ( .A(reg_file[1471]), .Y(n35903) );
  NOR2X1 U25273 ( .A(n25930), .B(n35904), .Y(n23656) );
  INVX1 U25274 ( .A(reg_file[1472]), .Y(n35904) );
  NOR2X1 U25275 ( .A(n25931), .B(n35905), .Y(n23655) );
  INVX1 U25276 ( .A(reg_file[1473]), .Y(n35905) );
  NOR2X1 U25277 ( .A(n25931), .B(n35906), .Y(n23654) );
  INVX1 U25278 ( .A(reg_file[1474]), .Y(n35906) );
  NOR2X1 U25279 ( .A(n25931), .B(n35907), .Y(n23653) );
  INVX1 U25280 ( .A(reg_file[1475]), .Y(n35907) );
  NOR2X1 U25281 ( .A(n25931), .B(n35908), .Y(n23652) );
  INVX1 U25282 ( .A(reg_file[1476]), .Y(n35908) );
  NOR2X1 U25283 ( .A(n25931), .B(n35909), .Y(n23651) );
  INVX1 U25284 ( .A(reg_file[1477]), .Y(n35909) );
  NOR2X1 U25285 ( .A(n25931), .B(n35910), .Y(n23650) );
  INVX1 U25286 ( .A(reg_file[1478]), .Y(n35910) );
  NOR2X1 U25287 ( .A(n25931), .B(n35911), .Y(n23649) );
  INVX1 U25288 ( .A(reg_file[1479]), .Y(n35911) );
  NOR2X1 U25289 ( .A(n25931), .B(n35912), .Y(n23648) );
  INVX1 U25290 ( .A(reg_file[1480]), .Y(n35912) );
  NOR2X1 U25291 ( .A(n25931), .B(n35913), .Y(n23647) );
  INVX1 U25292 ( .A(reg_file[1481]), .Y(n35913) );
  NOR2X1 U25293 ( .A(n25931), .B(n35914), .Y(n23646) );
  INVX1 U25294 ( .A(reg_file[1482]), .Y(n35914) );
  NOR2X1 U25295 ( .A(n25931), .B(n35915), .Y(n23645) );
  INVX1 U25296 ( .A(reg_file[1483]), .Y(n35915) );
  NOR2X1 U25297 ( .A(n25931), .B(n35916), .Y(n23644) );
  INVX1 U25298 ( .A(reg_file[1484]), .Y(n35916) );
  NOR2X1 U25299 ( .A(n25931), .B(n35917), .Y(n23643) );
  INVX1 U25300 ( .A(reg_file[1485]), .Y(n35917) );
  NOR2X1 U25301 ( .A(n25931), .B(n35918), .Y(n23642) );
  INVX1 U25302 ( .A(reg_file[1486]), .Y(n35918) );
  NOR2X1 U25303 ( .A(n25931), .B(n35919), .Y(n23641) );
  INVX1 U25304 ( .A(reg_file[1487]), .Y(n35919) );
  NOR2X1 U25305 ( .A(n25931), .B(n35920), .Y(n23640) );
  INVX1 U25306 ( .A(reg_file[1488]), .Y(n35920) );
  NOR2X1 U25307 ( .A(n25931), .B(n35921), .Y(n23639) );
  INVX1 U25308 ( .A(reg_file[1489]), .Y(n35921) );
  NOR2X1 U25309 ( .A(n25932), .B(n35922), .Y(n23638) );
  INVX1 U25310 ( .A(reg_file[1490]), .Y(n35922) );
  NOR2X1 U25311 ( .A(n25932), .B(n35923), .Y(n23637) );
  INVX1 U25312 ( .A(reg_file[1491]), .Y(n35923) );
  NOR2X1 U25313 ( .A(n25932), .B(n35924), .Y(n23636) );
  INVX1 U25314 ( .A(reg_file[1492]), .Y(n35924) );
  NOR2X1 U25315 ( .A(n25932), .B(n35925), .Y(n23635) );
  INVX1 U25316 ( .A(reg_file[1493]), .Y(n35925) );
  NOR2X1 U25317 ( .A(n25932), .B(n35926), .Y(n23634) );
  INVX1 U25318 ( .A(reg_file[1494]), .Y(n35926) );
  NOR2X1 U25319 ( .A(n25932), .B(n35927), .Y(n23633) );
  INVX1 U25320 ( .A(reg_file[1495]), .Y(n35927) );
  NOR2X1 U25321 ( .A(n25932), .B(n35928), .Y(n23632) );
  INVX1 U25322 ( .A(reg_file[1496]), .Y(n35928) );
  NOR2X1 U25323 ( .A(n25932), .B(n35929), .Y(n23631) );
  INVX1 U25324 ( .A(reg_file[1497]), .Y(n35929) );
  NOR2X1 U25325 ( .A(n25932), .B(n35930), .Y(n23630) );
  INVX1 U25326 ( .A(reg_file[1498]), .Y(n35930) );
  NOR2X1 U25327 ( .A(n25932), .B(n35931), .Y(n23629) );
  INVX1 U25328 ( .A(reg_file[1499]), .Y(n35931) );
  NOR2X1 U25329 ( .A(n25932), .B(n35932), .Y(n23628) );
  INVX1 U25330 ( .A(reg_file[1500]), .Y(n35932) );
  NOR2X1 U25331 ( .A(n25932), .B(n35933), .Y(n23627) );
  INVX1 U25332 ( .A(reg_file[1501]), .Y(n35933) );
  NOR2X1 U25333 ( .A(n25932), .B(n35934), .Y(n23626) );
  INVX1 U25334 ( .A(reg_file[1502]), .Y(n35934) );
  NOR2X1 U25335 ( .A(n25932), .B(n35935), .Y(n23625) );
  INVX1 U25336 ( .A(reg_file[1503]), .Y(n35935) );
  NOR2X1 U25337 ( .A(n25932), .B(n35936), .Y(n23624) );
  INVX1 U25338 ( .A(reg_file[1504]), .Y(n35936) );
  NOR2X1 U25339 ( .A(n25932), .B(n35937), .Y(n23623) );
  INVX1 U25340 ( .A(reg_file[1505]), .Y(n35937) );
  NOR2X1 U25341 ( .A(n25932), .B(n35938), .Y(n23622) );
  INVX1 U25342 ( .A(reg_file[1506]), .Y(n35938) );
  NOR2X1 U25343 ( .A(n25933), .B(n35939), .Y(n23621) );
  INVX1 U25344 ( .A(reg_file[1507]), .Y(n35939) );
  NOR2X1 U25345 ( .A(n25933), .B(n35940), .Y(n23620) );
  INVX1 U25346 ( .A(reg_file[1508]), .Y(n35940) );
  NOR2X1 U25347 ( .A(n25933), .B(n35941), .Y(n23619) );
  INVX1 U25348 ( .A(reg_file[1509]), .Y(n35941) );
  NOR2X1 U25349 ( .A(n25933), .B(n35942), .Y(n23618) );
  INVX1 U25350 ( .A(reg_file[1510]), .Y(n35942) );
  NOR2X1 U25351 ( .A(n25933), .B(n35943), .Y(n23617) );
  INVX1 U25352 ( .A(reg_file[1511]), .Y(n35943) );
  NOR2X1 U25353 ( .A(n25933), .B(n35944), .Y(n23616) );
  INVX1 U25354 ( .A(reg_file[1512]), .Y(n35944) );
  NOR2X1 U25355 ( .A(n25933), .B(n35945), .Y(n23615) );
  INVX1 U25356 ( .A(reg_file[1513]), .Y(n35945) );
  NOR2X1 U25357 ( .A(n25933), .B(n35946), .Y(n23614) );
  INVX1 U25358 ( .A(reg_file[1514]), .Y(n35946) );
  NOR2X1 U25359 ( .A(n25933), .B(n35947), .Y(n23613) );
  INVX1 U25360 ( .A(reg_file[1515]), .Y(n35947) );
  NOR2X1 U25361 ( .A(n25933), .B(n35948), .Y(n23612) );
  INVX1 U25362 ( .A(reg_file[1516]), .Y(n35948) );
  NOR2X1 U25363 ( .A(n25933), .B(n35949), .Y(n23611) );
  INVX1 U25364 ( .A(reg_file[1517]), .Y(n35949) );
  NOR2X1 U25365 ( .A(n25933), .B(n35950), .Y(n23610) );
  INVX1 U25366 ( .A(reg_file[1518]), .Y(n35950) );
  NOR2X1 U25367 ( .A(n25933), .B(n35951), .Y(n23609) );
  INVX1 U25368 ( .A(reg_file[1519]), .Y(n35951) );
  NOR2X1 U25369 ( .A(n25933), .B(n35952), .Y(n23608) );
  INVX1 U25370 ( .A(reg_file[1520]), .Y(n35952) );
  NOR2X1 U25371 ( .A(n25933), .B(n35953), .Y(n23607) );
  INVX1 U25372 ( .A(reg_file[1521]), .Y(n35953) );
  NOR2X1 U25373 ( .A(n25933), .B(n35954), .Y(n23606) );
  INVX1 U25374 ( .A(reg_file[1522]), .Y(n35954) );
  NOR2X1 U25375 ( .A(n25933), .B(n35955), .Y(n23605) );
  INVX1 U25376 ( .A(reg_file[1523]), .Y(n35955) );
  NOR2X1 U25377 ( .A(n25934), .B(n35956), .Y(n23604) );
  INVX1 U25378 ( .A(reg_file[1524]), .Y(n35956) );
  NOR2X1 U25379 ( .A(n25934), .B(n35957), .Y(n23603) );
  INVX1 U25380 ( .A(reg_file[1525]), .Y(n35957) );
  NOR2X1 U25381 ( .A(n25934), .B(n35958), .Y(n23602) );
  INVX1 U25382 ( .A(reg_file[1526]), .Y(n35958) );
  NOR2X1 U25383 ( .A(n25934), .B(n35959), .Y(n23601) );
  INVX1 U25384 ( .A(reg_file[1527]), .Y(n35959) );
  NOR2X1 U25385 ( .A(n25934), .B(n35960), .Y(n23600) );
  INVX1 U25386 ( .A(reg_file[1528]), .Y(n35960) );
  NOR2X1 U25387 ( .A(n25934), .B(n35961), .Y(n23599) );
  INVX1 U25388 ( .A(reg_file[1529]), .Y(n35961) );
  NOR2X1 U25389 ( .A(n25934), .B(n35962), .Y(n23598) );
  INVX1 U25390 ( .A(reg_file[1530]), .Y(n35962) );
  NOR2X1 U25391 ( .A(n25934), .B(n35963), .Y(n23597) );
  INVX1 U25392 ( .A(reg_file[1531]), .Y(n35963) );
  NOR2X1 U25393 ( .A(n25934), .B(n35964), .Y(n23596) );
  INVX1 U25394 ( .A(reg_file[1532]), .Y(n35964) );
  NOR2X1 U25395 ( .A(n25934), .B(n35965), .Y(n23595) );
  INVX1 U25396 ( .A(reg_file[1533]), .Y(n35965) );
  NOR2X1 U25397 ( .A(n25934), .B(n35966), .Y(n23594) );
  INVX1 U25398 ( .A(reg_file[1534]), .Y(n35966) );
  NOR2X1 U25399 ( .A(n25934), .B(n35967), .Y(n23593) );
  INVX1 U25400 ( .A(reg_file[1535]), .Y(n35967) );
  NOR2X1 U25401 ( .A(n35709), .B(n34927), .Y(n35840) );
  MUX2X1 U25402 ( .B(n31471), .A(n25129), .S(n25935), .Y(n23592) );
  INVX1 U25403 ( .A(reg_file[1536]), .Y(n31471) );
  MUX2X1 U25404 ( .B(n29833), .A(n25130), .S(n25935), .Y(n23591) );
  INVX1 U25405 ( .A(reg_file[1537]), .Y(n29833) );
  MUX2X1 U25406 ( .B(n29371), .A(n25131), .S(n25935), .Y(n23590) );
  INVX1 U25407 ( .A(reg_file[1538]), .Y(n29371) );
  MUX2X1 U25408 ( .B(n28909), .A(n25132), .S(n25935), .Y(n23589) );
  INVX1 U25409 ( .A(reg_file[1539]), .Y(n28909) );
  MUX2X1 U25410 ( .B(n28447), .A(n25133), .S(n25935), .Y(n23588) );
  INVX1 U25411 ( .A(reg_file[1540]), .Y(n28447) );
  MUX2X1 U25412 ( .B(n27985), .A(n25134), .S(n25935), .Y(n23587) );
  INVX1 U25413 ( .A(reg_file[1541]), .Y(n27985) );
  MUX2X1 U25414 ( .B(n27523), .A(n25135), .S(n25935), .Y(n23586) );
  INVX1 U25415 ( .A(reg_file[1542]), .Y(n27523) );
  MUX2X1 U25416 ( .B(n27061), .A(n25136), .S(n25935), .Y(n23585) );
  INVX1 U25417 ( .A(reg_file[1543]), .Y(n27061) );
  NOR2X1 U25418 ( .A(n25935), .B(n26599), .Y(n23584) );
  INVX1 U25419 ( .A(reg_file[1544]), .Y(n26599) );
  NOR2X1 U25420 ( .A(n25935), .B(n26106), .Y(n23583) );
  INVX1 U25421 ( .A(reg_file[1545]), .Y(n26106) );
  NOR2X1 U25422 ( .A(n25935), .B(n31009), .Y(n23582) );
  INVX1 U25423 ( .A(reg_file[1546]), .Y(n31009) );
  NOR2X1 U25424 ( .A(n25935), .B(n30547), .Y(n23581) );
  INVX1 U25425 ( .A(reg_file[1547]), .Y(n30547) );
  NOR2X1 U25426 ( .A(n25935), .B(n30169), .Y(n23580) );
  INVX1 U25427 ( .A(reg_file[1548]), .Y(n30169) );
  NOR2X1 U25428 ( .A(n25935), .B(n30127), .Y(n23579) );
  INVX1 U25429 ( .A(reg_file[1549]), .Y(n30127) );
  NOR2X1 U25430 ( .A(n25936), .B(n30085), .Y(n23578) );
  INVX1 U25431 ( .A(reg_file[1550]), .Y(n30085) );
  NOR2X1 U25432 ( .A(n25936), .B(n30043), .Y(n23577) );
  INVX1 U25433 ( .A(reg_file[1551]), .Y(n30043) );
  NOR2X1 U25434 ( .A(n25936), .B(n30001), .Y(n23576) );
  INVX1 U25435 ( .A(reg_file[1552]), .Y(n30001) );
  NOR2X1 U25436 ( .A(n25936), .B(n29959), .Y(n23575) );
  INVX1 U25437 ( .A(reg_file[1553]), .Y(n29959) );
  NOR2X1 U25438 ( .A(n25936), .B(n29917), .Y(n23574) );
  INVX1 U25439 ( .A(reg_file[1554]), .Y(n29917) );
  NOR2X1 U25440 ( .A(n25936), .B(n29875), .Y(n23573) );
  INVX1 U25441 ( .A(reg_file[1555]), .Y(n29875) );
  NOR2X1 U25442 ( .A(n25936), .B(n29791), .Y(n23572) );
  INVX1 U25443 ( .A(reg_file[1556]), .Y(n29791) );
  NOR2X1 U25444 ( .A(n25936), .B(n29749), .Y(n23571) );
  INVX1 U25445 ( .A(reg_file[1557]), .Y(n29749) );
  NOR2X1 U25446 ( .A(n25936), .B(n29707), .Y(n23570) );
  INVX1 U25447 ( .A(reg_file[1558]), .Y(n29707) );
  NOR2X1 U25448 ( .A(n25936), .B(n29665), .Y(n23569) );
  INVX1 U25449 ( .A(reg_file[1559]), .Y(n29665) );
  NOR2X1 U25450 ( .A(n25936), .B(n29623), .Y(n23568) );
  INVX1 U25451 ( .A(reg_file[1560]), .Y(n29623) );
  NOR2X1 U25452 ( .A(n25936), .B(n29581), .Y(n23567) );
  INVX1 U25453 ( .A(reg_file[1561]), .Y(n29581) );
  NOR2X1 U25454 ( .A(n25936), .B(n29539), .Y(n23566) );
  INVX1 U25455 ( .A(reg_file[1562]), .Y(n29539) );
  NOR2X1 U25456 ( .A(n25936), .B(n29497), .Y(n23565) );
  INVX1 U25457 ( .A(reg_file[1563]), .Y(n29497) );
  NOR2X1 U25458 ( .A(n25936), .B(n29455), .Y(n23564) );
  INVX1 U25459 ( .A(reg_file[1564]), .Y(n29455) );
  NOR2X1 U25460 ( .A(n25936), .B(n29413), .Y(n23563) );
  INVX1 U25461 ( .A(reg_file[1565]), .Y(n29413) );
  NOR2X1 U25462 ( .A(n25936), .B(n29329), .Y(n23562) );
  INVX1 U25463 ( .A(reg_file[1566]), .Y(n29329) );
  NOR2X1 U25464 ( .A(n25937), .B(n29287), .Y(n23561) );
  INVX1 U25465 ( .A(reg_file[1567]), .Y(n29287) );
  NOR2X1 U25466 ( .A(n25937), .B(n29245), .Y(n23560) );
  INVX1 U25467 ( .A(reg_file[1568]), .Y(n29245) );
  NOR2X1 U25468 ( .A(n25937), .B(n29203), .Y(n23559) );
  INVX1 U25469 ( .A(reg_file[1569]), .Y(n29203) );
  NOR2X1 U25470 ( .A(n25937), .B(n29161), .Y(n23558) );
  INVX1 U25471 ( .A(reg_file[1570]), .Y(n29161) );
  NOR2X1 U25472 ( .A(n25937), .B(n29119), .Y(n23557) );
  INVX1 U25473 ( .A(reg_file[1571]), .Y(n29119) );
  NOR2X1 U25474 ( .A(n25937), .B(n29077), .Y(n23556) );
  INVX1 U25475 ( .A(reg_file[1572]), .Y(n29077) );
  NOR2X1 U25476 ( .A(n25937), .B(n29035), .Y(n23555) );
  INVX1 U25477 ( .A(reg_file[1573]), .Y(n29035) );
  NOR2X1 U25478 ( .A(n25937), .B(n28993), .Y(n23554) );
  INVX1 U25479 ( .A(reg_file[1574]), .Y(n28993) );
  NOR2X1 U25480 ( .A(n25937), .B(n28951), .Y(n23553) );
  INVX1 U25481 ( .A(reg_file[1575]), .Y(n28951) );
  NOR2X1 U25482 ( .A(n25937), .B(n28867), .Y(n23552) );
  INVX1 U25483 ( .A(reg_file[1576]), .Y(n28867) );
  NOR2X1 U25484 ( .A(n25937), .B(n28825), .Y(n23551) );
  INVX1 U25485 ( .A(reg_file[1577]), .Y(n28825) );
  NOR2X1 U25486 ( .A(n25937), .B(n28783), .Y(n23550) );
  INVX1 U25487 ( .A(reg_file[1578]), .Y(n28783) );
  NOR2X1 U25488 ( .A(n25937), .B(n28741), .Y(n23549) );
  INVX1 U25489 ( .A(reg_file[1579]), .Y(n28741) );
  NOR2X1 U25490 ( .A(n25937), .B(n28699), .Y(n23548) );
  INVX1 U25491 ( .A(reg_file[1580]), .Y(n28699) );
  NOR2X1 U25492 ( .A(n25937), .B(n28657), .Y(n23547) );
  INVX1 U25493 ( .A(reg_file[1581]), .Y(n28657) );
  NOR2X1 U25494 ( .A(n25937), .B(n28615), .Y(n23546) );
  INVX1 U25495 ( .A(reg_file[1582]), .Y(n28615) );
  NOR2X1 U25496 ( .A(n25937), .B(n28573), .Y(n23545) );
  INVX1 U25497 ( .A(reg_file[1583]), .Y(n28573) );
  NOR2X1 U25498 ( .A(n25938), .B(n28531), .Y(n23544) );
  INVX1 U25499 ( .A(reg_file[1584]), .Y(n28531) );
  NOR2X1 U25500 ( .A(n25938), .B(n28489), .Y(n23543) );
  INVX1 U25501 ( .A(reg_file[1585]), .Y(n28489) );
  NOR2X1 U25502 ( .A(n25938), .B(n28405), .Y(n23542) );
  INVX1 U25503 ( .A(reg_file[1586]), .Y(n28405) );
  NOR2X1 U25504 ( .A(n25938), .B(n28363), .Y(n23541) );
  INVX1 U25505 ( .A(reg_file[1587]), .Y(n28363) );
  NOR2X1 U25506 ( .A(n25938), .B(n28321), .Y(n23540) );
  INVX1 U25507 ( .A(reg_file[1588]), .Y(n28321) );
  NOR2X1 U25508 ( .A(n25938), .B(n28279), .Y(n23539) );
  INVX1 U25509 ( .A(reg_file[1589]), .Y(n28279) );
  NOR2X1 U25510 ( .A(n25938), .B(n28237), .Y(n23538) );
  INVX1 U25511 ( .A(reg_file[1590]), .Y(n28237) );
  NOR2X1 U25512 ( .A(n25938), .B(n28195), .Y(n23537) );
  INVX1 U25513 ( .A(reg_file[1591]), .Y(n28195) );
  NOR2X1 U25514 ( .A(n25938), .B(n28153), .Y(n23536) );
  INVX1 U25515 ( .A(reg_file[1592]), .Y(n28153) );
  NOR2X1 U25516 ( .A(n25938), .B(n28111), .Y(n23535) );
  INVX1 U25517 ( .A(reg_file[1593]), .Y(n28111) );
  NOR2X1 U25518 ( .A(n25938), .B(n28069), .Y(n23534) );
  INVX1 U25519 ( .A(reg_file[1594]), .Y(n28069) );
  NOR2X1 U25520 ( .A(n25938), .B(n28027), .Y(n23533) );
  INVX1 U25521 ( .A(reg_file[1595]), .Y(n28027) );
  NOR2X1 U25522 ( .A(n25938), .B(n27943), .Y(n23532) );
  INVX1 U25523 ( .A(reg_file[1596]), .Y(n27943) );
  NOR2X1 U25524 ( .A(n25938), .B(n27901), .Y(n23531) );
  INVX1 U25525 ( .A(reg_file[1597]), .Y(n27901) );
  NOR2X1 U25526 ( .A(n25938), .B(n27859), .Y(n23530) );
  INVX1 U25527 ( .A(reg_file[1598]), .Y(n27859) );
  NOR2X1 U25528 ( .A(n25938), .B(n27817), .Y(n23529) );
  INVX1 U25529 ( .A(reg_file[1599]), .Y(n27817) );
  NOR2X1 U25530 ( .A(n25938), .B(n27775), .Y(n23528) );
  INVX1 U25531 ( .A(reg_file[1600]), .Y(n27775) );
  NOR2X1 U25532 ( .A(n25939), .B(n27733), .Y(n23527) );
  INVX1 U25533 ( .A(reg_file[1601]), .Y(n27733) );
  NOR2X1 U25534 ( .A(n25939), .B(n27691), .Y(n23526) );
  INVX1 U25535 ( .A(reg_file[1602]), .Y(n27691) );
  NOR2X1 U25536 ( .A(n25939), .B(n27649), .Y(n23525) );
  INVX1 U25537 ( .A(reg_file[1603]), .Y(n27649) );
  NOR2X1 U25538 ( .A(n25939), .B(n27607), .Y(n23524) );
  INVX1 U25539 ( .A(reg_file[1604]), .Y(n27607) );
  NOR2X1 U25540 ( .A(n25939), .B(n27565), .Y(n23523) );
  INVX1 U25541 ( .A(reg_file[1605]), .Y(n27565) );
  NOR2X1 U25542 ( .A(n25939), .B(n27481), .Y(n23522) );
  INVX1 U25543 ( .A(reg_file[1606]), .Y(n27481) );
  NOR2X1 U25544 ( .A(n25939), .B(n27439), .Y(n23521) );
  INVX1 U25545 ( .A(reg_file[1607]), .Y(n27439) );
  NOR2X1 U25546 ( .A(n25939), .B(n27397), .Y(n23520) );
  INVX1 U25547 ( .A(reg_file[1608]), .Y(n27397) );
  NOR2X1 U25548 ( .A(n25939), .B(n27355), .Y(n23519) );
  INVX1 U25549 ( .A(reg_file[1609]), .Y(n27355) );
  NOR2X1 U25550 ( .A(n25939), .B(n27313), .Y(n23518) );
  INVX1 U25551 ( .A(reg_file[1610]), .Y(n27313) );
  NOR2X1 U25552 ( .A(n25939), .B(n27271), .Y(n23517) );
  INVX1 U25553 ( .A(reg_file[1611]), .Y(n27271) );
  NOR2X1 U25554 ( .A(n25939), .B(n27229), .Y(n23516) );
  INVX1 U25555 ( .A(reg_file[1612]), .Y(n27229) );
  NOR2X1 U25556 ( .A(n25939), .B(n27187), .Y(n23515) );
  INVX1 U25557 ( .A(reg_file[1613]), .Y(n27187) );
  NOR2X1 U25558 ( .A(n25939), .B(n27145), .Y(n23514) );
  INVX1 U25559 ( .A(reg_file[1614]), .Y(n27145) );
  NOR2X1 U25560 ( .A(n25939), .B(n27103), .Y(n23513) );
  INVX1 U25561 ( .A(reg_file[1615]), .Y(n27103) );
  NOR2X1 U25562 ( .A(n25939), .B(n27019), .Y(n23512) );
  INVX1 U25563 ( .A(reg_file[1616]), .Y(n27019) );
  NOR2X1 U25564 ( .A(n25939), .B(n26977), .Y(n23511) );
  INVX1 U25565 ( .A(reg_file[1617]), .Y(n26977) );
  NOR2X1 U25566 ( .A(n25940), .B(n26935), .Y(n23510) );
  INVX1 U25567 ( .A(reg_file[1618]), .Y(n26935) );
  NOR2X1 U25568 ( .A(n25940), .B(n26893), .Y(n23509) );
  INVX1 U25569 ( .A(reg_file[1619]), .Y(n26893) );
  NOR2X1 U25570 ( .A(n25940), .B(n26851), .Y(n23508) );
  INVX1 U25571 ( .A(reg_file[1620]), .Y(n26851) );
  NOR2X1 U25572 ( .A(n25940), .B(n26809), .Y(n23507) );
  INVX1 U25573 ( .A(reg_file[1621]), .Y(n26809) );
  NOR2X1 U25574 ( .A(n25940), .B(n26767), .Y(n23506) );
  INVX1 U25575 ( .A(reg_file[1622]), .Y(n26767) );
  NOR2X1 U25576 ( .A(n25940), .B(n26725), .Y(n23505) );
  INVX1 U25577 ( .A(reg_file[1623]), .Y(n26725) );
  NOR2X1 U25578 ( .A(n25940), .B(n26683), .Y(n23504) );
  INVX1 U25579 ( .A(reg_file[1624]), .Y(n26683) );
  NOR2X1 U25580 ( .A(n25940), .B(n26641), .Y(n23503) );
  INVX1 U25581 ( .A(reg_file[1625]), .Y(n26641) );
  NOR2X1 U25582 ( .A(n25940), .B(n26557), .Y(n23502) );
  INVX1 U25583 ( .A(reg_file[1626]), .Y(n26557) );
  NOR2X1 U25584 ( .A(n25940), .B(n26515), .Y(n23501) );
  INVX1 U25585 ( .A(reg_file[1627]), .Y(n26515) );
  NOR2X1 U25586 ( .A(n25940), .B(n26473), .Y(n23500) );
  INVX1 U25587 ( .A(reg_file[1628]), .Y(n26473) );
  NOR2X1 U25588 ( .A(n25940), .B(n26431), .Y(n23499) );
  INVX1 U25589 ( .A(reg_file[1629]), .Y(n26431) );
  NOR2X1 U25590 ( .A(n25940), .B(n26389), .Y(n23498) );
  INVX1 U25591 ( .A(reg_file[1630]), .Y(n26389) );
  NOR2X1 U25592 ( .A(n25940), .B(n26347), .Y(n23497) );
  INVX1 U25593 ( .A(reg_file[1631]), .Y(n26347) );
  NOR2X1 U25594 ( .A(n25940), .B(n26305), .Y(n23496) );
  INVX1 U25595 ( .A(reg_file[1632]), .Y(n26305) );
  NOR2X1 U25596 ( .A(n25940), .B(n26263), .Y(n23495) );
  INVX1 U25597 ( .A(reg_file[1633]), .Y(n26263) );
  NOR2X1 U25598 ( .A(n25940), .B(n26221), .Y(n23494) );
  INVX1 U25599 ( .A(reg_file[1634]), .Y(n26221) );
  NOR2X1 U25600 ( .A(n25941), .B(n26179), .Y(n23493) );
  INVX1 U25601 ( .A(reg_file[1635]), .Y(n26179) );
  NOR2X1 U25602 ( .A(n25941), .B(n31429), .Y(n23492) );
  INVX1 U25603 ( .A(reg_file[1636]), .Y(n31429) );
  NOR2X1 U25604 ( .A(n25941), .B(n31387), .Y(n23491) );
  INVX1 U25605 ( .A(reg_file[1637]), .Y(n31387) );
  NOR2X1 U25606 ( .A(n25941), .B(n31345), .Y(n23490) );
  INVX1 U25607 ( .A(reg_file[1638]), .Y(n31345) );
  NOR2X1 U25608 ( .A(n25941), .B(n31303), .Y(n23489) );
  INVX1 U25609 ( .A(reg_file[1639]), .Y(n31303) );
  NOR2X1 U25610 ( .A(n25941), .B(n31261), .Y(n23488) );
  INVX1 U25611 ( .A(reg_file[1640]), .Y(n31261) );
  NOR2X1 U25612 ( .A(n25941), .B(n31219), .Y(n23487) );
  INVX1 U25613 ( .A(reg_file[1641]), .Y(n31219) );
  NOR2X1 U25614 ( .A(n25941), .B(n31177), .Y(n23486) );
  INVX1 U25615 ( .A(reg_file[1642]), .Y(n31177) );
  NOR2X1 U25616 ( .A(n25941), .B(n31135), .Y(n23485) );
  INVX1 U25617 ( .A(reg_file[1643]), .Y(n31135) );
  NOR2X1 U25618 ( .A(n25941), .B(n31093), .Y(n23484) );
  INVX1 U25619 ( .A(reg_file[1644]), .Y(n31093) );
  NOR2X1 U25620 ( .A(n25941), .B(n31051), .Y(n23483) );
  INVX1 U25621 ( .A(reg_file[1645]), .Y(n31051) );
  NOR2X1 U25622 ( .A(n25941), .B(n30967), .Y(n23482) );
  INVX1 U25623 ( .A(reg_file[1646]), .Y(n30967) );
  NOR2X1 U25624 ( .A(n25941), .B(n30925), .Y(n23481) );
  INVX1 U25625 ( .A(reg_file[1647]), .Y(n30925) );
  NOR2X1 U25626 ( .A(n25941), .B(n30883), .Y(n23480) );
  INVX1 U25627 ( .A(reg_file[1648]), .Y(n30883) );
  NOR2X1 U25628 ( .A(n25941), .B(n30841), .Y(n23479) );
  INVX1 U25629 ( .A(reg_file[1649]), .Y(n30841) );
  NOR2X1 U25630 ( .A(n25941), .B(n30799), .Y(n23478) );
  INVX1 U25631 ( .A(reg_file[1650]), .Y(n30799) );
  NOR2X1 U25632 ( .A(n25941), .B(n30757), .Y(n23477) );
  INVX1 U25633 ( .A(reg_file[1651]), .Y(n30757) );
  NOR2X1 U25634 ( .A(n25942), .B(n30715), .Y(n23476) );
  INVX1 U25635 ( .A(reg_file[1652]), .Y(n30715) );
  NOR2X1 U25636 ( .A(n25942), .B(n30673), .Y(n23475) );
  INVX1 U25637 ( .A(reg_file[1653]), .Y(n30673) );
  NOR2X1 U25638 ( .A(n25942), .B(n30631), .Y(n23474) );
  INVX1 U25639 ( .A(reg_file[1654]), .Y(n30631) );
  NOR2X1 U25640 ( .A(n25942), .B(n30589), .Y(n23473) );
  INVX1 U25641 ( .A(reg_file[1655]), .Y(n30589) );
  NOR2X1 U25642 ( .A(n25942), .B(n30505), .Y(n23472) );
  INVX1 U25643 ( .A(reg_file[1656]), .Y(n30505) );
  NOR2X1 U25644 ( .A(n25942), .B(n30463), .Y(n23471) );
  INVX1 U25645 ( .A(reg_file[1657]), .Y(n30463) );
  NOR2X1 U25646 ( .A(n25942), .B(n30421), .Y(n23470) );
  INVX1 U25647 ( .A(reg_file[1658]), .Y(n30421) );
  NOR2X1 U25648 ( .A(n25942), .B(n30379), .Y(n23469) );
  INVX1 U25649 ( .A(reg_file[1659]), .Y(n30379) );
  NOR2X1 U25650 ( .A(n25942), .B(n30337), .Y(n23468) );
  INVX1 U25651 ( .A(reg_file[1660]), .Y(n30337) );
  NOR2X1 U25652 ( .A(n25942), .B(n30295), .Y(n23467) );
  INVX1 U25653 ( .A(reg_file[1661]), .Y(n30295) );
  NOR2X1 U25654 ( .A(n25942), .B(n30253), .Y(n23466) );
  INVX1 U25655 ( .A(reg_file[1662]), .Y(n30253) );
  NOR2X1 U25656 ( .A(n25942), .B(n30211), .Y(n23465) );
  INVX1 U25657 ( .A(reg_file[1663]), .Y(n30211) );
  NOR2X1 U25658 ( .A(n35579), .B(n35058), .Y(n35968) );
  MUX2X1 U25659 ( .B(n31472), .A(n25129), .S(n25943), .Y(n23464) );
  INVX1 U25660 ( .A(reg_file[1664]), .Y(n31472) );
  MUX2X1 U25661 ( .B(n29834), .A(n25130), .S(n25943), .Y(n23463) );
  INVX1 U25662 ( .A(reg_file[1665]), .Y(n29834) );
  MUX2X1 U25663 ( .B(n29372), .A(n25131), .S(n25943), .Y(n23462) );
  INVX1 U25664 ( .A(reg_file[1666]), .Y(n29372) );
  MUX2X1 U25665 ( .B(n28910), .A(n25132), .S(n25943), .Y(n23461) );
  INVX1 U25666 ( .A(reg_file[1667]), .Y(n28910) );
  MUX2X1 U25667 ( .B(n28448), .A(n25133), .S(n25943), .Y(n23460) );
  INVX1 U25668 ( .A(reg_file[1668]), .Y(n28448) );
  MUX2X1 U25669 ( .B(n27986), .A(n25134), .S(n25943), .Y(n23459) );
  INVX1 U25670 ( .A(reg_file[1669]), .Y(n27986) );
  MUX2X1 U25671 ( .B(n27524), .A(n25135), .S(n25943), .Y(n23458) );
  INVX1 U25672 ( .A(reg_file[1670]), .Y(n27524) );
  MUX2X1 U25673 ( .B(n27062), .A(n25136), .S(n25943), .Y(n23457) );
  INVX1 U25674 ( .A(reg_file[1671]), .Y(n27062) );
  NOR2X1 U25675 ( .A(n25943), .B(n26600), .Y(n23456) );
  INVX1 U25676 ( .A(reg_file[1672]), .Y(n26600) );
  NOR2X1 U25677 ( .A(n25943), .B(n26108), .Y(n23455) );
  INVX1 U25678 ( .A(reg_file[1673]), .Y(n26108) );
  NOR2X1 U25679 ( .A(n25943), .B(n31010), .Y(n23454) );
  INVX1 U25680 ( .A(reg_file[1674]), .Y(n31010) );
  NOR2X1 U25681 ( .A(n25943), .B(n30548), .Y(n23453) );
  INVX1 U25682 ( .A(reg_file[1675]), .Y(n30548) );
  NOR2X1 U25683 ( .A(n25943), .B(n30170), .Y(n23452) );
  INVX1 U25684 ( .A(reg_file[1676]), .Y(n30170) );
  NOR2X1 U25685 ( .A(n25943), .B(n30128), .Y(n23451) );
  INVX1 U25686 ( .A(reg_file[1677]), .Y(n30128) );
  NOR2X1 U25687 ( .A(n25944), .B(n30086), .Y(n23450) );
  INVX1 U25688 ( .A(reg_file[1678]), .Y(n30086) );
  NOR2X1 U25689 ( .A(n25944), .B(n30044), .Y(n23449) );
  INVX1 U25690 ( .A(reg_file[1679]), .Y(n30044) );
  NOR2X1 U25691 ( .A(n25944), .B(n30002), .Y(n23448) );
  INVX1 U25692 ( .A(reg_file[1680]), .Y(n30002) );
  NOR2X1 U25693 ( .A(n25944), .B(n29960), .Y(n23447) );
  INVX1 U25694 ( .A(reg_file[1681]), .Y(n29960) );
  NOR2X1 U25695 ( .A(n25944), .B(n29918), .Y(n23446) );
  INVX1 U25696 ( .A(reg_file[1682]), .Y(n29918) );
  NOR2X1 U25697 ( .A(n25944), .B(n29876), .Y(n23445) );
  INVX1 U25698 ( .A(reg_file[1683]), .Y(n29876) );
  NOR2X1 U25699 ( .A(n25944), .B(n29792), .Y(n23444) );
  INVX1 U25700 ( .A(reg_file[1684]), .Y(n29792) );
  NOR2X1 U25701 ( .A(n25944), .B(n29750), .Y(n23443) );
  INVX1 U25702 ( .A(reg_file[1685]), .Y(n29750) );
  NOR2X1 U25703 ( .A(n25944), .B(n29708), .Y(n23442) );
  INVX1 U25704 ( .A(reg_file[1686]), .Y(n29708) );
  NOR2X1 U25705 ( .A(n25944), .B(n29666), .Y(n23441) );
  INVX1 U25706 ( .A(reg_file[1687]), .Y(n29666) );
  NOR2X1 U25707 ( .A(n25944), .B(n29624), .Y(n23440) );
  INVX1 U25708 ( .A(reg_file[1688]), .Y(n29624) );
  NOR2X1 U25709 ( .A(n25944), .B(n29582), .Y(n23439) );
  INVX1 U25710 ( .A(reg_file[1689]), .Y(n29582) );
  NOR2X1 U25711 ( .A(n25944), .B(n29540), .Y(n23438) );
  INVX1 U25712 ( .A(reg_file[1690]), .Y(n29540) );
  NOR2X1 U25713 ( .A(n25944), .B(n29498), .Y(n23437) );
  INVX1 U25714 ( .A(reg_file[1691]), .Y(n29498) );
  NOR2X1 U25715 ( .A(n25944), .B(n29456), .Y(n23436) );
  INVX1 U25716 ( .A(reg_file[1692]), .Y(n29456) );
  NOR2X1 U25717 ( .A(n25944), .B(n29414), .Y(n23435) );
  INVX1 U25718 ( .A(reg_file[1693]), .Y(n29414) );
  NOR2X1 U25719 ( .A(n25944), .B(n29330), .Y(n23434) );
  INVX1 U25720 ( .A(reg_file[1694]), .Y(n29330) );
  NOR2X1 U25721 ( .A(n25945), .B(n29288), .Y(n23433) );
  INVX1 U25722 ( .A(reg_file[1695]), .Y(n29288) );
  NOR2X1 U25723 ( .A(n25945), .B(n29246), .Y(n23432) );
  INVX1 U25724 ( .A(reg_file[1696]), .Y(n29246) );
  NOR2X1 U25725 ( .A(n25945), .B(n29204), .Y(n23431) );
  INVX1 U25726 ( .A(reg_file[1697]), .Y(n29204) );
  NOR2X1 U25727 ( .A(n25945), .B(n29162), .Y(n23430) );
  INVX1 U25728 ( .A(reg_file[1698]), .Y(n29162) );
  NOR2X1 U25729 ( .A(n25945), .B(n29120), .Y(n23429) );
  INVX1 U25730 ( .A(reg_file[1699]), .Y(n29120) );
  NOR2X1 U25731 ( .A(n25945), .B(n29078), .Y(n23428) );
  INVX1 U25732 ( .A(reg_file[1700]), .Y(n29078) );
  NOR2X1 U25733 ( .A(n25945), .B(n29036), .Y(n23427) );
  INVX1 U25734 ( .A(reg_file[1701]), .Y(n29036) );
  NOR2X1 U25735 ( .A(n25945), .B(n28994), .Y(n23426) );
  INVX1 U25736 ( .A(reg_file[1702]), .Y(n28994) );
  NOR2X1 U25737 ( .A(n25945), .B(n28952), .Y(n23425) );
  INVX1 U25738 ( .A(reg_file[1703]), .Y(n28952) );
  NOR2X1 U25739 ( .A(n25945), .B(n28868), .Y(n23424) );
  INVX1 U25740 ( .A(reg_file[1704]), .Y(n28868) );
  NOR2X1 U25741 ( .A(n25945), .B(n28826), .Y(n23423) );
  INVX1 U25742 ( .A(reg_file[1705]), .Y(n28826) );
  NOR2X1 U25743 ( .A(n25945), .B(n28784), .Y(n23422) );
  INVX1 U25744 ( .A(reg_file[1706]), .Y(n28784) );
  NOR2X1 U25745 ( .A(n25945), .B(n28742), .Y(n23421) );
  INVX1 U25746 ( .A(reg_file[1707]), .Y(n28742) );
  NOR2X1 U25747 ( .A(n25945), .B(n28700), .Y(n23420) );
  INVX1 U25748 ( .A(reg_file[1708]), .Y(n28700) );
  NOR2X1 U25749 ( .A(n25945), .B(n28658), .Y(n23419) );
  INVX1 U25750 ( .A(reg_file[1709]), .Y(n28658) );
  NOR2X1 U25751 ( .A(n25945), .B(n28616), .Y(n23418) );
  INVX1 U25752 ( .A(reg_file[1710]), .Y(n28616) );
  NOR2X1 U25753 ( .A(n25945), .B(n28574), .Y(n23417) );
  INVX1 U25754 ( .A(reg_file[1711]), .Y(n28574) );
  NOR2X1 U25755 ( .A(n25946), .B(n28532), .Y(n23416) );
  INVX1 U25756 ( .A(reg_file[1712]), .Y(n28532) );
  NOR2X1 U25757 ( .A(n25946), .B(n28490), .Y(n23415) );
  INVX1 U25758 ( .A(reg_file[1713]), .Y(n28490) );
  NOR2X1 U25759 ( .A(n25946), .B(n28406), .Y(n23414) );
  INVX1 U25760 ( .A(reg_file[1714]), .Y(n28406) );
  NOR2X1 U25761 ( .A(n25946), .B(n28364), .Y(n23413) );
  INVX1 U25762 ( .A(reg_file[1715]), .Y(n28364) );
  NOR2X1 U25763 ( .A(n25946), .B(n28322), .Y(n23412) );
  INVX1 U25764 ( .A(reg_file[1716]), .Y(n28322) );
  NOR2X1 U25765 ( .A(n25946), .B(n28280), .Y(n23411) );
  INVX1 U25766 ( .A(reg_file[1717]), .Y(n28280) );
  NOR2X1 U25767 ( .A(n25946), .B(n28238), .Y(n23410) );
  INVX1 U25768 ( .A(reg_file[1718]), .Y(n28238) );
  NOR2X1 U25769 ( .A(n25946), .B(n28196), .Y(n23409) );
  INVX1 U25770 ( .A(reg_file[1719]), .Y(n28196) );
  NOR2X1 U25771 ( .A(n25946), .B(n28154), .Y(n23408) );
  INVX1 U25772 ( .A(reg_file[1720]), .Y(n28154) );
  NOR2X1 U25773 ( .A(n25946), .B(n28112), .Y(n23407) );
  INVX1 U25774 ( .A(reg_file[1721]), .Y(n28112) );
  NOR2X1 U25775 ( .A(n25946), .B(n28070), .Y(n23406) );
  INVX1 U25776 ( .A(reg_file[1722]), .Y(n28070) );
  NOR2X1 U25777 ( .A(n25946), .B(n28028), .Y(n23405) );
  INVX1 U25778 ( .A(reg_file[1723]), .Y(n28028) );
  NOR2X1 U25779 ( .A(n25946), .B(n27944), .Y(n23404) );
  INVX1 U25780 ( .A(reg_file[1724]), .Y(n27944) );
  NOR2X1 U25781 ( .A(n25946), .B(n27902), .Y(n23403) );
  INVX1 U25782 ( .A(reg_file[1725]), .Y(n27902) );
  NOR2X1 U25783 ( .A(n25946), .B(n27860), .Y(n23402) );
  INVX1 U25784 ( .A(reg_file[1726]), .Y(n27860) );
  NOR2X1 U25785 ( .A(n25946), .B(n27818), .Y(n23401) );
  INVX1 U25786 ( .A(reg_file[1727]), .Y(n27818) );
  NOR2X1 U25787 ( .A(n25946), .B(n27776), .Y(n23400) );
  INVX1 U25788 ( .A(reg_file[1728]), .Y(n27776) );
  NOR2X1 U25789 ( .A(n25947), .B(n27734), .Y(n23399) );
  INVX1 U25790 ( .A(reg_file[1729]), .Y(n27734) );
  NOR2X1 U25791 ( .A(n25947), .B(n27692), .Y(n23398) );
  INVX1 U25792 ( .A(reg_file[1730]), .Y(n27692) );
  NOR2X1 U25793 ( .A(n25947), .B(n27650), .Y(n23397) );
  INVX1 U25794 ( .A(reg_file[1731]), .Y(n27650) );
  NOR2X1 U25795 ( .A(n25947), .B(n27608), .Y(n23396) );
  INVX1 U25796 ( .A(reg_file[1732]), .Y(n27608) );
  NOR2X1 U25797 ( .A(n25947), .B(n27566), .Y(n23395) );
  INVX1 U25798 ( .A(reg_file[1733]), .Y(n27566) );
  NOR2X1 U25799 ( .A(n25947), .B(n27482), .Y(n23394) );
  INVX1 U25800 ( .A(reg_file[1734]), .Y(n27482) );
  NOR2X1 U25801 ( .A(n25947), .B(n27440), .Y(n23393) );
  INVX1 U25802 ( .A(reg_file[1735]), .Y(n27440) );
  NOR2X1 U25803 ( .A(n25947), .B(n27398), .Y(n23392) );
  INVX1 U25804 ( .A(reg_file[1736]), .Y(n27398) );
  NOR2X1 U25805 ( .A(n25947), .B(n27356), .Y(n23391) );
  INVX1 U25806 ( .A(reg_file[1737]), .Y(n27356) );
  NOR2X1 U25807 ( .A(n25947), .B(n27314), .Y(n23390) );
  INVX1 U25808 ( .A(reg_file[1738]), .Y(n27314) );
  NOR2X1 U25809 ( .A(n25947), .B(n27272), .Y(n23389) );
  INVX1 U25810 ( .A(reg_file[1739]), .Y(n27272) );
  NOR2X1 U25811 ( .A(n25947), .B(n27230), .Y(n23388) );
  INVX1 U25812 ( .A(reg_file[1740]), .Y(n27230) );
  NOR2X1 U25813 ( .A(n25947), .B(n27188), .Y(n23387) );
  INVX1 U25814 ( .A(reg_file[1741]), .Y(n27188) );
  NOR2X1 U25815 ( .A(n25947), .B(n27146), .Y(n23386) );
  INVX1 U25816 ( .A(reg_file[1742]), .Y(n27146) );
  NOR2X1 U25817 ( .A(n25947), .B(n27104), .Y(n23385) );
  INVX1 U25818 ( .A(reg_file[1743]), .Y(n27104) );
  NOR2X1 U25819 ( .A(n25947), .B(n27020), .Y(n23384) );
  INVX1 U25820 ( .A(reg_file[1744]), .Y(n27020) );
  NOR2X1 U25821 ( .A(n25947), .B(n26978), .Y(n23383) );
  INVX1 U25822 ( .A(reg_file[1745]), .Y(n26978) );
  NOR2X1 U25823 ( .A(n25948), .B(n26936), .Y(n23382) );
  INVX1 U25824 ( .A(reg_file[1746]), .Y(n26936) );
  NOR2X1 U25825 ( .A(n25948), .B(n26894), .Y(n23381) );
  INVX1 U25826 ( .A(reg_file[1747]), .Y(n26894) );
  NOR2X1 U25827 ( .A(n25948), .B(n26852), .Y(n23380) );
  INVX1 U25828 ( .A(reg_file[1748]), .Y(n26852) );
  NOR2X1 U25829 ( .A(n25948), .B(n26810), .Y(n23379) );
  INVX1 U25830 ( .A(reg_file[1749]), .Y(n26810) );
  NOR2X1 U25831 ( .A(n25948), .B(n26768), .Y(n23378) );
  INVX1 U25832 ( .A(reg_file[1750]), .Y(n26768) );
  NOR2X1 U25833 ( .A(n25948), .B(n26726), .Y(n23377) );
  INVX1 U25834 ( .A(reg_file[1751]), .Y(n26726) );
  NOR2X1 U25835 ( .A(n25948), .B(n26684), .Y(n23376) );
  INVX1 U25836 ( .A(reg_file[1752]), .Y(n26684) );
  NOR2X1 U25837 ( .A(n25948), .B(n26642), .Y(n23375) );
  INVX1 U25838 ( .A(reg_file[1753]), .Y(n26642) );
  NOR2X1 U25839 ( .A(n25948), .B(n26558), .Y(n23374) );
  INVX1 U25840 ( .A(reg_file[1754]), .Y(n26558) );
  NOR2X1 U25841 ( .A(n25948), .B(n26516), .Y(n23373) );
  INVX1 U25842 ( .A(reg_file[1755]), .Y(n26516) );
  NOR2X1 U25843 ( .A(n25948), .B(n26474), .Y(n23372) );
  INVX1 U25844 ( .A(reg_file[1756]), .Y(n26474) );
  NOR2X1 U25845 ( .A(n25948), .B(n26432), .Y(n23371) );
  INVX1 U25846 ( .A(reg_file[1757]), .Y(n26432) );
  NOR2X1 U25847 ( .A(n25948), .B(n26390), .Y(n23370) );
  INVX1 U25848 ( .A(reg_file[1758]), .Y(n26390) );
  NOR2X1 U25849 ( .A(n25948), .B(n26348), .Y(n23369) );
  INVX1 U25850 ( .A(reg_file[1759]), .Y(n26348) );
  NOR2X1 U25851 ( .A(n25948), .B(n26306), .Y(n23368) );
  INVX1 U25852 ( .A(reg_file[1760]), .Y(n26306) );
  NOR2X1 U25853 ( .A(n25948), .B(n26264), .Y(n23367) );
  INVX1 U25854 ( .A(reg_file[1761]), .Y(n26264) );
  NOR2X1 U25855 ( .A(n25948), .B(n26222), .Y(n23366) );
  INVX1 U25856 ( .A(reg_file[1762]), .Y(n26222) );
  NOR2X1 U25857 ( .A(n25949), .B(n26180), .Y(n23365) );
  INVX1 U25858 ( .A(reg_file[1763]), .Y(n26180) );
  NOR2X1 U25859 ( .A(n25949), .B(n31430), .Y(n23364) );
  INVX1 U25860 ( .A(reg_file[1764]), .Y(n31430) );
  NOR2X1 U25861 ( .A(n25949), .B(n31388), .Y(n23363) );
  INVX1 U25862 ( .A(reg_file[1765]), .Y(n31388) );
  NOR2X1 U25863 ( .A(n25949), .B(n31346), .Y(n23362) );
  INVX1 U25864 ( .A(reg_file[1766]), .Y(n31346) );
  NOR2X1 U25865 ( .A(n25949), .B(n31304), .Y(n23361) );
  INVX1 U25866 ( .A(reg_file[1767]), .Y(n31304) );
  NOR2X1 U25867 ( .A(n25949), .B(n31262), .Y(n23360) );
  INVX1 U25868 ( .A(reg_file[1768]), .Y(n31262) );
  NOR2X1 U25869 ( .A(n25949), .B(n31220), .Y(n23359) );
  INVX1 U25870 ( .A(reg_file[1769]), .Y(n31220) );
  NOR2X1 U25871 ( .A(n25949), .B(n31178), .Y(n23358) );
  INVX1 U25872 ( .A(reg_file[1770]), .Y(n31178) );
  NOR2X1 U25873 ( .A(n25949), .B(n31136), .Y(n23357) );
  INVX1 U25874 ( .A(reg_file[1771]), .Y(n31136) );
  NOR2X1 U25875 ( .A(n25949), .B(n31094), .Y(n23356) );
  INVX1 U25876 ( .A(reg_file[1772]), .Y(n31094) );
  NOR2X1 U25877 ( .A(n25949), .B(n31052), .Y(n23355) );
  INVX1 U25878 ( .A(reg_file[1773]), .Y(n31052) );
  NOR2X1 U25879 ( .A(n25949), .B(n30968), .Y(n23354) );
  INVX1 U25880 ( .A(reg_file[1774]), .Y(n30968) );
  NOR2X1 U25881 ( .A(n25949), .B(n30926), .Y(n23353) );
  INVX1 U25882 ( .A(reg_file[1775]), .Y(n30926) );
  NOR2X1 U25883 ( .A(n25949), .B(n30884), .Y(n23352) );
  INVX1 U25884 ( .A(reg_file[1776]), .Y(n30884) );
  NOR2X1 U25885 ( .A(n25949), .B(n30842), .Y(n23351) );
  INVX1 U25886 ( .A(reg_file[1777]), .Y(n30842) );
  NOR2X1 U25887 ( .A(n25949), .B(n30800), .Y(n23350) );
  INVX1 U25888 ( .A(reg_file[1778]), .Y(n30800) );
  NOR2X1 U25889 ( .A(n25949), .B(n30758), .Y(n23349) );
  INVX1 U25890 ( .A(reg_file[1779]), .Y(n30758) );
  NOR2X1 U25891 ( .A(n25950), .B(n30716), .Y(n23348) );
  INVX1 U25892 ( .A(reg_file[1780]), .Y(n30716) );
  NOR2X1 U25893 ( .A(n25950), .B(n30674), .Y(n23347) );
  INVX1 U25894 ( .A(reg_file[1781]), .Y(n30674) );
  NOR2X1 U25895 ( .A(n25950), .B(n30632), .Y(n23346) );
  INVX1 U25896 ( .A(reg_file[1782]), .Y(n30632) );
  NOR2X1 U25897 ( .A(n25950), .B(n30590), .Y(n23345) );
  INVX1 U25898 ( .A(reg_file[1783]), .Y(n30590) );
  NOR2X1 U25899 ( .A(n25950), .B(n30506), .Y(n23344) );
  INVX1 U25900 ( .A(reg_file[1784]), .Y(n30506) );
  NOR2X1 U25901 ( .A(n25950), .B(n30464), .Y(n23343) );
  INVX1 U25902 ( .A(reg_file[1785]), .Y(n30464) );
  NOR2X1 U25903 ( .A(n25950), .B(n30422), .Y(n23342) );
  INVX1 U25904 ( .A(reg_file[1786]), .Y(n30422) );
  NOR2X1 U25905 ( .A(n25950), .B(n30380), .Y(n23341) );
  INVX1 U25906 ( .A(reg_file[1787]), .Y(n30380) );
  NOR2X1 U25907 ( .A(n25950), .B(n30338), .Y(n23340) );
  INVX1 U25908 ( .A(reg_file[1788]), .Y(n30338) );
  NOR2X1 U25909 ( .A(n25950), .B(n30296), .Y(n23339) );
  INVX1 U25910 ( .A(reg_file[1789]), .Y(n30296) );
  NOR2X1 U25911 ( .A(n25950), .B(n30254), .Y(n23338) );
  INVX1 U25912 ( .A(reg_file[1790]), .Y(n30254) );
  NOR2X1 U25913 ( .A(n25950), .B(n30212), .Y(n23337) );
  INVX1 U25914 ( .A(reg_file[1791]), .Y(n30212) );
  NOR2X1 U25915 ( .A(n35709), .B(n35058), .Y(n35969) );
  MUX2X1 U25916 ( .B(n31476), .A(n25129), .S(n25951), .Y(n23336) );
  INVX1 U25917 ( .A(reg_file[1792]), .Y(n31476) );
  MUX2X1 U25918 ( .B(n29835), .A(n25130), .S(n25951), .Y(n23335) );
  INVX1 U25919 ( .A(reg_file[1793]), .Y(n29835) );
  MUX2X1 U25920 ( .B(n29373), .A(n25131), .S(n25951), .Y(n23334) );
  INVX1 U25921 ( .A(reg_file[1794]), .Y(n29373) );
  MUX2X1 U25922 ( .B(n28911), .A(n25132), .S(n25951), .Y(n23333) );
  INVX1 U25923 ( .A(reg_file[1795]), .Y(n28911) );
  MUX2X1 U25924 ( .B(n28449), .A(n25133), .S(n25951), .Y(n23332) );
  INVX1 U25925 ( .A(reg_file[1796]), .Y(n28449) );
  MUX2X1 U25926 ( .B(n27987), .A(n25134), .S(n25951), .Y(n23331) );
  INVX1 U25927 ( .A(reg_file[1797]), .Y(n27987) );
  MUX2X1 U25928 ( .B(n27525), .A(n25135), .S(n25951), .Y(n23330) );
  INVX1 U25929 ( .A(reg_file[1798]), .Y(n27525) );
  MUX2X1 U25930 ( .B(n27063), .A(n25136), .S(n25951), .Y(n23329) );
  INVX1 U25931 ( .A(reg_file[1799]), .Y(n27063) );
  NOR2X1 U25932 ( .A(n25951), .B(n26601), .Y(n23328) );
  INVX1 U25933 ( .A(reg_file[1800]), .Y(n26601) );
  NOR2X1 U25934 ( .A(n25951), .B(n26110), .Y(n23327) );
  INVX1 U25935 ( .A(reg_file[1801]), .Y(n26110) );
  NOR2X1 U25936 ( .A(n25951), .B(n31011), .Y(n23326) );
  INVX1 U25937 ( .A(reg_file[1802]), .Y(n31011) );
  NOR2X1 U25938 ( .A(n25951), .B(n30549), .Y(n23325) );
  INVX1 U25939 ( .A(reg_file[1803]), .Y(n30549) );
  NOR2X1 U25940 ( .A(n25951), .B(n30171), .Y(n23324) );
  INVX1 U25941 ( .A(reg_file[1804]), .Y(n30171) );
  NOR2X1 U25942 ( .A(n25951), .B(n30129), .Y(n23323) );
  INVX1 U25943 ( .A(reg_file[1805]), .Y(n30129) );
  NOR2X1 U25944 ( .A(n25952), .B(n30087), .Y(n23322) );
  INVX1 U25945 ( .A(reg_file[1806]), .Y(n30087) );
  NOR2X1 U25946 ( .A(n25952), .B(n30045), .Y(n23321) );
  INVX1 U25947 ( .A(reg_file[1807]), .Y(n30045) );
  NOR2X1 U25948 ( .A(n25952), .B(n30003), .Y(n23320) );
  INVX1 U25949 ( .A(reg_file[1808]), .Y(n30003) );
  NOR2X1 U25950 ( .A(n25952), .B(n29961), .Y(n23319) );
  INVX1 U25951 ( .A(reg_file[1809]), .Y(n29961) );
  NOR2X1 U25952 ( .A(n25952), .B(n29919), .Y(n23318) );
  INVX1 U25953 ( .A(reg_file[1810]), .Y(n29919) );
  NOR2X1 U25954 ( .A(n25952), .B(n29877), .Y(n23317) );
  INVX1 U25955 ( .A(reg_file[1811]), .Y(n29877) );
  NOR2X1 U25956 ( .A(n25952), .B(n29793), .Y(n23316) );
  INVX1 U25957 ( .A(reg_file[1812]), .Y(n29793) );
  NOR2X1 U25958 ( .A(n25952), .B(n29751), .Y(n23315) );
  INVX1 U25959 ( .A(reg_file[1813]), .Y(n29751) );
  NOR2X1 U25960 ( .A(n25952), .B(n29709), .Y(n23314) );
  INVX1 U25961 ( .A(reg_file[1814]), .Y(n29709) );
  NOR2X1 U25962 ( .A(n25952), .B(n29667), .Y(n23313) );
  INVX1 U25963 ( .A(reg_file[1815]), .Y(n29667) );
  NOR2X1 U25964 ( .A(n25952), .B(n29625), .Y(n23312) );
  INVX1 U25965 ( .A(reg_file[1816]), .Y(n29625) );
  NOR2X1 U25966 ( .A(n25952), .B(n29583), .Y(n23311) );
  INVX1 U25967 ( .A(reg_file[1817]), .Y(n29583) );
  NOR2X1 U25968 ( .A(n25952), .B(n29541), .Y(n23310) );
  INVX1 U25969 ( .A(reg_file[1818]), .Y(n29541) );
  NOR2X1 U25970 ( .A(n25952), .B(n29499), .Y(n23309) );
  INVX1 U25971 ( .A(reg_file[1819]), .Y(n29499) );
  NOR2X1 U25972 ( .A(n25952), .B(n29457), .Y(n23308) );
  INVX1 U25973 ( .A(reg_file[1820]), .Y(n29457) );
  NOR2X1 U25974 ( .A(n25952), .B(n29415), .Y(n23307) );
  INVX1 U25975 ( .A(reg_file[1821]), .Y(n29415) );
  NOR2X1 U25976 ( .A(n25952), .B(n29331), .Y(n23306) );
  INVX1 U25977 ( .A(reg_file[1822]), .Y(n29331) );
  NOR2X1 U25978 ( .A(n25953), .B(n29289), .Y(n23305) );
  INVX1 U25979 ( .A(reg_file[1823]), .Y(n29289) );
  NOR2X1 U25980 ( .A(n25953), .B(n29247), .Y(n23304) );
  INVX1 U25981 ( .A(reg_file[1824]), .Y(n29247) );
  NOR2X1 U25982 ( .A(n25953), .B(n29205), .Y(n23303) );
  INVX1 U25983 ( .A(reg_file[1825]), .Y(n29205) );
  NOR2X1 U25984 ( .A(n25953), .B(n29163), .Y(n23302) );
  INVX1 U25985 ( .A(reg_file[1826]), .Y(n29163) );
  NOR2X1 U25986 ( .A(n25953), .B(n29121), .Y(n23301) );
  INVX1 U25987 ( .A(reg_file[1827]), .Y(n29121) );
  NOR2X1 U25988 ( .A(n25953), .B(n29079), .Y(n23300) );
  INVX1 U25989 ( .A(reg_file[1828]), .Y(n29079) );
  NOR2X1 U25990 ( .A(n25953), .B(n29037), .Y(n23299) );
  INVX1 U25991 ( .A(reg_file[1829]), .Y(n29037) );
  NOR2X1 U25992 ( .A(n25953), .B(n28995), .Y(n23298) );
  INVX1 U25993 ( .A(reg_file[1830]), .Y(n28995) );
  NOR2X1 U25994 ( .A(n25953), .B(n28953), .Y(n23297) );
  INVX1 U25995 ( .A(reg_file[1831]), .Y(n28953) );
  NOR2X1 U25996 ( .A(n25953), .B(n28869), .Y(n23296) );
  INVX1 U25997 ( .A(reg_file[1832]), .Y(n28869) );
  NOR2X1 U25998 ( .A(n25953), .B(n28827), .Y(n23295) );
  INVX1 U25999 ( .A(reg_file[1833]), .Y(n28827) );
  NOR2X1 U26000 ( .A(n25953), .B(n28785), .Y(n23294) );
  INVX1 U26001 ( .A(reg_file[1834]), .Y(n28785) );
  NOR2X1 U26002 ( .A(n25953), .B(n28743), .Y(n23293) );
  INVX1 U26003 ( .A(reg_file[1835]), .Y(n28743) );
  NOR2X1 U26004 ( .A(n25953), .B(n28701), .Y(n23292) );
  INVX1 U26005 ( .A(reg_file[1836]), .Y(n28701) );
  NOR2X1 U26006 ( .A(n25953), .B(n28659), .Y(n23291) );
  INVX1 U26007 ( .A(reg_file[1837]), .Y(n28659) );
  NOR2X1 U26008 ( .A(n25953), .B(n28617), .Y(n23290) );
  INVX1 U26009 ( .A(reg_file[1838]), .Y(n28617) );
  NOR2X1 U26010 ( .A(n25953), .B(n28575), .Y(n23289) );
  INVX1 U26011 ( .A(reg_file[1839]), .Y(n28575) );
  NOR2X1 U26012 ( .A(n25954), .B(n28533), .Y(n23288) );
  INVX1 U26013 ( .A(reg_file[1840]), .Y(n28533) );
  NOR2X1 U26014 ( .A(n25954), .B(n28491), .Y(n23287) );
  INVX1 U26015 ( .A(reg_file[1841]), .Y(n28491) );
  NOR2X1 U26016 ( .A(n25954), .B(n28407), .Y(n23286) );
  INVX1 U26017 ( .A(reg_file[1842]), .Y(n28407) );
  NOR2X1 U26018 ( .A(n25954), .B(n28365), .Y(n23285) );
  INVX1 U26019 ( .A(reg_file[1843]), .Y(n28365) );
  NOR2X1 U26020 ( .A(n25954), .B(n28323), .Y(n23284) );
  INVX1 U26021 ( .A(reg_file[1844]), .Y(n28323) );
  NOR2X1 U26022 ( .A(n25954), .B(n28281), .Y(n23283) );
  INVX1 U26023 ( .A(reg_file[1845]), .Y(n28281) );
  NOR2X1 U26024 ( .A(n25954), .B(n28239), .Y(n23282) );
  INVX1 U26025 ( .A(reg_file[1846]), .Y(n28239) );
  NOR2X1 U26026 ( .A(n25954), .B(n28197), .Y(n23281) );
  INVX1 U26027 ( .A(reg_file[1847]), .Y(n28197) );
  NOR2X1 U26028 ( .A(n25954), .B(n28155), .Y(n23280) );
  INVX1 U26029 ( .A(reg_file[1848]), .Y(n28155) );
  NOR2X1 U26030 ( .A(n25954), .B(n28113), .Y(n23279) );
  INVX1 U26031 ( .A(reg_file[1849]), .Y(n28113) );
  NOR2X1 U26032 ( .A(n25954), .B(n28071), .Y(n23278) );
  INVX1 U26033 ( .A(reg_file[1850]), .Y(n28071) );
  NOR2X1 U26034 ( .A(n25954), .B(n28029), .Y(n23277) );
  INVX1 U26035 ( .A(reg_file[1851]), .Y(n28029) );
  NOR2X1 U26036 ( .A(n25954), .B(n27945), .Y(n23276) );
  INVX1 U26037 ( .A(reg_file[1852]), .Y(n27945) );
  NOR2X1 U26038 ( .A(n25954), .B(n27903), .Y(n23275) );
  INVX1 U26039 ( .A(reg_file[1853]), .Y(n27903) );
  NOR2X1 U26040 ( .A(n25954), .B(n27861), .Y(n23274) );
  INVX1 U26041 ( .A(reg_file[1854]), .Y(n27861) );
  NOR2X1 U26042 ( .A(n25954), .B(n27819), .Y(n23273) );
  INVX1 U26043 ( .A(reg_file[1855]), .Y(n27819) );
  NOR2X1 U26044 ( .A(n25954), .B(n27777), .Y(n23272) );
  INVX1 U26045 ( .A(reg_file[1856]), .Y(n27777) );
  NOR2X1 U26046 ( .A(n25955), .B(n27735), .Y(n23271) );
  INVX1 U26047 ( .A(reg_file[1857]), .Y(n27735) );
  NOR2X1 U26048 ( .A(n25955), .B(n27693), .Y(n23270) );
  INVX1 U26049 ( .A(reg_file[1858]), .Y(n27693) );
  NOR2X1 U26050 ( .A(n25955), .B(n27651), .Y(n23269) );
  INVX1 U26051 ( .A(reg_file[1859]), .Y(n27651) );
  NOR2X1 U26052 ( .A(n25955), .B(n27609), .Y(n23268) );
  INVX1 U26053 ( .A(reg_file[1860]), .Y(n27609) );
  NOR2X1 U26054 ( .A(n25955), .B(n27567), .Y(n23267) );
  INVX1 U26055 ( .A(reg_file[1861]), .Y(n27567) );
  NOR2X1 U26056 ( .A(n25955), .B(n27483), .Y(n23266) );
  INVX1 U26057 ( .A(reg_file[1862]), .Y(n27483) );
  NOR2X1 U26058 ( .A(n25955), .B(n27441), .Y(n23265) );
  INVX1 U26059 ( .A(reg_file[1863]), .Y(n27441) );
  NOR2X1 U26060 ( .A(n25955), .B(n27399), .Y(n23264) );
  INVX1 U26061 ( .A(reg_file[1864]), .Y(n27399) );
  NOR2X1 U26062 ( .A(n25955), .B(n27357), .Y(n23263) );
  INVX1 U26063 ( .A(reg_file[1865]), .Y(n27357) );
  NOR2X1 U26064 ( .A(n25955), .B(n27315), .Y(n23262) );
  INVX1 U26065 ( .A(reg_file[1866]), .Y(n27315) );
  NOR2X1 U26066 ( .A(n25955), .B(n27273), .Y(n23261) );
  INVX1 U26067 ( .A(reg_file[1867]), .Y(n27273) );
  NOR2X1 U26068 ( .A(n25955), .B(n27231), .Y(n23260) );
  INVX1 U26069 ( .A(reg_file[1868]), .Y(n27231) );
  NOR2X1 U26070 ( .A(n25955), .B(n27189), .Y(n23259) );
  INVX1 U26071 ( .A(reg_file[1869]), .Y(n27189) );
  NOR2X1 U26072 ( .A(n25955), .B(n27147), .Y(n23258) );
  INVX1 U26073 ( .A(reg_file[1870]), .Y(n27147) );
  NOR2X1 U26074 ( .A(n25955), .B(n27105), .Y(n23257) );
  INVX1 U26075 ( .A(reg_file[1871]), .Y(n27105) );
  NOR2X1 U26076 ( .A(n25955), .B(n27021), .Y(n23256) );
  INVX1 U26077 ( .A(reg_file[1872]), .Y(n27021) );
  NOR2X1 U26078 ( .A(n25955), .B(n26979), .Y(n23255) );
  INVX1 U26079 ( .A(reg_file[1873]), .Y(n26979) );
  NOR2X1 U26080 ( .A(n25956), .B(n26937), .Y(n23254) );
  INVX1 U26081 ( .A(reg_file[1874]), .Y(n26937) );
  NOR2X1 U26082 ( .A(n25956), .B(n26895), .Y(n23253) );
  INVX1 U26083 ( .A(reg_file[1875]), .Y(n26895) );
  NOR2X1 U26084 ( .A(n25956), .B(n26853), .Y(n23252) );
  INVX1 U26085 ( .A(reg_file[1876]), .Y(n26853) );
  NOR2X1 U26086 ( .A(n25956), .B(n26811), .Y(n23251) );
  INVX1 U26087 ( .A(reg_file[1877]), .Y(n26811) );
  NOR2X1 U26088 ( .A(n25956), .B(n26769), .Y(n23250) );
  INVX1 U26089 ( .A(reg_file[1878]), .Y(n26769) );
  NOR2X1 U26090 ( .A(n25956), .B(n26727), .Y(n23249) );
  INVX1 U26091 ( .A(reg_file[1879]), .Y(n26727) );
  NOR2X1 U26092 ( .A(n25956), .B(n26685), .Y(n23248) );
  INVX1 U26093 ( .A(reg_file[1880]), .Y(n26685) );
  NOR2X1 U26094 ( .A(n25956), .B(n26643), .Y(n23247) );
  INVX1 U26095 ( .A(reg_file[1881]), .Y(n26643) );
  NOR2X1 U26096 ( .A(n25956), .B(n26559), .Y(n23246) );
  INVX1 U26097 ( .A(reg_file[1882]), .Y(n26559) );
  NOR2X1 U26098 ( .A(n25956), .B(n26517), .Y(n23245) );
  INVX1 U26099 ( .A(reg_file[1883]), .Y(n26517) );
  NOR2X1 U26100 ( .A(n25956), .B(n26475), .Y(n23244) );
  INVX1 U26101 ( .A(reg_file[1884]), .Y(n26475) );
  NOR2X1 U26102 ( .A(n25956), .B(n26433), .Y(n23243) );
  INVX1 U26103 ( .A(reg_file[1885]), .Y(n26433) );
  NOR2X1 U26104 ( .A(n25956), .B(n26391), .Y(n23242) );
  INVX1 U26105 ( .A(reg_file[1886]), .Y(n26391) );
  NOR2X1 U26106 ( .A(n25956), .B(n26349), .Y(n23241) );
  INVX1 U26107 ( .A(reg_file[1887]), .Y(n26349) );
  NOR2X1 U26108 ( .A(n25956), .B(n26307), .Y(n23240) );
  INVX1 U26109 ( .A(reg_file[1888]), .Y(n26307) );
  NOR2X1 U26110 ( .A(n25956), .B(n26265), .Y(n23239) );
  INVX1 U26111 ( .A(reg_file[1889]), .Y(n26265) );
  NOR2X1 U26112 ( .A(n25956), .B(n26223), .Y(n23238) );
  INVX1 U26113 ( .A(reg_file[1890]), .Y(n26223) );
  NOR2X1 U26114 ( .A(n25957), .B(n26181), .Y(n23237) );
  INVX1 U26115 ( .A(reg_file[1891]), .Y(n26181) );
  NOR2X1 U26116 ( .A(n25957), .B(n31431), .Y(n23236) );
  INVX1 U26117 ( .A(reg_file[1892]), .Y(n31431) );
  NOR2X1 U26118 ( .A(n25957), .B(n31389), .Y(n23235) );
  INVX1 U26119 ( .A(reg_file[1893]), .Y(n31389) );
  NOR2X1 U26120 ( .A(n25957), .B(n31347), .Y(n23234) );
  INVX1 U26121 ( .A(reg_file[1894]), .Y(n31347) );
  NOR2X1 U26122 ( .A(n25957), .B(n31305), .Y(n23233) );
  INVX1 U26123 ( .A(reg_file[1895]), .Y(n31305) );
  NOR2X1 U26124 ( .A(n25957), .B(n31263), .Y(n23232) );
  INVX1 U26125 ( .A(reg_file[1896]), .Y(n31263) );
  NOR2X1 U26126 ( .A(n25957), .B(n31221), .Y(n23231) );
  INVX1 U26127 ( .A(reg_file[1897]), .Y(n31221) );
  NOR2X1 U26128 ( .A(n25957), .B(n31179), .Y(n23230) );
  INVX1 U26129 ( .A(reg_file[1898]), .Y(n31179) );
  NOR2X1 U26130 ( .A(n25957), .B(n31137), .Y(n23229) );
  INVX1 U26131 ( .A(reg_file[1899]), .Y(n31137) );
  NOR2X1 U26132 ( .A(n25957), .B(n31095), .Y(n23228) );
  INVX1 U26133 ( .A(reg_file[1900]), .Y(n31095) );
  NOR2X1 U26134 ( .A(n25957), .B(n31053), .Y(n23227) );
  INVX1 U26135 ( .A(reg_file[1901]), .Y(n31053) );
  NOR2X1 U26136 ( .A(n25957), .B(n30969), .Y(n23226) );
  INVX1 U26137 ( .A(reg_file[1902]), .Y(n30969) );
  NOR2X1 U26138 ( .A(n25957), .B(n30927), .Y(n23225) );
  INVX1 U26139 ( .A(reg_file[1903]), .Y(n30927) );
  NOR2X1 U26140 ( .A(n25957), .B(n30885), .Y(n23224) );
  INVX1 U26141 ( .A(reg_file[1904]), .Y(n30885) );
  NOR2X1 U26142 ( .A(n25957), .B(n30843), .Y(n23223) );
  INVX1 U26143 ( .A(reg_file[1905]), .Y(n30843) );
  NOR2X1 U26144 ( .A(n25957), .B(n30801), .Y(n23222) );
  INVX1 U26145 ( .A(reg_file[1906]), .Y(n30801) );
  NOR2X1 U26146 ( .A(n25957), .B(n30759), .Y(n23221) );
  INVX1 U26147 ( .A(reg_file[1907]), .Y(n30759) );
  NOR2X1 U26148 ( .A(n25958), .B(n30717), .Y(n23220) );
  INVX1 U26149 ( .A(reg_file[1908]), .Y(n30717) );
  NOR2X1 U26150 ( .A(n25958), .B(n30675), .Y(n23219) );
  INVX1 U26151 ( .A(reg_file[1909]), .Y(n30675) );
  NOR2X1 U26152 ( .A(n25958), .B(n30633), .Y(n23218) );
  INVX1 U26153 ( .A(reg_file[1910]), .Y(n30633) );
  NOR2X1 U26154 ( .A(n25958), .B(n30591), .Y(n23217) );
  INVX1 U26155 ( .A(reg_file[1911]), .Y(n30591) );
  NOR2X1 U26156 ( .A(n25958), .B(n30507), .Y(n23216) );
  INVX1 U26157 ( .A(reg_file[1912]), .Y(n30507) );
  NOR2X1 U26158 ( .A(n25958), .B(n30465), .Y(n23215) );
  INVX1 U26159 ( .A(reg_file[1913]), .Y(n30465) );
  NOR2X1 U26160 ( .A(n25958), .B(n30423), .Y(n23214) );
  INVX1 U26161 ( .A(reg_file[1914]), .Y(n30423) );
  NOR2X1 U26162 ( .A(n25958), .B(n30381), .Y(n23213) );
  INVX1 U26163 ( .A(reg_file[1915]), .Y(n30381) );
  NOR2X1 U26164 ( .A(n25958), .B(n30339), .Y(n23212) );
  INVX1 U26165 ( .A(reg_file[1916]), .Y(n30339) );
  NOR2X1 U26166 ( .A(n25958), .B(n30297), .Y(n23211) );
  INVX1 U26167 ( .A(reg_file[1917]), .Y(n30297) );
  NOR2X1 U26168 ( .A(n25958), .B(n30255), .Y(n23210) );
  INVX1 U26169 ( .A(reg_file[1918]), .Y(n30255) );
  NOR2X1 U26170 ( .A(n25958), .B(n30213), .Y(n23209) );
  INVX1 U26171 ( .A(reg_file[1919]), .Y(n30213) );
  NOR2X1 U26172 ( .A(n35579), .B(n35317), .Y(n35970) );
  NAND3X1 U26173 ( .A(n35320), .B(n35319), .C(wraddr[3]), .Y(n35579) );
  MUX2X1 U26174 ( .B(n31477), .A(n25129), .S(n25959), .Y(n23208) );
  INVX1 U26175 ( .A(reg_file[1920]), .Y(n31477) );
  MUX2X1 U26176 ( .B(n29836), .A(n25130), .S(n25959), .Y(n23207) );
  INVX1 U26177 ( .A(reg_file[1921]), .Y(n29836) );
  MUX2X1 U26178 ( .B(n29374), .A(n25131), .S(n25959), .Y(n23206) );
  INVX1 U26179 ( .A(reg_file[1922]), .Y(n29374) );
  MUX2X1 U26180 ( .B(n28912), .A(n25132), .S(n25959), .Y(n23205) );
  INVX1 U26181 ( .A(reg_file[1923]), .Y(n28912) );
  MUX2X1 U26182 ( .B(n28450), .A(n25133), .S(n25959), .Y(n23204) );
  INVX1 U26183 ( .A(reg_file[1924]), .Y(n28450) );
  MUX2X1 U26184 ( .B(n27988), .A(n25134), .S(n25959), .Y(n23203) );
  INVX1 U26185 ( .A(reg_file[1925]), .Y(n27988) );
  MUX2X1 U26186 ( .B(n27526), .A(n25135), .S(n25959), .Y(n23202) );
  INVX1 U26187 ( .A(reg_file[1926]), .Y(n27526) );
  MUX2X1 U26188 ( .B(n27064), .A(n25136), .S(n25959), .Y(n23201) );
  INVX1 U26189 ( .A(reg_file[1927]), .Y(n27064) );
  NOR2X1 U26190 ( .A(n25959), .B(n26602), .Y(n23200) );
  INVX1 U26191 ( .A(reg_file[1928]), .Y(n26602) );
  NOR2X1 U26192 ( .A(n25959), .B(n26112), .Y(n23199) );
  INVX1 U26193 ( .A(reg_file[1929]), .Y(n26112) );
  NOR2X1 U26194 ( .A(n25959), .B(n31012), .Y(n23198) );
  INVX1 U26195 ( .A(reg_file[1930]), .Y(n31012) );
  NOR2X1 U26196 ( .A(n25959), .B(n30550), .Y(n23197) );
  INVX1 U26197 ( .A(reg_file[1931]), .Y(n30550) );
  NOR2X1 U26198 ( .A(n25959), .B(n30172), .Y(n23196) );
  INVX1 U26199 ( .A(reg_file[1932]), .Y(n30172) );
  NOR2X1 U26200 ( .A(n25959), .B(n30130), .Y(n23195) );
  INVX1 U26201 ( .A(reg_file[1933]), .Y(n30130) );
  NOR2X1 U26202 ( .A(n25960), .B(n30088), .Y(n23194) );
  INVX1 U26203 ( .A(reg_file[1934]), .Y(n30088) );
  NOR2X1 U26204 ( .A(n25960), .B(n30046), .Y(n23193) );
  INVX1 U26205 ( .A(reg_file[1935]), .Y(n30046) );
  NOR2X1 U26206 ( .A(n25960), .B(n30004), .Y(n23192) );
  INVX1 U26207 ( .A(reg_file[1936]), .Y(n30004) );
  NOR2X1 U26208 ( .A(n25960), .B(n29962), .Y(n23191) );
  INVX1 U26209 ( .A(reg_file[1937]), .Y(n29962) );
  NOR2X1 U26210 ( .A(n25960), .B(n29920), .Y(n23190) );
  INVX1 U26211 ( .A(reg_file[1938]), .Y(n29920) );
  NOR2X1 U26212 ( .A(n25960), .B(n29878), .Y(n23189) );
  INVX1 U26213 ( .A(reg_file[1939]), .Y(n29878) );
  NOR2X1 U26214 ( .A(n25960), .B(n29794), .Y(n23188) );
  INVX1 U26215 ( .A(reg_file[1940]), .Y(n29794) );
  NOR2X1 U26216 ( .A(n25960), .B(n29752), .Y(n23187) );
  INVX1 U26217 ( .A(reg_file[1941]), .Y(n29752) );
  NOR2X1 U26218 ( .A(n25960), .B(n29710), .Y(n23186) );
  INVX1 U26219 ( .A(reg_file[1942]), .Y(n29710) );
  NOR2X1 U26220 ( .A(n25960), .B(n29668), .Y(n23185) );
  INVX1 U26221 ( .A(reg_file[1943]), .Y(n29668) );
  NOR2X1 U26222 ( .A(n25960), .B(n29626), .Y(n23184) );
  INVX1 U26223 ( .A(reg_file[1944]), .Y(n29626) );
  NOR2X1 U26224 ( .A(n25960), .B(n29584), .Y(n23183) );
  INVX1 U26225 ( .A(reg_file[1945]), .Y(n29584) );
  NOR2X1 U26226 ( .A(n25960), .B(n29542), .Y(n23182) );
  INVX1 U26227 ( .A(reg_file[1946]), .Y(n29542) );
  NOR2X1 U26228 ( .A(n25960), .B(n29500), .Y(n23181) );
  INVX1 U26229 ( .A(reg_file[1947]), .Y(n29500) );
  NOR2X1 U26230 ( .A(n25960), .B(n29458), .Y(n23180) );
  INVX1 U26231 ( .A(reg_file[1948]), .Y(n29458) );
  NOR2X1 U26232 ( .A(n25960), .B(n29416), .Y(n23179) );
  INVX1 U26233 ( .A(reg_file[1949]), .Y(n29416) );
  NOR2X1 U26234 ( .A(n25960), .B(n29332), .Y(n23178) );
  INVX1 U26235 ( .A(reg_file[1950]), .Y(n29332) );
  NOR2X1 U26236 ( .A(n25961), .B(n29290), .Y(n23177) );
  INVX1 U26237 ( .A(reg_file[1951]), .Y(n29290) );
  NOR2X1 U26238 ( .A(n25961), .B(n29248), .Y(n23176) );
  INVX1 U26239 ( .A(reg_file[1952]), .Y(n29248) );
  NOR2X1 U26240 ( .A(n25961), .B(n29206), .Y(n23175) );
  INVX1 U26241 ( .A(reg_file[1953]), .Y(n29206) );
  NOR2X1 U26242 ( .A(n25961), .B(n29164), .Y(n23174) );
  INVX1 U26243 ( .A(reg_file[1954]), .Y(n29164) );
  NOR2X1 U26244 ( .A(n25961), .B(n29122), .Y(n23173) );
  INVX1 U26245 ( .A(reg_file[1955]), .Y(n29122) );
  NOR2X1 U26246 ( .A(n25961), .B(n29080), .Y(n23172) );
  INVX1 U26247 ( .A(reg_file[1956]), .Y(n29080) );
  NOR2X1 U26248 ( .A(n25961), .B(n29038), .Y(n23171) );
  INVX1 U26249 ( .A(reg_file[1957]), .Y(n29038) );
  NOR2X1 U26250 ( .A(n25961), .B(n28996), .Y(n23170) );
  INVX1 U26251 ( .A(reg_file[1958]), .Y(n28996) );
  NOR2X1 U26252 ( .A(n25961), .B(n28954), .Y(n23169) );
  INVX1 U26253 ( .A(reg_file[1959]), .Y(n28954) );
  NOR2X1 U26254 ( .A(n25961), .B(n28870), .Y(n23168) );
  INVX1 U26255 ( .A(reg_file[1960]), .Y(n28870) );
  NOR2X1 U26256 ( .A(n25961), .B(n28828), .Y(n23167) );
  INVX1 U26257 ( .A(reg_file[1961]), .Y(n28828) );
  NOR2X1 U26258 ( .A(n25961), .B(n28786), .Y(n23166) );
  INVX1 U26259 ( .A(reg_file[1962]), .Y(n28786) );
  NOR2X1 U26260 ( .A(n25961), .B(n28744), .Y(n23165) );
  INVX1 U26261 ( .A(reg_file[1963]), .Y(n28744) );
  NOR2X1 U26262 ( .A(n25961), .B(n28702), .Y(n23164) );
  INVX1 U26263 ( .A(reg_file[1964]), .Y(n28702) );
  NOR2X1 U26264 ( .A(n25961), .B(n28660), .Y(n23163) );
  INVX1 U26265 ( .A(reg_file[1965]), .Y(n28660) );
  NOR2X1 U26266 ( .A(n25961), .B(n28618), .Y(n23162) );
  INVX1 U26267 ( .A(reg_file[1966]), .Y(n28618) );
  NOR2X1 U26268 ( .A(n25961), .B(n28576), .Y(n23161) );
  INVX1 U26269 ( .A(reg_file[1967]), .Y(n28576) );
  NOR2X1 U26270 ( .A(n25962), .B(n28534), .Y(n23160) );
  INVX1 U26271 ( .A(reg_file[1968]), .Y(n28534) );
  NOR2X1 U26272 ( .A(n25962), .B(n28492), .Y(n23159) );
  INVX1 U26273 ( .A(reg_file[1969]), .Y(n28492) );
  NOR2X1 U26274 ( .A(n25962), .B(n28408), .Y(n23158) );
  INVX1 U26275 ( .A(reg_file[1970]), .Y(n28408) );
  NOR2X1 U26276 ( .A(n25962), .B(n28366), .Y(n23157) );
  INVX1 U26277 ( .A(reg_file[1971]), .Y(n28366) );
  NOR2X1 U26278 ( .A(n25962), .B(n28324), .Y(n23156) );
  INVX1 U26279 ( .A(reg_file[1972]), .Y(n28324) );
  NOR2X1 U26280 ( .A(n25962), .B(n28282), .Y(n23155) );
  INVX1 U26281 ( .A(reg_file[1973]), .Y(n28282) );
  NOR2X1 U26282 ( .A(n25962), .B(n28240), .Y(n23154) );
  INVX1 U26283 ( .A(reg_file[1974]), .Y(n28240) );
  NOR2X1 U26284 ( .A(n25962), .B(n28198), .Y(n23153) );
  INVX1 U26285 ( .A(reg_file[1975]), .Y(n28198) );
  NOR2X1 U26286 ( .A(n25962), .B(n28156), .Y(n23152) );
  INVX1 U26287 ( .A(reg_file[1976]), .Y(n28156) );
  NOR2X1 U26288 ( .A(n25962), .B(n28114), .Y(n23151) );
  INVX1 U26289 ( .A(reg_file[1977]), .Y(n28114) );
  NOR2X1 U26290 ( .A(n25962), .B(n28072), .Y(n23150) );
  INVX1 U26291 ( .A(reg_file[1978]), .Y(n28072) );
  NOR2X1 U26292 ( .A(n25962), .B(n28030), .Y(n23149) );
  INVX1 U26293 ( .A(reg_file[1979]), .Y(n28030) );
  NOR2X1 U26294 ( .A(n25962), .B(n27946), .Y(n23148) );
  INVX1 U26295 ( .A(reg_file[1980]), .Y(n27946) );
  NOR2X1 U26296 ( .A(n25962), .B(n27904), .Y(n23147) );
  INVX1 U26297 ( .A(reg_file[1981]), .Y(n27904) );
  NOR2X1 U26298 ( .A(n25962), .B(n27862), .Y(n23146) );
  INVX1 U26299 ( .A(reg_file[1982]), .Y(n27862) );
  NOR2X1 U26300 ( .A(n25962), .B(n27820), .Y(n23145) );
  INVX1 U26301 ( .A(reg_file[1983]), .Y(n27820) );
  NOR2X1 U26302 ( .A(n25962), .B(n27778), .Y(n23144) );
  INVX1 U26303 ( .A(reg_file[1984]), .Y(n27778) );
  NOR2X1 U26304 ( .A(n25963), .B(n27736), .Y(n23143) );
  INVX1 U26305 ( .A(reg_file[1985]), .Y(n27736) );
  NOR2X1 U26306 ( .A(n25963), .B(n27694), .Y(n23142) );
  INVX1 U26307 ( .A(reg_file[1986]), .Y(n27694) );
  NOR2X1 U26308 ( .A(n25963), .B(n27652), .Y(n23141) );
  INVX1 U26309 ( .A(reg_file[1987]), .Y(n27652) );
  NOR2X1 U26310 ( .A(n25963), .B(n27610), .Y(n23140) );
  INVX1 U26311 ( .A(reg_file[1988]), .Y(n27610) );
  NOR2X1 U26312 ( .A(n25963), .B(n27568), .Y(n23139) );
  INVX1 U26313 ( .A(reg_file[1989]), .Y(n27568) );
  NOR2X1 U26314 ( .A(n25963), .B(n27484), .Y(n23138) );
  INVX1 U26315 ( .A(reg_file[1990]), .Y(n27484) );
  NOR2X1 U26316 ( .A(n25963), .B(n27442), .Y(n23137) );
  INVX1 U26317 ( .A(reg_file[1991]), .Y(n27442) );
  NOR2X1 U26318 ( .A(n25963), .B(n27400), .Y(n23136) );
  INVX1 U26319 ( .A(reg_file[1992]), .Y(n27400) );
  NOR2X1 U26320 ( .A(n25963), .B(n27358), .Y(n23135) );
  INVX1 U26321 ( .A(reg_file[1993]), .Y(n27358) );
  NOR2X1 U26322 ( .A(n25963), .B(n27316), .Y(n23134) );
  INVX1 U26323 ( .A(reg_file[1994]), .Y(n27316) );
  NOR2X1 U26324 ( .A(n25963), .B(n27274), .Y(n23133) );
  INVX1 U26325 ( .A(reg_file[1995]), .Y(n27274) );
  NOR2X1 U26326 ( .A(n25963), .B(n27232), .Y(n23132) );
  INVX1 U26327 ( .A(reg_file[1996]), .Y(n27232) );
  NOR2X1 U26328 ( .A(n25963), .B(n27190), .Y(n23131) );
  INVX1 U26329 ( .A(reg_file[1997]), .Y(n27190) );
  NOR2X1 U26330 ( .A(n25963), .B(n27148), .Y(n23130) );
  INVX1 U26331 ( .A(reg_file[1998]), .Y(n27148) );
  NOR2X1 U26332 ( .A(n25963), .B(n27106), .Y(n23129) );
  INVX1 U26333 ( .A(reg_file[1999]), .Y(n27106) );
  NOR2X1 U26334 ( .A(n25963), .B(n27022), .Y(n23128) );
  INVX1 U26335 ( .A(reg_file[2000]), .Y(n27022) );
  NOR2X1 U26336 ( .A(n25963), .B(n26980), .Y(n23127) );
  INVX1 U26337 ( .A(reg_file[2001]), .Y(n26980) );
  NOR2X1 U26338 ( .A(n25964), .B(n26938), .Y(n23126) );
  INVX1 U26339 ( .A(reg_file[2002]), .Y(n26938) );
  NOR2X1 U26340 ( .A(n25964), .B(n26896), .Y(n23125) );
  INVX1 U26341 ( .A(reg_file[2003]), .Y(n26896) );
  NOR2X1 U26342 ( .A(n25964), .B(n26854), .Y(n23124) );
  INVX1 U26343 ( .A(reg_file[2004]), .Y(n26854) );
  NOR2X1 U26344 ( .A(n25964), .B(n26812), .Y(n23123) );
  INVX1 U26345 ( .A(reg_file[2005]), .Y(n26812) );
  NOR2X1 U26346 ( .A(n25964), .B(n26770), .Y(n23122) );
  INVX1 U26347 ( .A(reg_file[2006]), .Y(n26770) );
  NOR2X1 U26348 ( .A(n25964), .B(n26728), .Y(n23121) );
  INVX1 U26349 ( .A(reg_file[2007]), .Y(n26728) );
  NOR2X1 U26350 ( .A(n25964), .B(n26686), .Y(n23120) );
  INVX1 U26351 ( .A(reg_file[2008]), .Y(n26686) );
  NOR2X1 U26352 ( .A(n25964), .B(n26644), .Y(n23119) );
  INVX1 U26353 ( .A(reg_file[2009]), .Y(n26644) );
  NOR2X1 U26354 ( .A(n25964), .B(n26560), .Y(n23118) );
  INVX1 U26355 ( .A(reg_file[2010]), .Y(n26560) );
  NOR2X1 U26356 ( .A(n25964), .B(n26518), .Y(n23117) );
  INVX1 U26357 ( .A(reg_file[2011]), .Y(n26518) );
  NOR2X1 U26358 ( .A(n25964), .B(n26476), .Y(n23116) );
  INVX1 U26359 ( .A(reg_file[2012]), .Y(n26476) );
  NOR2X1 U26360 ( .A(n25964), .B(n26434), .Y(n23115) );
  INVX1 U26361 ( .A(reg_file[2013]), .Y(n26434) );
  NOR2X1 U26362 ( .A(n25964), .B(n26392), .Y(n23114) );
  INVX1 U26363 ( .A(reg_file[2014]), .Y(n26392) );
  NOR2X1 U26364 ( .A(n25964), .B(n26350), .Y(n23113) );
  INVX1 U26365 ( .A(reg_file[2015]), .Y(n26350) );
  NOR2X1 U26366 ( .A(n25964), .B(n26308), .Y(n23112) );
  INVX1 U26367 ( .A(reg_file[2016]), .Y(n26308) );
  NOR2X1 U26368 ( .A(n25964), .B(n26266), .Y(n23111) );
  INVX1 U26369 ( .A(reg_file[2017]), .Y(n26266) );
  NOR2X1 U26370 ( .A(n25964), .B(n26224), .Y(n23110) );
  INVX1 U26371 ( .A(reg_file[2018]), .Y(n26224) );
  NOR2X1 U26372 ( .A(n25965), .B(n26182), .Y(n23109) );
  INVX1 U26373 ( .A(reg_file[2019]), .Y(n26182) );
  NOR2X1 U26374 ( .A(n25965), .B(n31432), .Y(n23108) );
  INVX1 U26375 ( .A(reg_file[2020]), .Y(n31432) );
  NOR2X1 U26376 ( .A(n25965), .B(n31390), .Y(n23107) );
  INVX1 U26377 ( .A(reg_file[2021]), .Y(n31390) );
  NOR2X1 U26378 ( .A(n25965), .B(n31348), .Y(n23106) );
  INVX1 U26379 ( .A(reg_file[2022]), .Y(n31348) );
  NOR2X1 U26380 ( .A(n25965), .B(n31306), .Y(n23105) );
  INVX1 U26381 ( .A(reg_file[2023]), .Y(n31306) );
  NOR2X1 U26382 ( .A(n25965), .B(n31264), .Y(n23104) );
  INVX1 U26383 ( .A(reg_file[2024]), .Y(n31264) );
  NOR2X1 U26384 ( .A(n25965), .B(n31222), .Y(n23103) );
  INVX1 U26385 ( .A(reg_file[2025]), .Y(n31222) );
  NOR2X1 U26386 ( .A(n25965), .B(n31180), .Y(n23102) );
  INVX1 U26387 ( .A(reg_file[2026]), .Y(n31180) );
  NOR2X1 U26388 ( .A(n25965), .B(n31138), .Y(n23101) );
  INVX1 U26389 ( .A(reg_file[2027]), .Y(n31138) );
  NOR2X1 U26390 ( .A(n25965), .B(n31096), .Y(n23100) );
  INVX1 U26391 ( .A(reg_file[2028]), .Y(n31096) );
  NOR2X1 U26392 ( .A(n25965), .B(n31054), .Y(n23099) );
  INVX1 U26393 ( .A(reg_file[2029]), .Y(n31054) );
  NOR2X1 U26394 ( .A(n25965), .B(n30970), .Y(n23098) );
  INVX1 U26395 ( .A(reg_file[2030]), .Y(n30970) );
  NOR2X1 U26396 ( .A(n25965), .B(n30928), .Y(n23097) );
  INVX1 U26397 ( .A(reg_file[2031]), .Y(n30928) );
  NOR2X1 U26398 ( .A(n25965), .B(n30886), .Y(n23096) );
  INVX1 U26399 ( .A(reg_file[2032]), .Y(n30886) );
  NOR2X1 U26400 ( .A(n25965), .B(n30844), .Y(n23095) );
  INVX1 U26401 ( .A(reg_file[2033]), .Y(n30844) );
  NOR2X1 U26402 ( .A(n25965), .B(n30802), .Y(n23094) );
  INVX1 U26403 ( .A(reg_file[2034]), .Y(n30802) );
  NOR2X1 U26404 ( .A(n25965), .B(n30760), .Y(n23093) );
  INVX1 U26405 ( .A(reg_file[2035]), .Y(n30760) );
  NOR2X1 U26406 ( .A(n25966), .B(n30718), .Y(n23092) );
  INVX1 U26407 ( .A(reg_file[2036]), .Y(n30718) );
  NOR2X1 U26408 ( .A(n25966), .B(n30676), .Y(n23091) );
  INVX1 U26409 ( .A(reg_file[2037]), .Y(n30676) );
  NOR2X1 U26410 ( .A(n25966), .B(n30634), .Y(n23090) );
  INVX1 U26411 ( .A(reg_file[2038]), .Y(n30634) );
  NOR2X1 U26412 ( .A(n25966), .B(n30592), .Y(n23089) );
  INVX1 U26413 ( .A(reg_file[2039]), .Y(n30592) );
  NOR2X1 U26414 ( .A(n25966), .B(n30508), .Y(n23088) );
  INVX1 U26415 ( .A(reg_file[2040]), .Y(n30508) );
  NOR2X1 U26416 ( .A(n25966), .B(n30466), .Y(n23087) );
  INVX1 U26417 ( .A(reg_file[2041]), .Y(n30466) );
  NOR2X1 U26418 ( .A(n25966), .B(n30424), .Y(n23086) );
  INVX1 U26419 ( .A(reg_file[2042]), .Y(n30424) );
  NOR2X1 U26420 ( .A(n25966), .B(n30382), .Y(n23085) );
  INVX1 U26421 ( .A(reg_file[2043]), .Y(n30382) );
  NOR2X1 U26422 ( .A(n25966), .B(n30340), .Y(n23084) );
  INVX1 U26423 ( .A(reg_file[2044]), .Y(n30340) );
  NOR2X1 U26424 ( .A(n25966), .B(n30298), .Y(n23083) );
  INVX1 U26425 ( .A(reg_file[2045]), .Y(n30298) );
  NOR2X1 U26426 ( .A(n25966), .B(n30256), .Y(n23082) );
  INVX1 U26427 ( .A(reg_file[2046]), .Y(n30256) );
  NOR2X1 U26428 ( .A(n25966), .B(n30214), .Y(n23081) );
  INVX1 U26429 ( .A(reg_file[2047]), .Y(n30214) );
  NOR2X1 U26430 ( .A(n35709), .B(n35317), .Y(n35971) );
  NAND3X1 U26431 ( .A(wraddr[0]), .B(n35319), .C(wraddr[3]), .Y(n35709) );
  INVX1 U26432 ( .A(wraddr[4]), .Y(n35319) );
  MUX2X1 U26433 ( .B(n35972), .A(n25129), .S(n25967), .Y(n23080) );
  INVX1 U26434 ( .A(reg_file[2048]), .Y(n35972) );
  MUX2X1 U26435 ( .B(n35974), .A(n25130), .S(n25967), .Y(n23079) );
  INVX1 U26436 ( .A(reg_file[2049]), .Y(n35974) );
  MUX2X1 U26437 ( .B(n35975), .A(n25131), .S(n25967), .Y(n23078) );
  INVX1 U26438 ( .A(reg_file[2050]), .Y(n35975) );
  MUX2X1 U26439 ( .B(n35976), .A(n25132), .S(n25967), .Y(n23077) );
  INVX1 U26440 ( .A(reg_file[2051]), .Y(n35976) );
  MUX2X1 U26441 ( .B(n35977), .A(n25133), .S(n25967), .Y(n23076) );
  INVX1 U26442 ( .A(reg_file[2052]), .Y(n35977) );
  MUX2X1 U26443 ( .B(n35978), .A(n25134), .S(n25967), .Y(n23075) );
  INVX1 U26444 ( .A(reg_file[2053]), .Y(n35978) );
  MUX2X1 U26445 ( .B(n35979), .A(n25135), .S(n25967), .Y(n23074) );
  INVX1 U26446 ( .A(reg_file[2054]), .Y(n35979) );
  MUX2X1 U26447 ( .B(n35980), .A(n25136), .S(n25967), .Y(n23073) );
  INVX1 U26448 ( .A(reg_file[2055]), .Y(n35980) );
  NOR2X1 U26449 ( .A(n25967), .B(n35981), .Y(n23072) );
  INVX1 U26450 ( .A(reg_file[2056]), .Y(n35981) );
  NOR2X1 U26451 ( .A(n25967), .B(n35982), .Y(n23071) );
  INVX1 U26452 ( .A(reg_file[2057]), .Y(n35982) );
  NOR2X1 U26453 ( .A(n25967), .B(n35983), .Y(n23070) );
  INVX1 U26454 ( .A(reg_file[2058]), .Y(n35983) );
  NOR2X1 U26455 ( .A(n25967), .B(n35984), .Y(n23069) );
  INVX1 U26456 ( .A(reg_file[2059]), .Y(n35984) );
  NOR2X1 U26457 ( .A(n25967), .B(n35985), .Y(n23068) );
  INVX1 U26458 ( .A(reg_file[2060]), .Y(n35985) );
  NOR2X1 U26459 ( .A(n25967), .B(n35986), .Y(n23067) );
  INVX1 U26460 ( .A(reg_file[2061]), .Y(n35986) );
  NOR2X1 U26461 ( .A(n25968), .B(n35987), .Y(n23066) );
  INVX1 U26462 ( .A(reg_file[2062]), .Y(n35987) );
  NOR2X1 U26463 ( .A(n25968), .B(n35988), .Y(n23065) );
  INVX1 U26464 ( .A(reg_file[2063]), .Y(n35988) );
  NOR2X1 U26465 ( .A(n25968), .B(n35989), .Y(n23064) );
  INVX1 U26466 ( .A(reg_file[2064]), .Y(n35989) );
  NOR2X1 U26467 ( .A(n25968), .B(n35990), .Y(n23063) );
  INVX1 U26468 ( .A(reg_file[2065]), .Y(n35990) );
  NOR2X1 U26469 ( .A(n25968), .B(n35991), .Y(n23062) );
  INVX1 U26470 ( .A(reg_file[2066]), .Y(n35991) );
  NOR2X1 U26471 ( .A(n25968), .B(n35992), .Y(n23061) );
  INVX1 U26472 ( .A(reg_file[2067]), .Y(n35992) );
  NOR2X1 U26473 ( .A(n25968), .B(n35993), .Y(n23060) );
  INVX1 U26474 ( .A(reg_file[2068]), .Y(n35993) );
  NOR2X1 U26475 ( .A(n25968), .B(n35994), .Y(n23059) );
  INVX1 U26476 ( .A(reg_file[2069]), .Y(n35994) );
  NOR2X1 U26477 ( .A(n25968), .B(n35995), .Y(n23058) );
  INVX1 U26478 ( .A(reg_file[2070]), .Y(n35995) );
  NOR2X1 U26479 ( .A(n25968), .B(n35996), .Y(n23057) );
  INVX1 U26480 ( .A(reg_file[2071]), .Y(n35996) );
  NOR2X1 U26481 ( .A(n25968), .B(n35997), .Y(n23056) );
  INVX1 U26482 ( .A(reg_file[2072]), .Y(n35997) );
  NOR2X1 U26483 ( .A(n25968), .B(n35998), .Y(n23055) );
  INVX1 U26484 ( .A(reg_file[2073]), .Y(n35998) );
  NOR2X1 U26485 ( .A(n25968), .B(n35999), .Y(n23054) );
  INVX1 U26486 ( .A(reg_file[2074]), .Y(n35999) );
  NOR2X1 U26487 ( .A(n25968), .B(n36000), .Y(n23053) );
  INVX1 U26488 ( .A(reg_file[2075]), .Y(n36000) );
  NOR2X1 U26489 ( .A(n25968), .B(n36001), .Y(n23052) );
  INVX1 U26490 ( .A(reg_file[2076]), .Y(n36001) );
  NOR2X1 U26491 ( .A(n25968), .B(n36002), .Y(n23051) );
  INVX1 U26492 ( .A(reg_file[2077]), .Y(n36002) );
  NOR2X1 U26493 ( .A(n25968), .B(n36003), .Y(n23050) );
  INVX1 U26494 ( .A(reg_file[2078]), .Y(n36003) );
  NOR2X1 U26495 ( .A(n25969), .B(n36004), .Y(n23049) );
  INVX1 U26496 ( .A(reg_file[2079]), .Y(n36004) );
  NOR2X1 U26497 ( .A(n25969), .B(n36005), .Y(n23048) );
  INVX1 U26498 ( .A(reg_file[2080]), .Y(n36005) );
  NOR2X1 U26499 ( .A(n25969), .B(n36006), .Y(n23047) );
  INVX1 U26500 ( .A(reg_file[2081]), .Y(n36006) );
  NOR2X1 U26501 ( .A(n25969), .B(n36007), .Y(n23046) );
  INVX1 U26502 ( .A(reg_file[2082]), .Y(n36007) );
  NOR2X1 U26503 ( .A(n25969), .B(n36008), .Y(n23045) );
  INVX1 U26504 ( .A(reg_file[2083]), .Y(n36008) );
  NOR2X1 U26505 ( .A(n25969), .B(n36009), .Y(n23044) );
  INVX1 U26506 ( .A(reg_file[2084]), .Y(n36009) );
  NOR2X1 U26507 ( .A(n25969), .B(n36010), .Y(n23043) );
  INVX1 U26508 ( .A(reg_file[2085]), .Y(n36010) );
  NOR2X1 U26509 ( .A(n25969), .B(n36011), .Y(n23042) );
  INVX1 U26510 ( .A(reg_file[2086]), .Y(n36011) );
  NOR2X1 U26511 ( .A(n25969), .B(n36012), .Y(n23041) );
  INVX1 U26512 ( .A(reg_file[2087]), .Y(n36012) );
  NOR2X1 U26513 ( .A(n25969), .B(n36013), .Y(n23040) );
  INVX1 U26514 ( .A(reg_file[2088]), .Y(n36013) );
  NOR2X1 U26515 ( .A(n25969), .B(n36014), .Y(n23039) );
  INVX1 U26516 ( .A(reg_file[2089]), .Y(n36014) );
  NOR2X1 U26517 ( .A(n25969), .B(n36015), .Y(n23038) );
  INVX1 U26518 ( .A(reg_file[2090]), .Y(n36015) );
  NOR2X1 U26519 ( .A(n25969), .B(n36016), .Y(n23037) );
  INVX1 U26520 ( .A(reg_file[2091]), .Y(n36016) );
  NOR2X1 U26521 ( .A(n25969), .B(n36017), .Y(n23036) );
  INVX1 U26522 ( .A(reg_file[2092]), .Y(n36017) );
  NOR2X1 U26523 ( .A(n25969), .B(n36018), .Y(n23035) );
  INVX1 U26524 ( .A(reg_file[2093]), .Y(n36018) );
  NOR2X1 U26525 ( .A(n25969), .B(n36019), .Y(n23034) );
  INVX1 U26526 ( .A(reg_file[2094]), .Y(n36019) );
  NOR2X1 U26527 ( .A(n25969), .B(n36020), .Y(n23033) );
  INVX1 U26528 ( .A(reg_file[2095]), .Y(n36020) );
  NOR2X1 U26529 ( .A(n25970), .B(n36021), .Y(n23032) );
  INVX1 U26530 ( .A(reg_file[2096]), .Y(n36021) );
  NOR2X1 U26531 ( .A(n25970), .B(n36022), .Y(n23031) );
  INVX1 U26532 ( .A(reg_file[2097]), .Y(n36022) );
  NOR2X1 U26533 ( .A(n25970), .B(n36023), .Y(n23030) );
  INVX1 U26534 ( .A(reg_file[2098]), .Y(n36023) );
  NOR2X1 U26535 ( .A(n25970), .B(n36024), .Y(n23029) );
  INVX1 U26536 ( .A(reg_file[2099]), .Y(n36024) );
  NOR2X1 U26537 ( .A(n25970), .B(n36025), .Y(n23028) );
  INVX1 U26538 ( .A(reg_file[2100]), .Y(n36025) );
  NOR2X1 U26539 ( .A(n25970), .B(n36026), .Y(n23027) );
  INVX1 U26540 ( .A(reg_file[2101]), .Y(n36026) );
  NOR2X1 U26541 ( .A(n25970), .B(n36027), .Y(n23026) );
  INVX1 U26542 ( .A(reg_file[2102]), .Y(n36027) );
  NOR2X1 U26543 ( .A(n25970), .B(n36028), .Y(n23025) );
  INVX1 U26544 ( .A(reg_file[2103]), .Y(n36028) );
  NOR2X1 U26545 ( .A(n25970), .B(n36029), .Y(n23024) );
  INVX1 U26546 ( .A(reg_file[2104]), .Y(n36029) );
  NOR2X1 U26547 ( .A(n25970), .B(n36030), .Y(n23023) );
  INVX1 U26548 ( .A(reg_file[2105]), .Y(n36030) );
  NOR2X1 U26549 ( .A(n25970), .B(n36031), .Y(n23022) );
  INVX1 U26550 ( .A(reg_file[2106]), .Y(n36031) );
  NOR2X1 U26551 ( .A(n25970), .B(n36032), .Y(n23021) );
  INVX1 U26552 ( .A(reg_file[2107]), .Y(n36032) );
  NOR2X1 U26553 ( .A(n25970), .B(n36033), .Y(n23020) );
  INVX1 U26554 ( .A(reg_file[2108]), .Y(n36033) );
  NOR2X1 U26555 ( .A(n25970), .B(n36034), .Y(n23019) );
  INVX1 U26556 ( .A(reg_file[2109]), .Y(n36034) );
  NOR2X1 U26557 ( .A(n25970), .B(n36035), .Y(n23018) );
  INVX1 U26558 ( .A(reg_file[2110]), .Y(n36035) );
  NOR2X1 U26559 ( .A(n25970), .B(n36036), .Y(n23017) );
  INVX1 U26560 ( .A(reg_file[2111]), .Y(n36036) );
  NOR2X1 U26561 ( .A(n25970), .B(n36037), .Y(n23016) );
  INVX1 U26562 ( .A(reg_file[2112]), .Y(n36037) );
  NOR2X1 U26563 ( .A(n25971), .B(n36038), .Y(n23015) );
  INVX1 U26564 ( .A(reg_file[2113]), .Y(n36038) );
  NOR2X1 U26565 ( .A(n25971), .B(n36039), .Y(n23014) );
  INVX1 U26566 ( .A(reg_file[2114]), .Y(n36039) );
  NOR2X1 U26567 ( .A(n25971), .B(n36040), .Y(n23013) );
  INVX1 U26568 ( .A(reg_file[2115]), .Y(n36040) );
  NOR2X1 U26569 ( .A(n25971), .B(n36041), .Y(n23012) );
  INVX1 U26570 ( .A(reg_file[2116]), .Y(n36041) );
  NOR2X1 U26571 ( .A(n25971), .B(n36042), .Y(n23011) );
  INVX1 U26572 ( .A(reg_file[2117]), .Y(n36042) );
  NOR2X1 U26573 ( .A(n25971), .B(n36043), .Y(n23010) );
  INVX1 U26574 ( .A(reg_file[2118]), .Y(n36043) );
  NOR2X1 U26575 ( .A(n25971), .B(n36044), .Y(n23009) );
  INVX1 U26576 ( .A(reg_file[2119]), .Y(n36044) );
  NOR2X1 U26577 ( .A(n25971), .B(n36045), .Y(n23008) );
  INVX1 U26578 ( .A(reg_file[2120]), .Y(n36045) );
  NOR2X1 U26579 ( .A(n25971), .B(n36046), .Y(n23007) );
  INVX1 U26580 ( .A(reg_file[2121]), .Y(n36046) );
  NOR2X1 U26581 ( .A(n25971), .B(n36047), .Y(n23006) );
  INVX1 U26582 ( .A(reg_file[2122]), .Y(n36047) );
  NOR2X1 U26583 ( .A(n25971), .B(n36048), .Y(n23005) );
  INVX1 U26584 ( .A(reg_file[2123]), .Y(n36048) );
  NOR2X1 U26585 ( .A(n25971), .B(n36049), .Y(n23004) );
  INVX1 U26586 ( .A(reg_file[2124]), .Y(n36049) );
  NOR2X1 U26587 ( .A(n25971), .B(n36050), .Y(n23003) );
  INVX1 U26588 ( .A(reg_file[2125]), .Y(n36050) );
  NOR2X1 U26589 ( .A(n25971), .B(n36051), .Y(n23002) );
  INVX1 U26590 ( .A(reg_file[2126]), .Y(n36051) );
  NOR2X1 U26591 ( .A(n25971), .B(n36052), .Y(n23001) );
  INVX1 U26592 ( .A(reg_file[2127]), .Y(n36052) );
  NOR2X1 U26593 ( .A(n25971), .B(n36053), .Y(n23000) );
  INVX1 U26594 ( .A(reg_file[2128]), .Y(n36053) );
  NOR2X1 U26595 ( .A(n25971), .B(n36054), .Y(n22999) );
  INVX1 U26596 ( .A(reg_file[2129]), .Y(n36054) );
  NOR2X1 U26597 ( .A(n25972), .B(n36055), .Y(n22998) );
  INVX1 U26598 ( .A(reg_file[2130]), .Y(n36055) );
  NOR2X1 U26599 ( .A(n25972), .B(n36056), .Y(n22997) );
  INVX1 U26600 ( .A(reg_file[2131]), .Y(n36056) );
  NOR2X1 U26601 ( .A(n25972), .B(n36057), .Y(n22996) );
  INVX1 U26602 ( .A(reg_file[2132]), .Y(n36057) );
  NOR2X1 U26603 ( .A(n25972), .B(n36058), .Y(n22995) );
  INVX1 U26604 ( .A(reg_file[2133]), .Y(n36058) );
  NOR2X1 U26605 ( .A(n25972), .B(n36059), .Y(n22994) );
  INVX1 U26606 ( .A(reg_file[2134]), .Y(n36059) );
  NOR2X1 U26607 ( .A(n25972), .B(n36060), .Y(n22993) );
  INVX1 U26608 ( .A(reg_file[2135]), .Y(n36060) );
  NOR2X1 U26609 ( .A(n25972), .B(n36061), .Y(n22992) );
  INVX1 U26610 ( .A(reg_file[2136]), .Y(n36061) );
  NOR2X1 U26611 ( .A(n25972), .B(n36062), .Y(n22991) );
  INVX1 U26612 ( .A(reg_file[2137]), .Y(n36062) );
  NOR2X1 U26613 ( .A(n25972), .B(n36063), .Y(n22990) );
  INVX1 U26614 ( .A(reg_file[2138]), .Y(n36063) );
  NOR2X1 U26615 ( .A(n25972), .B(n36064), .Y(n22989) );
  INVX1 U26616 ( .A(reg_file[2139]), .Y(n36064) );
  NOR2X1 U26617 ( .A(n25972), .B(n36065), .Y(n22988) );
  INVX1 U26618 ( .A(reg_file[2140]), .Y(n36065) );
  NOR2X1 U26619 ( .A(n25972), .B(n36066), .Y(n22987) );
  INVX1 U26620 ( .A(reg_file[2141]), .Y(n36066) );
  NOR2X1 U26621 ( .A(n25972), .B(n36067), .Y(n22986) );
  INVX1 U26622 ( .A(reg_file[2142]), .Y(n36067) );
  NOR2X1 U26623 ( .A(n25972), .B(n36068), .Y(n22985) );
  INVX1 U26624 ( .A(reg_file[2143]), .Y(n36068) );
  NOR2X1 U26625 ( .A(n25972), .B(n36069), .Y(n22984) );
  INVX1 U26626 ( .A(reg_file[2144]), .Y(n36069) );
  NOR2X1 U26627 ( .A(n25972), .B(n36070), .Y(n22983) );
  INVX1 U26628 ( .A(reg_file[2145]), .Y(n36070) );
  NOR2X1 U26629 ( .A(n25972), .B(n36071), .Y(n22982) );
  INVX1 U26630 ( .A(reg_file[2146]), .Y(n36071) );
  NOR2X1 U26631 ( .A(n25973), .B(n36072), .Y(n22981) );
  INVX1 U26632 ( .A(reg_file[2147]), .Y(n36072) );
  NOR2X1 U26633 ( .A(n25973), .B(n36073), .Y(n22980) );
  INVX1 U26634 ( .A(reg_file[2148]), .Y(n36073) );
  NOR2X1 U26635 ( .A(n25973), .B(n36074), .Y(n22979) );
  INVX1 U26636 ( .A(reg_file[2149]), .Y(n36074) );
  NOR2X1 U26637 ( .A(n25973), .B(n36075), .Y(n22978) );
  INVX1 U26638 ( .A(reg_file[2150]), .Y(n36075) );
  NOR2X1 U26639 ( .A(n25973), .B(n36076), .Y(n22977) );
  INVX1 U26640 ( .A(reg_file[2151]), .Y(n36076) );
  NOR2X1 U26641 ( .A(n25973), .B(n36077), .Y(n22976) );
  INVX1 U26642 ( .A(reg_file[2152]), .Y(n36077) );
  NOR2X1 U26643 ( .A(n25973), .B(n36078), .Y(n22975) );
  INVX1 U26644 ( .A(reg_file[2153]), .Y(n36078) );
  NOR2X1 U26645 ( .A(n25973), .B(n36079), .Y(n22974) );
  INVX1 U26646 ( .A(reg_file[2154]), .Y(n36079) );
  NOR2X1 U26647 ( .A(n25973), .B(n36080), .Y(n22973) );
  INVX1 U26648 ( .A(reg_file[2155]), .Y(n36080) );
  NOR2X1 U26649 ( .A(n25973), .B(n36081), .Y(n22972) );
  INVX1 U26650 ( .A(reg_file[2156]), .Y(n36081) );
  NOR2X1 U26651 ( .A(n25973), .B(n36082), .Y(n22971) );
  INVX1 U26652 ( .A(reg_file[2157]), .Y(n36082) );
  NOR2X1 U26653 ( .A(n25973), .B(n36083), .Y(n22970) );
  INVX1 U26654 ( .A(reg_file[2158]), .Y(n36083) );
  NOR2X1 U26655 ( .A(n25973), .B(n36084), .Y(n22969) );
  INVX1 U26656 ( .A(reg_file[2159]), .Y(n36084) );
  NOR2X1 U26657 ( .A(n25973), .B(n36085), .Y(n22968) );
  INVX1 U26658 ( .A(reg_file[2160]), .Y(n36085) );
  NOR2X1 U26659 ( .A(n25973), .B(n36086), .Y(n22967) );
  INVX1 U26660 ( .A(reg_file[2161]), .Y(n36086) );
  NOR2X1 U26661 ( .A(n25973), .B(n36087), .Y(n22966) );
  INVX1 U26662 ( .A(reg_file[2162]), .Y(n36087) );
  NOR2X1 U26663 ( .A(n25973), .B(n36088), .Y(n22965) );
  INVX1 U26664 ( .A(reg_file[2163]), .Y(n36088) );
  NOR2X1 U26665 ( .A(n25974), .B(n36089), .Y(n22964) );
  INVX1 U26666 ( .A(reg_file[2164]), .Y(n36089) );
  NOR2X1 U26667 ( .A(n25974), .B(n36090), .Y(n22963) );
  INVX1 U26668 ( .A(reg_file[2165]), .Y(n36090) );
  NOR2X1 U26669 ( .A(n25974), .B(n36091), .Y(n22962) );
  INVX1 U26670 ( .A(reg_file[2166]), .Y(n36091) );
  NOR2X1 U26671 ( .A(n25974), .B(n36092), .Y(n22961) );
  INVX1 U26672 ( .A(reg_file[2167]), .Y(n36092) );
  NOR2X1 U26673 ( .A(n25974), .B(n36093), .Y(n22960) );
  INVX1 U26674 ( .A(reg_file[2168]), .Y(n36093) );
  NOR2X1 U26675 ( .A(n25974), .B(n36094), .Y(n22959) );
  INVX1 U26676 ( .A(reg_file[2169]), .Y(n36094) );
  NOR2X1 U26677 ( .A(n25974), .B(n36095), .Y(n22958) );
  INVX1 U26678 ( .A(reg_file[2170]), .Y(n36095) );
  NOR2X1 U26679 ( .A(n25974), .B(n36096), .Y(n22957) );
  INVX1 U26680 ( .A(reg_file[2171]), .Y(n36096) );
  NOR2X1 U26681 ( .A(n25974), .B(n36097), .Y(n22956) );
  INVX1 U26682 ( .A(reg_file[2172]), .Y(n36097) );
  NOR2X1 U26683 ( .A(n25974), .B(n36098), .Y(n22955) );
  INVX1 U26684 ( .A(reg_file[2173]), .Y(n36098) );
  NOR2X1 U26685 ( .A(n25974), .B(n36099), .Y(n22954) );
  INVX1 U26686 ( .A(reg_file[2174]), .Y(n36099) );
  NOR2X1 U26687 ( .A(n25974), .B(n36100), .Y(n22953) );
  INVX1 U26688 ( .A(reg_file[2175]), .Y(n36100) );
  NOR2X1 U26689 ( .A(n36101), .B(n34923), .Y(n35973) );
  MUX2X1 U26690 ( .B(n36102), .A(n25129), .S(n25975), .Y(n22952) );
  INVX1 U26691 ( .A(reg_file[2176]), .Y(n36102) );
  MUX2X1 U26692 ( .B(n36104), .A(n25130), .S(n25975), .Y(n22951) );
  INVX1 U26693 ( .A(reg_file[2177]), .Y(n36104) );
  MUX2X1 U26694 ( .B(n36105), .A(n25131), .S(n25975), .Y(n22950) );
  INVX1 U26695 ( .A(reg_file[2178]), .Y(n36105) );
  MUX2X1 U26696 ( .B(n36106), .A(n25132), .S(n25975), .Y(n22949) );
  INVX1 U26697 ( .A(reg_file[2179]), .Y(n36106) );
  MUX2X1 U26698 ( .B(n36107), .A(n25133), .S(n25975), .Y(n22948) );
  INVX1 U26699 ( .A(reg_file[2180]), .Y(n36107) );
  MUX2X1 U26700 ( .B(n36108), .A(n25134), .S(n25975), .Y(n22947) );
  INVX1 U26701 ( .A(reg_file[2181]), .Y(n36108) );
  MUX2X1 U26702 ( .B(n36109), .A(n25135), .S(n25975), .Y(n22946) );
  INVX1 U26703 ( .A(reg_file[2182]), .Y(n36109) );
  MUX2X1 U26704 ( .B(n36110), .A(n25136), .S(n25975), .Y(n22945) );
  INVX1 U26705 ( .A(reg_file[2183]), .Y(n36110) );
  NOR2X1 U26706 ( .A(n25975), .B(n36111), .Y(n22944) );
  INVX1 U26707 ( .A(reg_file[2184]), .Y(n36111) );
  NOR2X1 U26708 ( .A(n25975), .B(n36112), .Y(n22943) );
  INVX1 U26709 ( .A(reg_file[2185]), .Y(n36112) );
  NOR2X1 U26710 ( .A(n25975), .B(n36113), .Y(n22942) );
  INVX1 U26711 ( .A(reg_file[2186]), .Y(n36113) );
  NOR2X1 U26712 ( .A(n25975), .B(n36114), .Y(n22941) );
  INVX1 U26713 ( .A(reg_file[2187]), .Y(n36114) );
  NOR2X1 U26714 ( .A(n25975), .B(n36115), .Y(n22940) );
  INVX1 U26715 ( .A(reg_file[2188]), .Y(n36115) );
  NOR2X1 U26716 ( .A(n25975), .B(n36116), .Y(n22939) );
  INVX1 U26717 ( .A(reg_file[2189]), .Y(n36116) );
  NOR2X1 U26718 ( .A(n25976), .B(n36117), .Y(n22938) );
  INVX1 U26719 ( .A(reg_file[2190]), .Y(n36117) );
  NOR2X1 U26720 ( .A(n25976), .B(n36118), .Y(n22937) );
  INVX1 U26721 ( .A(reg_file[2191]), .Y(n36118) );
  NOR2X1 U26722 ( .A(n25976), .B(n36119), .Y(n22936) );
  INVX1 U26723 ( .A(reg_file[2192]), .Y(n36119) );
  NOR2X1 U26724 ( .A(n25976), .B(n36120), .Y(n22935) );
  INVX1 U26725 ( .A(reg_file[2193]), .Y(n36120) );
  NOR2X1 U26726 ( .A(n25976), .B(n36121), .Y(n22934) );
  INVX1 U26727 ( .A(reg_file[2194]), .Y(n36121) );
  NOR2X1 U26728 ( .A(n25976), .B(n36122), .Y(n22933) );
  INVX1 U26729 ( .A(reg_file[2195]), .Y(n36122) );
  NOR2X1 U26730 ( .A(n25976), .B(n36123), .Y(n22932) );
  INVX1 U26731 ( .A(reg_file[2196]), .Y(n36123) );
  NOR2X1 U26732 ( .A(n25976), .B(n36124), .Y(n22931) );
  INVX1 U26733 ( .A(reg_file[2197]), .Y(n36124) );
  NOR2X1 U26734 ( .A(n25976), .B(n36125), .Y(n22930) );
  INVX1 U26735 ( .A(reg_file[2198]), .Y(n36125) );
  NOR2X1 U26736 ( .A(n25976), .B(n36126), .Y(n22929) );
  INVX1 U26737 ( .A(reg_file[2199]), .Y(n36126) );
  NOR2X1 U26738 ( .A(n25976), .B(n36127), .Y(n22928) );
  INVX1 U26739 ( .A(reg_file[2200]), .Y(n36127) );
  NOR2X1 U26740 ( .A(n25976), .B(n36128), .Y(n22927) );
  INVX1 U26741 ( .A(reg_file[2201]), .Y(n36128) );
  NOR2X1 U26742 ( .A(n25976), .B(n36129), .Y(n22926) );
  INVX1 U26743 ( .A(reg_file[2202]), .Y(n36129) );
  NOR2X1 U26744 ( .A(n25976), .B(n36130), .Y(n22925) );
  INVX1 U26745 ( .A(reg_file[2203]), .Y(n36130) );
  NOR2X1 U26746 ( .A(n25976), .B(n36131), .Y(n22924) );
  INVX1 U26747 ( .A(reg_file[2204]), .Y(n36131) );
  NOR2X1 U26748 ( .A(n25976), .B(n36132), .Y(n22923) );
  INVX1 U26749 ( .A(reg_file[2205]), .Y(n36132) );
  NOR2X1 U26750 ( .A(n25976), .B(n36133), .Y(n22922) );
  INVX1 U26751 ( .A(reg_file[2206]), .Y(n36133) );
  NOR2X1 U26752 ( .A(n25977), .B(n36134), .Y(n22921) );
  INVX1 U26753 ( .A(reg_file[2207]), .Y(n36134) );
  NOR2X1 U26754 ( .A(n25977), .B(n36135), .Y(n22920) );
  INVX1 U26755 ( .A(reg_file[2208]), .Y(n36135) );
  NOR2X1 U26756 ( .A(n25977), .B(n36136), .Y(n22919) );
  INVX1 U26757 ( .A(reg_file[2209]), .Y(n36136) );
  NOR2X1 U26758 ( .A(n25977), .B(n36137), .Y(n22918) );
  INVX1 U26759 ( .A(reg_file[2210]), .Y(n36137) );
  NOR2X1 U26760 ( .A(n25977), .B(n36138), .Y(n22917) );
  INVX1 U26761 ( .A(reg_file[2211]), .Y(n36138) );
  NOR2X1 U26762 ( .A(n25977), .B(n36139), .Y(n22916) );
  INVX1 U26763 ( .A(reg_file[2212]), .Y(n36139) );
  NOR2X1 U26764 ( .A(n25977), .B(n36140), .Y(n22915) );
  INVX1 U26765 ( .A(reg_file[2213]), .Y(n36140) );
  NOR2X1 U26766 ( .A(n25977), .B(n36141), .Y(n22914) );
  INVX1 U26767 ( .A(reg_file[2214]), .Y(n36141) );
  NOR2X1 U26768 ( .A(n25977), .B(n36142), .Y(n22913) );
  INVX1 U26769 ( .A(reg_file[2215]), .Y(n36142) );
  NOR2X1 U26770 ( .A(n25977), .B(n36143), .Y(n22912) );
  INVX1 U26771 ( .A(reg_file[2216]), .Y(n36143) );
  NOR2X1 U26772 ( .A(n25977), .B(n36144), .Y(n22911) );
  INVX1 U26773 ( .A(reg_file[2217]), .Y(n36144) );
  NOR2X1 U26774 ( .A(n25977), .B(n36145), .Y(n22910) );
  INVX1 U26775 ( .A(reg_file[2218]), .Y(n36145) );
  NOR2X1 U26776 ( .A(n25977), .B(n36146), .Y(n22909) );
  INVX1 U26777 ( .A(reg_file[2219]), .Y(n36146) );
  NOR2X1 U26778 ( .A(n25977), .B(n36147), .Y(n22908) );
  INVX1 U26779 ( .A(reg_file[2220]), .Y(n36147) );
  NOR2X1 U26780 ( .A(n25977), .B(n36148), .Y(n22907) );
  INVX1 U26781 ( .A(reg_file[2221]), .Y(n36148) );
  NOR2X1 U26782 ( .A(n25977), .B(n36149), .Y(n22906) );
  INVX1 U26783 ( .A(reg_file[2222]), .Y(n36149) );
  NOR2X1 U26784 ( .A(n25977), .B(n36150), .Y(n22905) );
  INVX1 U26785 ( .A(reg_file[2223]), .Y(n36150) );
  NOR2X1 U26786 ( .A(n25978), .B(n36151), .Y(n22904) );
  INVX1 U26787 ( .A(reg_file[2224]), .Y(n36151) );
  NOR2X1 U26788 ( .A(n25978), .B(n36152), .Y(n22903) );
  INVX1 U26789 ( .A(reg_file[2225]), .Y(n36152) );
  NOR2X1 U26790 ( .A(n25978), .B(n36153), .Y(n22902) );
  INVX1 U26791 ( .A(reg_file[2226]), .Y(n36153) );
  NOR2X1 U26792 ( .A(n25978), .B(n36154), .Y(n22901) );
  INVX1 U26793 ( .A(reg_file[2227]), .Y(n36154) );
  NOR2X1 U26794 ( .A(n25978), .B(n36155), .Y(n22900) );
  INVX1 U26795 ( .A(reg_file[2228]), .Y(n36155) );
  NOR2X1 U26796 ( .A(n25978), .B(n36156), .Y(n22899) );
  INVX1 U26797 ( .A(reg_file[2229]), .Y(n36156) );
  NOR2X1 U26798 ( .A(n25978), .B(n36157), .Y(n22898) );
  INVX1 U26799 ( .A(reg_file[2230]), .Y(n36157) );
  NOR2X1 U26800 ( .A(n25978), .B(n36158), .Y(n22897) );
  INVX1 U26801 ( .A(reg_file[2231]), .Y(n36158) );
  NOR2X1 U26802 ( .A(n25978), .B(n36159), .Y(n22896) );
  INVX1 U26803 ( .A(reg_file[2232]), .Y(n36159) );
  NOR2X1 U26804 ( .A(n25978), .B(n36160), .Y(n22895) );
  INVX1 U26805 ( .A(reg_file[2233]), .Y(n36160) );
  NOR2X1 U26806 ( .A(n25978), .B(n36161), .Y(n22894) );
  INVX1 U26807 ( .A(reg_file[2234]), .Y(n36161) );
  NOR2X1 U26808 ( .A(n25978), .B(n36162), .Y(n22893) );
  INVX1 U26809 ( .A(reg_file[2235]), .Y(n36162) );
  NOR2X1 U26810 ( .A(n25978), .B(n36163), .Y(n22892) );
  INVX1 U26811 ( .A(reg_file[2236]), .Y(n36163) );
  NOR2X1 U26812 ( .A(n25978), .B(n36164), .Y(n22891) );
  INVX1 U26813 ( .A(reg_file[2237]), .Y(n36164) );
  NOR2X1 U26814 ( .A(n25978), .B(n36165), .Y(n22890) );
  INVX1 U26815 ( .A(reg_file[2238]), .Y(n36165) );
  NOR2X1 U26816 ( .A(n25978), .B(n36166), .Y(n22889) );
  INVX1 U26817 ( .A(reg_file[2239]), .Y(n36166) );
  NOR2X1 U26818 ( .A(n25978), .B(n36167), .Y(n22888) );
  INVX1 U26819 ( .A(reg_file[2240]), .Y(n36167) );
  NOR2X1 U26820 ( .A(n25979), .B(n36168), .Y(n22887) );
  INVX1 U26821 ( .A(reg_file[2241]), .Y(n36168) );
  NOR2X1 U26822 ( .A(n25979), .B(n36169), .Y(n22886) );
  INVX1 U26823 ( .A(reg_file[2242]), .Y(n36169) );
  NOR2X1 U26824 ( .A(n25979), .B(n36170), .Y(n22885) );
  INVX1 U26825 ( .A(reg_file[2243]), .Y(n36170) );
  NOR2X1 U26826 ( .A(n25979), .B(n36171), .Y(n22884) );
  INVX1 U26827 ( .A(reg_file[2244]), .Y(n36171) );
  NOR2X1 U26828 ( .A(n25979), .B(n36172), .Y(n22883) );
  INVX1 U26829 ( .A(reg_file[2245]), .Y(n36172) );
  NOR2X1 U26830 ( .A(n25979), .B(n36173), .Y(n22882) );
  INVX1 U26831 ( .A(reg_file[2246]), .Y(n36173) );
  NOR2X1 U26832 ( .A(n25979), .B(n36174), .Y(n22881) );
  INVX1 U26833 ( .A(reg_file[2247]), .Y(n36174) );
  NOR2X1 U26834 ( .A(n25979), .B(n36175), .Y(n22880) );
  INVX1 U26835 ( .A(reg_file[2248]), .Y(n36175) );
  NOR2X1 U26836 ( .A(n25979), .B(n36176), .Y(n22879) );
  INVX1 U26837 ( .A(reg_file[2249]), .Y(n36176) );
  NOR2X1 U26838 ( .A(n25979), .B(n36177), .Y(n22878) );
  INVX1 U26839 ( .A(reg_file[2250]), .Y(n36177) );
  NOR2X1 U26840 ( .A(n25979), .B(n36178), .Y(n22877) );
  INVX1 U26841 ( .A(reg_file[2251]), .Y(n36178) );
  NOR2X1 U26842 ( .A(n25979), .B(n36179), .Y(n22876) );
  INVX1 U26843 ( .A(reg_file[2252]), .Y(n36179) );
  NOR2X1 U26844 ( .A(n25979), .B(n36180), .Y(n22875) );
  INVX1 U26845 ( .A(reg_file[2253]), .Y(n36180) );
  NOR2X1 U26846 ( .A(n25979), .B(n36181), .Y(n22874) );
  INVX1 U26847 ( .A(reg_file[2254]), .Y(n36181) );
  NOR2X1 U26848 ( .A(n25979), .B(n36182), .Y(n22873) );
  INVX1 U26849 ( .A(reg_file[2255]), .Y(n36182) );
  NOR2X1 U26850 ( .A(n25979), .B(n36183), .Y(n22872) );
  INVX1 U26851 ( .A(reg_file[2256]), .Y(n36183) );
  NOR2X1 U26852 ( .A(n25979), .B(n36184), .Y(n22871) );
  INVX1 U26853 ( .A(reg_file[2257]), .Y(n36184) );
  NOR2X1 U26854 ( .A(n25980), .B(n36185), .Y(n22870) );
  INVX1 U26855 ( .A(reg_file[2258]), .Y(n36185) );
  NOR2X1 U26856 ( .A(n25980), .B(n36186), .Y(n22869) );
  INVX1 U26857 ( .A(reg_file[2259]), .Y(n36186) );
  NOR2X1 U26858 ( .A(n25980), .B(n36187), .Y(n22868) );
  INVX1 U26859 ( .A(reg_file[2260]), .Y(n36187) );
  NOR2X1 U26860 ( .A(n25980), .B(n36188), .Y(n22867) );
  INVX1 U26861 ( .A(reg_file[2261]), .Y(n36188) );
  NOR2X1 U26862 ( .A(n25980), .B(n36189), .Y(n22866) );
  INVX1 U26863 ( .A(reg_file[2262]), .Y(n36189) );
  NOR2X1 U26864 ( .A(n25980), .B(n36190), .Y(n22865) );
  INVX1 U26865 ( .A(reg_file[2263]), .Y(n36190) );
  NOR2X1 U26866 ( .A(n25980), .B(n36191), .Y(n22864) );
  INVX1 U26867 ( .A(reg_file[2264]), .Y(n36191) );
  NOR2X1 U26868 ( .A(n25980), .B(n36192), .Y(n22863) );
  INVX1 U26869 ( .A(reg_file[2265]), .Y(n36192) );
  NOR2X1 U26870 ( .A(n25980), .B(n36193), .Y(n22862) );
  INVX1 U26871 ( .A(reg_file[2266]), .Y(n36193) );
  NOR2X1 U26872 ( .A(n25980), .B(n36194), .Y(n22861) );
  INVX1 U26873 ( .A(reg_file[2267]), .Y(n36194) );
  NOR2X1 U26874 ( .A(n25980), .B(n36195), .Y(n22860) );
  INVX1 U26875 ( .A(reg_file[2268]), .Y(n36195) );
  NOR2X1 U26876 ( .A(n25980), .B(n36196), .Y(n22859) );
  INVX1 U26877 ( .A(reg_file[2269]), .Y(n36196) );
  NOR2X1 U26878 ( .A(n25980), .B(n36197), .Y(n22858) );
  INVX1 U26879 ( .A(reg_file[2270]), .Y(n36197) );
  NOR2X1 U26880 ( .A(n25980), .B(n36198), .Y(n22857) );
  INVX1 U26881 ( .A(reg_file[2271]), .Y(n36198) );
  NOR2X1 U26882 ( .A(n25980), .B(n36199), .Y(n22856) );
  INVX1 U26883 ( .A(reg_file[2272]), .Y(n36199) );
  NOR2X1 U26884 ( .A(n25980), .B(n36200), .Y(n22855) );
  INVX1 U26885 ( .A(reg_file[2273]), .Y(n36200) );
  NOR2X1 U26886 ( .A(n25980), .B(n36201), .Y(n22854) );
  INVX1 U26887 ( .A(reg_file[2274]), .Y(n36201) );
  NOR2X1 U26888 ( .A(n25981), .B(n36202), .Y(n22853) );
  INVX1 U26889 ( .A(reg_file[2275]), .Y(n36202) );
  NOR2X1 U26890 ( .A(n25981), .B(n36203), .Y(n22852) );
  INVX1 U26891 ( .A(reg_file[2276]), .Y(n36203) );
  NOR2X1 U26892 ( .A(n25981), .B(n36204), .Y(n22851) );
  INVX1 U26893 ( .A(reg_file[2277]), .Y(n36204) );
  NOR2X1 U26894 ( .A(n25981), .B(n36205), .Y(n22850) );
  INVX1 U26895 ( .A(reg_file[2278]), .Y(n36205) );
  NOR2X1 U26896 ( .A(n25981), .B(n36206), .Y(n22849) );
  INVX1 U26897 ( .A(reg_file[2279]), .Y(n36206) );
  NOR2X1 U26898 ( .A(n25981), .B(n36207), .Y(n22848) );
  INVX1 U26899 ( .A(reg_file[2280]), .Y(n36207) );
  NOR2X1 U26900 ( .A(n25981), .B(n36208), .Y(n22847) );
  INVX1 U26901 ( .A(reg_file[2281]), .Y(n36208) );
  NOR2X1 U26902 ( .A(n25981), .B(n36209), .Y(n22846) );
  INVX1 U26903 ( .A(reg_file[2282]), .Y(n36209) );
  NOR2X1 U26904 ( .A(n25981), .B(n36210), .Y(n22845) );
  INVX1 U26905 ( .A(reg_file[2283]), .Y(n36210) );
  NOR2X1 U26906 ( .A(n25981), .B(n36211), .Y(n22844) );
  INVX1 U26907 ( .A(reg_file[2284]), .Y(n36211) );
  NOR2X1 U26908 ( .A(n25981), .B(n36212), .Y(n22843) );
  INVX1 U26909 ( .A(reg_file[2285]), .Y(n36212) );
  NOR2X1 U26910 ( .A(n25981), .B(n36213), .Y(n22842) );
  INVX1 U26911 ( .A(reg_file[2286]), .Y(n36213) );
  NOR2X1 U26912 ( .A(n25981), .B(n36214), .Y(n22841) );
  INVX1 U26913 ( .A(reg_file[2287]), .Y(n36214) );
  NOR2X1 U26914 ( .A(n25981), .B(n36215), .Y(n22840) );
  INVX1 U26915 ( .A(reg_file[2288]), .Y(n36215) );
  NOR2X1 U26916 ( .A(n25981), .B(n36216), .Y(n22839) );
  INVX1 U26917 ( .A(reg_file[2289]), .Y(n36216) );
  NOR2X1 U26918 ( .A(n25981), .B(n36217), .Y(n22838) );
  INVX1 U26919 ( .A(reg_file[2290]), .Y(n36217) );
  NOR2X1 U26920 ( .A(n25981), .B(n36218), .Y(n22837) );
  INVX1 U26921 ( .A(reg_file[2291]), .Y(n36218) );
  NOR2X1 U26922 ( .A(n25982), .B(n36219), .Y(n22836) );
  INVX1 U26923 ( .A(reg_file[2292]), .Y(n36219) );
  NOR2X1 U26924 ( .A(n25982), .B(n36220), .Y(n22835) );
  INVX1 U26925 ( .A(reg_file[2293]), .Y(n36220) );
  NOR2X1 U26926 ( .A(n25982), .B(n36221), .Y(n22834) );
  INVX1 U26927 ( .A(reg_file[2294]), .Y(n36221) );
  NOR2X1 U26928 ( .A(n25982), .B(n36222), .Y(n22833) );
  INVX1 U26929 ( .A(reg_file[2295]), .Y(n36222) );
  NOR2X1 U26930 ( .A(n25982), .B(n36223), .Y(n22832) );
  INVX1 U26931 ( .A(reg_file[2296]), .Y(n36223) );
  NOR2X1 U26932 ( .A(n25982), .B(n36224), .Y(n22831) );
  INVX1 U26933 ( .A(reg_file[2297]), .Y(n36224) );
  NOR2X1 U26934 ( .A(n25982), .B(n36225), .Y(n22830) );
  INVX1 U26935 ( .A(reg_file[2298]), .Y(n36225) );
  NOR2X1 U26936 ( .A(n25982), .B(n36226), .Y(n22829) );
  INVX1 U26937 ( .A(reg_file[2299]), .Y(n36226) );
  NOR2X1 U26938 ( .A(n25982), .B(n36227), .Y(n22828) );
  INVX1 U26939 ( .A(reg_file[2300]), .Y(n36227) );
  NOR2X1 U26940 ( .A(n25982), .B(n36228), .Y(n22827) );
  INVX1 U26941 ( .A(reg_file[2301]), .Y(n36228) );
  NOR2X1 U26942 ( .A(n25982), .B(n36229), .Y(n22826) );
  INVX1 U26943 ( .A(reg_file[2302]), .Y(n36229) );
  NOR2X1 U26944 ( .A(n25982), .B(n36230), .Y(n22825) );
  INVX1 U26945 ( .A(reg_file[2303]), .Y(n36230) );
  NOR2X1 U26946 ( .A(n36231), .B(n34923), .Y(n36103) );
  MUX2X1 U26947 ( .B(n36232), .A(n25129), .S(n25983), .Y(n22824) );
  INVX1 U26948 ( .A(reg_file[2304]), .Y(n36232) );
  MUX2X1 U26949 ( .B(n36234), .A(n25130), .S(n25983), .Y(n22823) );
  INVX1 U26950 ( .A(reg_file[2305]), .Y(n36234) );
  MUX2X1 U26951 ( .B(n36235), .A(n25131), .S(n25983), .Y(n22822) );
  INVX1 U26952 ( .A(reg_file[2306]), .Y(n36235) );
  MUX2X1 U26953 ( .B(n36236), .A(n25132), .S(n25983), .Y(n22821) );
  INVX1 U26954 ( .A(reg_file[2307]), .Y(n36236) );
  MUX2X1 U26955 ( .B(n36237), .A(n25133), .S(n25983), .Y(n22820) );
  INVX1 U26956 ( .A(reg_file[2308]), .Y(n36237) );
  MUX2X1 U26957 ( .B(n36238), .A(n25134), .S(n25983), .Y(n22819) );
  INVX1 U26958 ( .A(reg_file[2309]), .Y(n36238) );
  MUX2X1 U26959 ( .B(n36239), .A(n25135), .S(n25983), .Y(n22818) );
  INVX1 U26960 ( .A(reg_file[2310]), .Y(n36239) );
  MUX2X1 U26961 ( .B(n36240), .A(n25136), .S(n25983), .Y(n22817) );
  INVX1 U26962 ( .A(reg_file[2311]), .Y(n36240) );
  NOR2X1 U26963 ( .A(n25983), .B(n36241), .Y(n22816) );
  INVX1 U26964 ( .A(reg_file[2312]), .Y(n36241) );
  NOR2X1 U26965 ( .A(n25983), .B(n36242), .Y(n22815) );
  INVX1 U26966 ( .A(reg_file[2313]), .Y(n36242) );
  NOR2X1 U26967 ( .A(n25983), .B(n36243), .Y(n22814) );
  INVX1 U26968 ( .A(reg_file[2314]), .Y(n36243) );
  NOR2X1 U26969 ( .A(n25983), .B(n36244), .Y(n22813) );
  INVX1 U26970 ( .A(reg_file[2315]), .Y(n36244) );
  NOR2X1 U26971 ( .A(n25983), .B(n36245), .Y(n22812) );
  INVX1 U26972 ( .A(reg_file[2316]), .Y(n36245) );
  NOR2X1 U26973 ( .A(n25983), .B(n36246), .Y(n22811) );
  INVX1 U26974 ( .A(reg_file[2317]), .Y(n36246) );
  NOR2X1 U26975 ( .A(n25984), .B(n36247), .Y(n22810) );
  INVX1 U26976 ( .A(reg_file[2318]), .Y(n36247) );
  NOR2X1 U26977 ( .A(n25984), .B(n36248), .Y(n22809) );
  INVX1 U26978 ( .A(reg_file[2319]), .Y(n36248) );
  NOR2X1 U26979 ( .A(n25984), .B(n36249), .Y(n22808) );
  INVX1 U26980 ( .A(reg_file[2320]), .Y(n36249) );
  NOR2X1 U26981 ( .A(n25984), .B(n36250), .Y(n22807) );
  INVX1 U26982 ( .A(reg_file[2321]), .Y(n36250) );
  NOR2X1 U26983 ( .A(n25984), .B(n36251), .Y(n22806) );
  INVX1 U26984 ( .A(reg_file[2322]), .Y(n36251) );
  NOR2X1 U26985 ( .A(n25984), .B(n36252), .Y(n22805) );
  INVX1 U26986 ( .A(reg_file[2323]), .Y(n36252) );
  NOR2X1 U26987 ( .A(n25984), .B(n36253), .Y(n22804) );
  INVX1 U26988 ( .A(reg_file[2324]), .Y(n36253) );
  NOR2X1 U26989 ( .A(n25984), .B(n36254), .Y(n22803) );
  INVX1 U26990 ( .A(reg_file[2325]), .Y(n36254) );
  NOR2X1 U26991 ( .A(n25984), .B(n36255), .Y(n22802) );
  INVX1 U26992 ( .A(reg_file[2326]), .Y(n36255) );
  NOR2X1 U26993 ( .A(n25984), .B(n36256), .Y(n22801) );
  INVX1 U26994 ( .A(reg_file[2327]), .Y(n36256) );
  NOR2X1 U26995 ( .A(n25984), .B(n36257), .Y(n22800) );
  INVX1 U26996 ( .A(reg_file[2328]), .Y(n36257) );
  NOR2X1 U26997 ( .A(n25984), .B(n36258), .Y(n22799) );
  INVX1 U26998 ( .A(reg_file[2329]), .Y(n36258) );
  NOR2X1 U26999 ( .A(n25984), .B(n36259), .Y(n22798) );
  INVX1 U27000 ( .A(reg_file[2330]), .Y(n36259) );
  NOR2X1 U27001 ( .A(n25984), .B(n36260), .Y(n22797) );
  INVX1 U27002 ( .A(reg_file[2331]), .Y(n36260) );
  NOR2X1 U27003 ( .A(n25984), .B(n36261), .Y(n22796) );
  INVX1 U27004 ( .A(reg_file[2332]), .Y(n36261) );
  NOR2X1 U27005 ( .A(n25984), .B(n36262), .Y(n22795) );
  INVX1 U27006 ( .A(reg_file[2333]), .Y(n36262) );
  NOR2X1 U27007 ( .A(n25984), .B(n36263), .Y(n22794) );
  INVX1 U27008 ( .A(reg_file[2334]), .Y(n36263) );
  NOR2X1 U27009 ( .A(n25985), .B(n36264), .Y(n22793) );
  INVX1 U27010 ( .A(reg_file[2335]), .Y(n36264) );
  NOR2X1 U27011 ( .A(n25985), .B(n36265), .Y(n22792) );
  INVX1 U27012 ( .A(reg_file[2336]), .Y(n36265) );
  NOR2X1 U27013 ( .A(n25985), .B(n36266), .Y(n22791) );
  INVX1 U27014 ( .A(reg_file[2337]), .Y(n36266) );
  NOR2X1 U27015 ( .A(n25985), .B(n36267), .Y(n22790) );
  INVX1 U27016 ( .A(reg_file[2338]), .Y(n36267) );
  NOR2X1 U27017 ( .A(n25985), .B(n36268), .Y(n22789) );
  INVX1 U27018 ( .A(reg_file[2339]), .Y(n36268) );
  NOR2X1 U27019 ( .A(n25985), .B(n36269), .Y(n22788) );
  INVX1 U27020 ( .A(reg_file[2340]), .Y(n36269) );
  NOR2X1 U27021 ( .A(n25985), .B(n36270), .Y(n22787) );
  INVX1 U27022 ( .A(reg_file[2341]), .Y(n36270) );
  NOR2X1 U27023 ( .A(n25985), .B(n36271), .Y(n22786) );
  INVX1 U27024 ( .A(reg_file[2342]), .Y(n36271) );
  NOR2X1 U27025 ( .A(n25985), .B(n36272), .Y(n22785) );
  INVX1 U27026 ( .A(reg_file[2343]), .Y(n36272) );
  NOR2X1 U27027 ( .A(n25985), .B(n36273), .Y(n22784) );
  INVX1 U27028 ( .A(reg_file[2344]), .Y(n36273) );
  NOR2X1 U27029 ( .A(n25985), .B(n36274), .Y(n22783) );
  INVX1 U27030 ( .A(reg_file[2345]), .Y(n36274) );
  NOR2X1 U27031 ( .A(n25985), .B(n36275), .Y(n22782) );
  INVX1 U27032 ( .A(reg_file[2346]), .Y(n36275) );
  NOR2X1 U27033 ( .A(n25985), .B(n36276), .Y(n22781) );
  INVX1 U27034 ( .A(reg_file[2347]), .Y(n36276) );
  NOR2X1 U27035 ( .A(n25985), .B(n36277), .Y(n22780) );
  INVX1 U27036 ( .A(reg_file[2348]), .Y(n36277) );
  NOR2X1 U27037 ( .A(n25985), .B(n36278), .Y(n22779) );
  INVX1 U27038 ( .A(reg_file[2349]), .Y(n36278) );
  NOR2X1 U27039 ( .A(n25985), .B(n36279), .Y(n22778) );
  INVX1 U27040 ( .A(reg_file[2350]), .Y(n36279) );
  NOR2X1 U27041 ( .A(n25985), .B(n36280), .Y(n22777) );
  INVX1 U27042 ( .A(reg_file[2351]), .Y(n36280) );
  NOR2X1 U27043 ( .A(n25986), .B(n36281), .Y(n22776) );
  INVX1 U27044 ( .A(reg_file[2352]), .Y(n36281) );
  NOR2X1 U27045 ( .A(n25986), .B(n36282), .Y(n22775) );
  INVX1 U27046 ( .A(reg_file[2353]), .Y(n36282) );
  NOR2X1 U27047 ( .A(n25986), .B(n36283), .Y(n22774) );
  INVX1 U27048 ( .A(reg_file[2354]), .Y(n36283) );
  NOR2X1 U27049 ( .A(n25986), .B(n36284), .Y(n22773) );
  INVX1 U27050 ( .A(reg_file[2355]), .Y(n36284) );
  NOR2X1 U27051 ( .A(n25986), .B(n36285), .Y(n22772) );
  INVX1 U27052 ( .A(reg_file[2356]), .Y(n36285) );
  NOR2X1 U27053 ( .A(n25986), .B(n36286), .Y(n22771) );
  INVX1 U27054 ( .A(reg_file[2357]), .Y(n36286) );
  NOR2X1 U27055 ( .A(n25986), .B(n36287), .Y(n22770) );
  INVX1 U27056 ( .A(reg_file[2358]), .Y(n36287) );
  NOR2X1 U27057 ( .A(n25986), .B(n36288), .Y(n22769) );
  INVX1 U27058 ( .A(reg_file[2359]), .Y(n36288) );
  NOR2X1 U27059 ( .A(n25986), .B(n36289), .Y(n22768) );
  INVX1 U27060 ( .A(reg_file[2360]), .Y(n36289) );
  NOR2X1 U27061 ( .A(n25986), .B(n36290), .Y(n22767) );
  INVX1 U27062 ( .A(reg_file[2361]), .Y(n36290) );
  NOR2X1 U27063 ( .A(n25986), .B(n36291), .Y(n22766) );
  INVX1 U27064 ( .A(reg_file[2362]), .Y(n36291) );
  NOR2X1 U27065 ( .A(n25986), .B(n36292), .Y(n22765) );
  INVX1 U27066 ( .A(reg_file[2363]), .Y(n36292) );
  NOR2X1 U27067 ( .A(n25986), .B(n36293), .Y(n22764) );
  INVX1 U27068 ( .A(reg_file[2364]), .Y(n36293) );
  NOR2X1 U27069 ( .A(n25986), .B(n36294), .Y(n22763) );
  INVX1 U27070 ( .A(reg_file[2365]), .Y(n36294) );
  NOR2X1 U27071 ( .A(n25986), .B(n36295), .Y(n22762) );
  INVX1 U27072 ( .A(reg_file[2366]), .Y(n36295) );
  NOR2X1 U27073 ( .A(n25986), .B(n36296), .Y(n22761) );
  INVX1 U27074 ( .A(reg_file[2367]), .Y(n36296) );
  NOR2X1 U27075 ( .A(n25986), .B(n36297), .Y(n22760) );
  INVX1 U27076 ( .A(reg_file[2368]), .Y(n36297) );
  NOR2X1 U27077 ( .A(n25987), .B(n36298), .Y(n22759) );
  INVX1 U27078 ( .A(reg_file[2369]), .Y(n36298) );
  NOR2X1 U27079 ( .A(n25987), .B(n36299), .Y(n22758) );
  INVX1 U27080 ( .A(reg_file[2370]), .Y(n36299) );
  NOR2X1 U27081 ( .A(n25987), .B(n36300), .Y(n22757) );
  INVX1 U27082 ( .A(reg_file[2371]), .Y(n36300) );
  NOR2X1 U27083 ( .A(n25987), .B(n36301), .Y(n22756) );
  INVX1 U27084 ( .A(reg_file[2372]), .Y(n36301) );
  NOR2X1 U27085 ( .A(n25987), .B(n36302), .Y(n22755) );
  INVX1 U27086 ( .A(reg_file[2373]), .Y(n36302) );
  NOR2X1 U27087 ( .A(n25987), .B(n36303), .Y(n22754) );
  INVX1 U27088 ( .A(reg_file[2374]), .Y(n36303) );
  NOR2X1 U27089 ( .A(n25987), .B(n36304), .Y(n22753) );
  INVX1 U27090 ( .A(reg_file[2375]), .Y(n36304) );
  NOR2X1 U27091 ( .A(n25987), .B(n36305), .Y(n22752) );
  INVX1 U27092 ( .A(reg_file[2376]), .Y(n36305) );
  NOR2X1 U27093 ( .A(n25987), .B(n36306), .Y(n22751) );
  INVX1 U27094 ( .A(reg_file[2377]), .Y(n36306) );
  NOR2X1 U27095 ( .A(n25987), .B(n36307), .Y(n22750) );
  INVX1 U27096 ( .A(reg_file[2378]), .Y(n36307) );
  NOR2X1 U27097 ( .A(n25987), .B(n36308), .Y(n22749) );
  INVX1 U27098 ( .A(reg_file[2379]), .Y(n36308) );
  NOR2X1 U27099 ( .A(n25987), .B(n36309), .Y(n22748) );
  INVX1 U27100 ( .A(reg_file[2380]), .Y(n36309) );
  NOR2X1 U27101 ( .A(n25987), .B(n36310), .Y(n22747) );
  INVX1 U27102 ( .A(reg_file[2381]), .Y(n36310) );
  NOR2X1 U27103 ( .A(n25987), .B(n36311), .Y(n22746) );
  INVX1 U27104 ( .A(reg_file[2382]), .Y(n36311) );
  NOR2X1 U27105 ( .A(n25987), .B(n36312), .Y(n22745) );
  INVX1 U27106 ( .A(reg_file[2383]), .Y(n36312) );
  NOR2X1 U27107 ( .A(n25987), .B(n36313), .Y(n22744) );
  INVX1 U27108 ( .A(reg_file[2384]), .Y(n36313) );
  NOR2X1 U27109 ( .A(n25987), .B(n36314), .Y(n22743) );
  INVX1 U27110 ( .A(reg_file[2385]), .Y(n36314) );
  NOR2X1 U27111 ( .A(n25988), .B(n36315), .Y(n22742) );
  INVX1 U27112 ( .A(reg_file[2386]), .Y(n36315) );
  NOR2X1 U27113 ( .A(n25988), .B(n36316), .Y(n22741) );
  INVX1 U27114 ( .A(reg_file[2387]), .Y(n36316) );
  NOR2X1 U27115 ( .A(n25988), .B(n36317), .Y(n22740) );
  INVX1 U27116 ( .A(reg_file[2388]), .Y(n36317) );
  NOR2X1 U27117 ( .A(n25988), .B(n36318), .Y(n22739) );
  INVX1 U27118 ( .A(reg_file[2389]), .Y(n36318) );
  NOR2X1 U27119 ( .A(n25988), .B(n36319), .Y(n22738) );
  INVX1 U27120 ( .A(reg_file[2390]), .Y(n36319) );
  NOR2X1 U27121 ( .A(n25988), .B(n36320), .Y(n22737) );
  INVX1 U27122 ( .A(reg_file[2391]), .Y(n36320) );
  NOR2X1 U27123 ( .A(n25988), .B(n36321), .Y(n22736) );
  INVX1 U27124 ( .A(reg_file[2392]), .Y(n36321) );
  NOR2X1 U27125 ( .A(n25988), .B(n36322), .Y(n22735) );
  INVX1 U27126 ( .A(reg_file[2393]), .Y(n36322) );
  NOR2X1 U27127 ( .A(n25988), .B(n36323), .Y(n22734) );
  INVX1 U27128 ( .A(reg_file[2394]), .Y(n36323) );
  NOR2X1 U27129 ( .A(n25988), .B(n36324), .Y(n22733) );
  INVX1 U27130 ( .A(reg_file[2395]), .Y(n36324) );
  NOR2X1 U27131 ( .A(n25988), .B(n36325), .Y(n22732) );
  INVX1 U27132 ( .A(reg_file[2396]), .Y(n36325) );
  NOR2X1 U27133 ( .A(n25988), .B(n36326), .Y(n22731) );
  INVX1 U27134 ( .A(reg_file[2397]), .Y(n36326) );
  NOR2X1 U27135 ( .A(n25988), .B(n36327), .Y(n22730) );
  INVX1 U27136 ( .A(reg_file[2398]), .Y(n36327) );
  NOR2X1 U27137 ( .A(n25988), .B(n36328), .Y(n22729) );
  INVX1 U27138 ( .A(reg_file[2399]), .Y(n36328) );
  NOR2X1 U27139 ( .A(n25988), .B(n36329), .Y(n22728) );
  INVX1 U27140 ( .A(reg_file[2400]), .Y(n36329) );
  NOR2X1 U27141 ( .A(n25988), .B(n36330), .Y(n22727) );
  INVX1 U27142 ( .A(reg_file[2401]), .Y(n36330) );
  NOR2X1 U27143 ( .A(n25988), .B(n36331), .Y(n22726) );
  INVX1 U27144 ( .A(reg_file[2402]), .Y(n36331) );
  NOR2X1 U27145 ( .A(n25989), .B(n36332), .Y(n22725) );
  INVX1 U27146 ( .A(reg_file[2403]), .Y(n36332) );
  NOR2X1 U27147 ( .A(n25989), .B(n36333), .Y(n22724) );
  INVX1 U27148 ( .A(reg_file[2404]), .Y(n36333) );
  NOR2X1 U27149 ( .A(n25989), .B(n36334), .Y(n22723) );
  INVX1 U27150 ( .A(reg_file[2405]), .Y(n36334) );
  NOR2X1 U27151 ( .A(n25989), .B(n36335), .Y(n22722) );
  INVX1 U27152 ( .A(reg_file[2406]), .Y(n36335) );
  NOR2X1 U27153 ( .A(n25989), .B(n36336), .Y(n22721) );
  INVX1 U27154 ( .A(reg_file[2407]), .Y(n36336) );
  NOR2X1 U27155 ( .A(n25989), .B(n36337), .Y(n22720) );
  INVX1 U27156 ( .A(reg_file[2408]), .Y(n36337) );
  NOR2X1 U27157 ( .A(n25989), .B(n36338), .Y(n22719) );
  INVX1 U27158 ( .A(reg_file[2409]), .Y(n36338) );
  NOR2X1 U27159 ( .A(n25989), .B(n36339), .Y(n22718) );
  INVX1 U27160 ( .A(reg_file[2410]), .Y(n36339) );
  NOR2X1 U27161 ( .A(n25989), .B(n36340), .Y(n22717) );
  INVX1 U27162 ( .A(reg_file[2411]), .Y(n36340) );
  NOR2X1 U27163 ( .A(n25989), .B(n36341), .Y(n22716) );
  INVX1 U27164 ( .A(reg_file[2412]), .Y(n36341) );
  NOR2X1 U27165 ( .A(n25989), .B(n36342), .Y(n22715) );
  INVX1 U27166 ( .A(reg_file[2413]), .Y(n36342) );
  NOR2X1 U27167 ( .A(n25989), .B(n36343), .Y(n22714) );
  INVX1 U27168 ( .A(reg_file[2414]), .Y(n36343) );
  NOR2X1 U27169 ( .A(n25989), .B(n36344), .Y(n22713) );
  INVX1 U27170 ( .A(reg_file[2415]), .Y(n36344) );
  NOR2X1 U27171 ( .A(n25989), .B(n36345), .Y(n22712) );
  INVX1 U27172 ( .A(reg_file[2416]), .Y(n36345) );
  NOR2X1 U27173 ( .A(n25989), .B(n36346), .Y(n22711) );
  INVX1 U27174 ( .A(reg_file[2417]), .Y(n36346) );
  NOR2X1 U27175 ( .A(n25989), .B(n36347), .Y(n22710) );
  INVX1 U27176 ( .A(reg_file[2418]), .Y(n36347) );
  NOR2X1 U27177 ( .A(n25989), .B(n36348), .Y(n22709) );
  INVX1 U27178 ( .A(reg_file[2419]), .Y(n36348) );
  NOR2X1 U27179 ( .A(n25990), .B(n36349), .Y(n22708) );
  INVX1 U27180 ( .A(reg_file[2420]), .Y(n36349) );
  NOR2X1 U27181 ( .A(n25990), .B(n36350), .Y(n22707) );
  INVX1 U27182 ( .A(reg_file[2421]), .Y(n36350) );
  NOR2X1 U27183 ( .A(n25990), .B(n36351), .Y(n22706) );
  INVX1 U27184 ( .A(reg_file[2422]), .Y(n36351) );
  NOR2X1 U27185 ( .A(n25990), .B(n36352), .Y(n22705) );
  INVX1 U27186 ( .A(reg_file[2423]), .Y(n36352) );
  NOR2X1 U27187 ( .A(n25990), .B(n36353), .Y(n22704) );
  INVX1 U27188 ( .A(reg_file[2424]), .Y(n36353) );
  NOR2X1 U27189 ( .A(n25990), .B(n36354), .Y(n22703) );
  INVX1 U27190 ( .A(reg_file[2425]), .Y(n36354) );
  NOR2X1 U27191 ( .A(n25990), .B(n36355), .Y(n22702) );
  INVX1 U27192 ( .A(reg_file[2426]), .Y(n36355) );
  NOR2X1 U27193 ( .A(n25990), .B(n36356), .Y(n22701) );
  INVX1 U27194 ( .A(reg_file[2427]), .Y(n36356) );
  NOR2X1 U27195 ( .A(n25990), .B(n36357), .Y(n22700) );
  INVX1 U27196 ( .A(reg_file[2428]), .Y(n36357) );
  NOR2X1 U27197 ( .A(n25990), .B(n36358), .Y(n22699) );
  INVX1 U27198 ( .A(reg_file[2429]), .Y(n36358) );
  NOR2X1 U27199 ( .A(n25990), .B(n36359), .Y(n22698) );
  INVX1 U27200 ( .A(reg_file[2430]), .Y(n36359) );
  NOR2X1 U27201 ( .A(n25990), .B(n36360), .Y(n22697) );
  INVX1 U27202 ( .A(reg_file[2431]), .Y(n36360) );
  NOR2X1 U27203 ( .A(n36101), .B(n34927), .Y(n36233) );
  MUX2X1 U27204 ( .B(n36361), .A(n25129), .S(n25991), .Y(n22696) );
  INVX1 U27205 ( .A(reg_file[2432]), .Y(n36361) );
  MUX2X1 U27206 ( .B(n36363), .A(n25130), .S(n25991), .Y(n22695) );
  INVX1 U27207 ( .A(reg_file[2433]), .Y(n36363) );
  MUX2X1 U27208 ( .B(n36364), .A(n25131), .S(n25991), .Y(n22694) );
  INVX1 U27209 ( .A(reg_file[2434]), .Y(n36364) );
  MUX2X1 U27210 ( .B(n36365), .A(n25132), .S(n25991), .Y(n22693) );
  INVX1 U27211 ( .A(reg_file[2435]), .Y(n36365) );
  MUX2X1 U27212 ( .B(n36366), .A(n25133), .S(n25991), .Y(n22692) );
  INVX1 U27213 ( .A(reg_file[2436]), .Y(n36366) );
  MUX2X1 U27214 ( .B(n36367), .A(n25134), .S(n25991), .Y(n22691) );
  INVX1 U27215 ( .A(reg_file[2437]), .Y(n36367) );
  MUX2X1 U27216 ( .B(n36368), .A(n25135), .S(n25991), .Y(n22690) );
  INVX1 U27217 ( .A(reg_file[2438]), .Y(n36368) );
  MUX2X1 U27218 ( .B(n36369), .A(n25136), .S(n25991), .Y(n22689) );
  INVX1 U27219 ( .A(reg_file[2439]), .Y(n36369) );
  NOR2X1 U27220 ( .A(n25991), .B(n36370), .Y(n22688) );
  INVX1 U27221 ( .A(reg_file[2440]), .Y(n36370) );
  NOR2X1 U27222 ( .A(n25991), .B(n36371), .Y(n22687) );
  INVX1 U27223 ( .A(reg_file[2441]), .Y(n36371) );
  NOR2X1 U27224 ( .A(n25991), .B(n36372), .Y(n22686) );
  INVX1 U27225 ( .A(reg_file[2442]), .Y(n36372) );
  NOR2X1 U27226 ( .A(n25991), .B(n36373), .Y(n22685) );
  INVX1 U27227 ( .A(reg_file[2443]), .Y(n36373) );
  NOR2X1 U27228 ( .A(n25991), .B(n36374), .Y(n22684) );
  INVX1 U27229 ( .A(reg_file[2444]), .Y(n36374) );
  NOR2X1 U27230 ( .A(n25991), .B(n36375), .Y(n22683) );
  INVX1 U27231 ( .A(reg_file[2445]), .Y(n36375) );
  NOR2X1 U27232 ( .A(n25992), .B(n36376), .Y(n22682) );
  INVX1 U27233 ( .A(reg_file[2446]), .Y(n36376) );
  NOR2X1 U27234 ( .A(n25992), .B(n36377), .Y(n22681) );
  INVX1 U27235 ( .A(reg_file[2447]), .Y(n36377) );
  NOR2X1 U27236 ( .A(n25992), .B(n36378), .Y(n22680) );
  INVX1 U27237 ( .A(reg_file[2448]), .Y(n36378) );
  NOR2X1 U27238 ( .A(n25992), .B(n36379), .Y(n22679) );
  INVX1 U27239 ( .A(reg_file[2449]), .Y(n36379) );
  NOR2X1 U27240 ( .A(n25992), .B(n36380), .Y(n22678) );
  INVX1 U27241 ( .A(reg_file[2450]), .Y(n36380) );
  NOR2X1 U27242 ( .A(n25992), .B(n36381), .Y(n22677) );
  INVX1 U27243 ( .A(reg_file[2451]), .Y(n36381) );
  NOR2X1 U27244 ( .A(n25992), .B(n36382), .Y(n22676) );
  INVX1 U27245 ( .A(reg_file[2452]), .Y(n36382) );
  NOR2X1 U27246 ( .A(n25992), .B(n36383), .Y(n22675) );
  INVX1 U27247 ( .A(reg_file[2453]), .Y(n36383) );
  NOR2X1 U27248 ( .A(n25992), .B(n36384), .Y(n22674) );
  INVX1 U27249 ( .A(reg_file[2454]), .Y(n36384) );
  NOR2X1 U27250 ( .A(n25992), .B(n36385), .Y(n22673) );
  INVX1 U27251 ( .A(reg_file[2455]), .Y(n36385) );
  NOR2X1 U27252 ( .A(n25992), .B(n36386), .Y(n22672) );
  INVX1 U27253 ( .A(reg_file[2456]), .Y(n36386) );
  NOR2X1 U27254 ( .A(n25992), .B(n36387), .Y(n22671) );
  INVX1 U27255 ( .A(reg_file[2457]), .Y(n36387) );
  NOR2X1 U27256 ( .A(n25992), .B(n36388), .Y(n22670) );
  INVX1 U27257 ( .A(reg_file[2458]), .Y(n36388) );
  NOR2X1 U27258 ( .A(n25992), .B(n36389), .Y(n22669) );
  INVX1 U27259 ( .A(reg_file[2459]), .Y(n36389) );
  NOR2X1 U27260 ( .A(n25992), .B(n36390), .Y(n22668) );
  INVX1 U27261 ( .A(reg_file[2460]), .Y(n36390) );
  NOR2X1 U27262 ( .A(n25992), .B(n36391), .Y(n22667) );
  INVX1 U27263 ( .A(reg_file[2461]), .Y(n36391) );
  NOR2X1 U27264 ( .A(n25992), .B(n36392), .Y(n22666) );
  INVX1 U27265 ( .A(reg_file[2462]), .Y(n36392) );
  NOR2X1 U27266 ( .A(n25993), .B(n36393), .Y(n22665) );
  INVX1 U27267 ( .A(reg_file[2463]), .Y(n36393) );
  NOR2X1 U27268 ( .A(n25993), .B(n36394), .Y(n22664) );
  INVX1 U27269 ( .A(reg_file[2464]), .Y(n36394) );
  NOR2X1 U27270 ( .A(n25993), .B(n36395), .Y(n22663) );
  INVX1 U27271 ( .A(reg_file[2465]), .Y(n36395) );
  NOR2X1 U27272 ( .A(n25993), .B(n36396), .Y(n22662) );
  INVX1 U27273 ( .A(reg_file[2466]), .Y(n36396) );
  NOR2X1 U27274 ( .A(n25993), .B(n36397), .Y(n22661) );
  INVX1 U27275 ( .A(reg_file[2467]), .Y(n36397) );
  NOR2X1 U27276 ( .A(n25993), .B(n36398), .Y(n22660) );
  INVX1 U27277 ( .A(reg_file[2468]), .Y(n36398) );
  NOR2X1 U27278 ( .A(n25993), .B(n36399), .Y(n22659) );
  INVX1 U27279 ( .A(reg_file[2469]), .Y(n36399) );
  NOR2X1 U27280 ( .A(n25993), .B(n36400), .Y(n22658) );
  INVX1 U27281 ( .A(reg_file[2470]), .Y(n36400) );
  NOR2X1 U27282 ( .A(n25993), .B(n36401), .Y(n22657) );
  INVX1 U27283 ( .A(reg_file[2471]), .Y(n36401) );
  NOR2X1 U27284 ( .A(n25993), .B(n36402), .Y(n22656) );
  INVX1 U27285 ( .A(reg_file[2472]), .Y(n36402) );
  NOR2X1 U27286 ( .A(n25993), .B(n36403), .Y(n22655) );
  INVX1 U27287 ( .A(reg_file[2473]), .Y(n36403) );
  NOR2X1 U27288 ( .A(n25993), .B(n36404), .Y(n22654) );
  INVX1 U27289 ( .A(reg_file[2474]), .Y(n36404) );
  NOR2X1 U27290 ( .A(n25993), .B(n36405), .Y(n22653) );
  INVX1 U27291 ( .A(reg_file[2475]), .Y(n36405) );
  NOR2X1 U27292 ( .A(n25993), .B(n36406), .Y(n22652) );
  INVX1 U27293 ( .A(reg_file[2476]), .Y(n36406) );
  NOR2X1 U27294 ( .A(n25993), .B(n36407), .Y(n22651) );
  INVX1 U27295 ( .A(reg_file[2477]), .Y(n36407) );
  NOR2X1 U27296 ( .A(n25993), .B(n36408), .Y(n22650) );
  INVX1 U27297 ( .A(reg_file[2478]), .Y(n36408) );
  NOR2X1 U27298 ( .A(n25993), .B(n36409), .Y(n22649) );
  INVX1 U27299 ( .A(reg_file[2479]), .Y(n36409) );
  NOR2X1 U27300 ( .A(n25994), .B(n36410), .Y(n22648) );
  INVX1 U27301 ( .A(reg_file[2480]), .Y(n36410) );
  NOR2X1 U27302 ( .A(n25994), .B(n36411), .Y(n22647) );
  INVX1 U27303 ( .A(reg_file[2481]), .Y(n36411) );
  NOR2X1 U27304 ( .A(n25994), .B(n36412), .Y(n22646) );
  INVX1 U27305 ( .A(reg_file[2482]), .Y(n36412) );
  NOR2X1 U27306 ( .A(n25994), .B(n36413), .Y(n22645) );
  INVX1 U27307 ( .A(reg_file[2483]), .Y(n36413) );
  NOR2X1 U27308 ( .A(n25994), .B(n36414), .Y(n22644) );
  INVX1 U27309 ( .A(reg_file[2484]), .Y(n36414) );
  NOR2X1 U27310 ( .A(n25994), .B(n36415), .Y(n22643) );
  INVX1 U27311 ( .A(reg_file[2485]), .Y(n36415) );
  NOR2X1 U27312 ( .A(n25994), .B(n36416), .Y(n22642) );
  INVX1 U27313 ( .A(reg_file[2486]), .Y(n36416) );
  NOR2X1 U27314 ( .A(n25994), .B(n36417), .Y(n22641) );
  INVX1 U27315 ( .A(reg_file[2487]), .Y(n36417) );
  NOR2X1 U27316 ( .A(n25994), .B(n36418), .Y(n22640) );
  INVX1 U27317 ( .A(reg_file[2488]), .Y(n36418) );
  NOR2X1 U27318 ( .A(n25994), .B(n36419), .Y(n22639) );
  INVX1 U27319 ( .A(reg_file[2489]), .Y(n36419) );
  NOR2X1 U27320 ( .A(n25994), .B(n36420), .Y(n22638) );
  INVX1 U27321 ( .A(reg_file[2490]), .Y(n36420) );
  NOR2X1 U27322 ( .A(n25994), .B(n36421), .Y(n22637) );
  INVX1 U27323 ( .A(reg_file[2491]), .Y(n36421) );
  NOR2X1 U27324 ( .A(n25994), .B(n36422), .Y(n22636) );
  INVX1 U27325 ( .A(reg_file[2492]), .Y(n36422) );
  NOR2X1 U27326 ( .A(n25994), .B(n36423), .Y(n22635) );
  INVX1 U27327 ( .A(reg_file[2493]), .Y(n36423) );
  NOR2X1 U27328 ( .A(n25994), .B(n36424), .Y(n22634) );
  INVX1 U27329 ( .A(reg_file[2494]), .Y(n36424) );
  NOR2X1 U27330 ( .A(n25994), .B(n36425), .Y(n22633) );
  INVX1 U27331 ( .A(reg_file[2495]), .Y(n36425) );
  NOR2X1 U27332 ( .A(n25994), .B(n36426), .Y(n22632) );
  INVX1 U27333 ( .A(reg_file[2496]), .Y(n36426) );
  NOR2X1 U27334 ( .A(n25995), .B(n36427), .Y(n22631) );
  INVX1 U27335 ( .A(reg_file[2497]), .Y(n36427) );
  NOR2X1 U27336 ( .A(n25995), .B(n36428), .Y(n22630) );
  INVX1 U27337 ( .A(reg_file[2498]), .Y(n36428) );
  NOR2X1 U27338 ( .A(n25995), .B(n36429), .Y(n22629) );
  INVX1 U27339 ( .A(reg_file[2499]), .Y(n36429) );
  NOR2X1 U27340 ( .A(n25995), .B(n36430), .Y(n22628) );
  INVX1 U27341 ( .A(reg_file[2500]), .Y(n36430) );
  NOR2X1 U27342 ( .A(n25995), .B(n36431), .Y(n22627) );
  INVX1 U27343 ( .A(reg_file[2501]), .Y(n36431) );
  NOR2X1 U27344 ( .A(n25995), .B(n36432), .Y(n22626) );
  INVX1 U27345 ( .A(reg_file[2502]), .Y(n36432) );
  NOR2X1 U27346 ( .A(n25995), .B(n36433), .Y(n22625) );
  INVX1 U27347 ( .A(reg_file[2503]), .Y(n36433) );
  NOR2X1 U27348 ( .A(n25995), .B(n36434), .Y(n22624) );
  INVX1 U27349 ( .A(reg_file[2504]), .Y(n36434) );
  NOR2X1 U27350 ( .A(n25995), .B(n36435), .Y(n22623) );
  INVX1 U27351 ( .A(reg_file[2505]), .Y(n36435) );
  NOR2X1 U27352 ( .A(n25995), .B(n36436), .Y(n22622) );
  INVX1 U27353 ( .A(reg_file[2506]), .Y(n36436) );
  NOR2X1 U27354 ( .A(n25995), .B(n36437), .Y(n22621) );
  INVX1 U27355 ( .A(reg_file[2507]), .Y(n36437) );
  NOR2X1 U27356 ( .A(n25995), .B(n36438), .Y(n22620) );
  INVX1 U27357 ( .A(reg_file[2508]), .Y(n36438) );
  NOR2X1 U27358 ( .A(n25995), .B(n36439), .Y(n22619) );
  INVX1 U27359 ( .A(reg_file[2509]), .Y(n36439) );
  NOR2X1 U27360 ( .A(n25995), .B(n36440), .Y(n22618) );
  INVX1 U27361 ( .A(reg_file[2510]), .Y(n36440) );
  NOR2X1 U27362 ( .A(n25995), .B(n36441), .Y(n22617) );
  INVX1 U27363 ( .A(reg_file[2511]), .Y(n36441) );
  NOR2X1 U27364 ( .A(n25995), .B(n36442), .Y(n22616) );
  INVX1 U27365 ( .A(reg_file[2512]), .Y(n36442) );
  NOR2X1 U27366 ( .A(n25995), .B(n36443), .Y(n22615) );
  INVX1 U27367 ( .A(reg_file[2513]), .Y(n36443) );
  NOR2X1 U27368 ( .A(n25996), .B(n36444), .Y(n22614) );
  INVX1 U27369 ( .A(reg_file[2514]), .Y(n36444) );
  NOR2X1 U27370 ( .A(n25996), .B(n36445), .Y(n22613) );
  INVX1 U27371 ( .A(reg_file[2515]), .Y(n36445) );
  NOR2X1 U27372 ( .A(n25996), .B(n36446), .Y(n22612) );
  INVX1 U27373 ( .A(reg_file[2516]), .Y(n36446) );
  NOR2X1 U27374 ( .A(n25996), .B(n36447), .Y(n22611) );
  INVX1 U27375 ( .A(reg_file[2517]), .Y(n36447) );
  NOR2X1 U27376 ( .A(n25996), .B(n36448), .Y(n22610) );
  INVX1 U27377 ( .A(reg_file[2518]), .Y(n36448) );
  NOR2X1 U27378 ( .A(n25996), .B(n36449), .Y(n22609) );
  INVX1 U27379 ( .A(reg_file[2519]), .Y(n36449) );
  NOR2X1 U27380 ( .A(n25996), .B(n36450), .Y(n22608) );
  INVX1 U27381 ( .A(reg_file[2520]), .Y(n36450) );
  NOR2X1 U27382 ( .A(n25996), .B(n36451), .Y(n22607) );
  INVX1 U27383 ( .A(reg_file[2521]), .Y(n36451) );
  NOR2X1 U27384 ( .A(n25996), .B(n36452), .Y(n22606) );
  INVX1 U27385 ( .A(reg_file[2522]), .Y(n36452) );
  NOR2X1 U27386 ( .A(n25996), .B(n36453), .Y(n22605) );
  INVX1 U27387 ( .A(reg_file[2523]), .Y(n36453) );
  NOR2X1 U27388 ( .A(n25996), .B(n36454), .Y(n22604) );
  INVX1 U27389 ( .A(reg_file[2524]), .Y(n36454) );
  NOR2X1 U27390 ( .A(n25996), .B(n36455), .Y(n22603) );
  INVX1 U27391 ( .A(reg_file[2525]), .Y(n36455) );
  NOR2X1 U27392 ( .A(n25996), .B(n36456), .Y(n22602) );
  INVX1 U27393 ( .A(reg_file[2526]), .Y(n36456) );
  NOR2X1 U27394 ( .A(n25996), .B(n36457), .Y(n22601) );
  INVX1 U27395 ( .A(reg_file[2527]), .Y(n36457) );
  NOR2X1 U27396 ( .A(n25996), .B(n36458), .Y(n22600) );
  INVX1 U27397 ( .A(reg_file[2528]), .Y(n36458) );
  NOR2X1 U27398 ( .A(n25996), .B(n36459), .Y(n22599) );
  INVX1 U27399 ( .A(reg_file[2529]), .Y(n36459) );
  NOR2X1 U27400 ( .A(n25996), .B(n36460), .Y(n22598) );
  INVX1 U27401 ( .A(reg_file[2530]), .Y(n36460) );
  NOR2X1 U27402 ( .A(n25997), .B(n36461), .Y(n22597) );
  INVX1 U27403 ( .A(reg_file[2531]), .Y(n36461) );
  NOR2X1 U27404 ( .A(n25997), .B(n36462), .Y(n22596) );
  INVX1 U27405 ( .A(reg_file[2532]), .Y(n36462) );
  NOR2X1 U27406 ( .A(n25997), .B(n36463), .Y(n22595) );
  INVX1 U27407 ( .A(reg_file[2533]), .Y(n36463) );
  NOR2X1 U27408 ( .A(n25997), .B(n36464), .Y(n22594) );
  INVX1 U27409 ( .A(reg_file[2534]), .Y(n36464) );
  NOR2X1 U27410 ( .A(n25997), .B(n36465), .Y(n22593) );
  INVX1 U27411 ( .A(reg_file[2535]), .Y(n36465) );
  NOR2X1 U27412 ( .A(n25997), .B(n36466), .Y(n22592) );
  INVX1 U27413 ( .A(reg_file[2536]), .Y(n36466) );
  NOR2X1 U27414 ( .A(n25997), .B(n36467), .Y(n22591) );
  INVX1 U27415 ( .A(reg_file[2537]), .Y(n36467) );
  NOR2X1 U27416 ( .A(n25997), .B(n36468), .Y(n22590) );
  INVX1 U27417 ( .A(reg_file[2538]), .Y(n36468) );
  NOR2X1 U27418 ( .A(n25997), .B(n36469), .Y(n22589) );
  INVX1 U27419 ( .A(reg_file[2539]), .Y(n36469) );
  NOR2X1 U27420 ( .A(n25997), .B(n36470), .Y(n22588) );
  INVX1 U27421 ( .A(reg_file[2540]), .Y(n36470) );
  NOR2X1 U27422 ( .A(n25997), .B(n36471), .Y(n22587) );
  INVX1 U27423 ( .A(reg_file[2541]), .Y(n36471) );
  NOR2X1 U27424 ( .A(n25997), .B(n36472), .Y(n22586) );
  INVX1 U27425 ( .A(reg_file[2542]), .Y(n36472) );
  NOR2X1 U27426 ( .A(n25997), .B(n36473), .Y(n22585) );
  INVX1 U27427 ( .A(reg_file[2543]), .Y(n36473) );
  NOR2X1 U27428 ( .A(n25997), .B(n36474), .Y(n22584) );
  INVX1 U27429 ( .A(reg_file[2544]), .Y(n36474) );
  NOR2X1 U27430 ( .A(n25997), .B(n36475), .Y(n22583) );
  INVX1 U27431 ( .A(reg_file[2545]), .Y(n36475) );
  NOR2X1 U27432 ( .A(n25997), .B(n36476), .Y(n22582) );
  INVX1 U27433 ( .A(reg_file[2546]), .Y(n36476) );
  NOR2X1 U27434 ( .A(n25997), .B(n36477), .Y(n22581) );
  INVX1 U27435 ( .A(reg_file[2547]), .Y(n36477) );
  NOR2X1 U27436 ( .A(n25998), .B(n36478), .Y(n22580) );
  INVX1 U27437 ( .A(reg_file[2548]), .Y(n36478) );
  NOR2X1 U27438 ( .A(n25998), .B(n36479), .Y(n22579) );
  INVX1 U27439 ( .A(reg_file[2549]), .Y(n36479) );
  NOR2X1 U27440 ( .A(n25998), .B(n36480), .Y(n22578) );
  INVX1 U27441 ( .A(reg_file[2550]), .Y(n36480) );
  NOR2X1 U27442 ( .A(n25998), .B(n36481), .Y(n22577) );
  INVX1 U27443 ( .A(reg_file[2551]), .Y(n36481) );
  NOR2X1 U27444 ( .A(n25998), .B(n36482), .Y(n22576) );
  INVX1 U27445 ( .A(reg_file[2552]), .Y(n36482) );
  NOR2X1 U27446 ( .A(n25998), .B(n36483), .Y(n22575) );
  INVX1 U27447 ( .A(reg_file[2553]), .Y(n36483) );
  NOR2X1 U27448 ( .A(n25998), .B(n36484), .Y(n22574) );
  INVX1 U27449 ( .A(reg_file[2554]), .Y(n36484) );
  NOR2X1 U27450 ( .A(n25998), .B(n36485), .Y(n22573) );
  INVX1 U27451 ( .A(reg_file[2555]), .Y(n36485) );
  NOR2X1 U27452 ( .A(n25998), .B(n36486), .Y(n22572) );
  INVX1 U27453 ( .A(reg_file[2556]), .Y(n36486) );
  NOR2X1 U27454 ( .A(n25998), .B(n36487), .Y(n22571) );
  INVX1 U27455 ( .A(reg_file[2557]), .Y(n36487) );
  NOR2X1 U27456 ( .A(n25998), .B(n36488), .Y(n22570) );
  INVX1 U27457 ( .A(reg_file[2558]), .Y(n36488) );
  NOR2X1 U27458 ( .A(n25998), .B(n36489), .Y(n22569) );
  INVX1 U27459 ( .A(reg_file[2559]), .Y(n36489) );
  NOR2X1 U27460 ( .A(n36231), .B(n34927), .Y(n36362) );
  MUX2X1 U27461 ( .B(n31519), .A(n25129), .S(n25999), .Y(n22568) );
  INVX1 U27462 ( .A(reg_file[2560]), .Y(n31519) );
  MUX2X1 U27463 ( .B(n29862), .A(n25130), .S(n25999), .Y(n22567) );
  INVX1 U27464 ( .A(reg_file[2561]), .Y(n29862) );
  MUX2X1 U27465 ( .B(n29400), .A(n25131), .S(n25999), .Y(n22566) );
  INVX1 U27466 ( .A(reg_file[2562]), .Y(n29400) );
  MUX2X1 U27467 ( .B(n28938), .A(n25132), .S(n25999), .Y(n22565) );
  INVX1 U27468 ( .A(reg_file[2563]), .Y(n28938) );
  MUX2X1 U27469 ( .B(n28476), .A(n25133), .S(n25999), .Y(n22564) );
  INVX1 U27470 ( .A(reg_file[2564]), .Y(n28476) );
  MUX2X1 U27471 ( .B(n28014), .A(n25134), .S(n25999), .Y(n22563) );
  INVX1 U27472 ( .A(reg_file[2565]), .Y(n28014) );
  MUX2X1 U27473 ( .B(n27552), .A(n25135), .S(n25999), .Y(n22562) );
  INVX1 U27474 ( .A(reg_file[2566]), .Y(n27552) );
  MUX2X1 U27475 ( .B(n27090), .A(n25136), .S(n25999), .Y(n22561) );
  INVX1 U27476 ( .A(reg_file[2567]), .Y(n27090) );
  NOR2X1 U27477 ( .A(n25999), .B(n26628), .Y(n22560) );
  INVX1 U27478 ( .A(reg_file[2568]), .Y(n26628) );
  NOR2X1 U27479 ( .A(n25999), .B(n26159), .Y(n22559) );
  INVX1 U27480 ( .A(reg_file[2569]), .Y(n26159) );
  NOR2X1 U27481 ( .A(n25999), .B(n31038), .Y(n22558) );
  INVX1 U27482 ( .A(reg_file[2570]), .Y(n31038) );
  NOR2X1 U27483 ( .A(n25999), .B(n30576), .Y(n22557) );
  INVX1 U27484 ( .A(reg_file[2571]), .Y(n30576) );
  NOR2X1 U27485 ( .A(n25999), .B(n30198), .Y(n22556) );
  INVX1 U27486 ( .A(reg_file[2572]), .Y(n30198) );
  NOR2X1 U27487 ( .A(n25999), .B(n30156), .Y(n22555) );
  INVX1 U27488 ( .A(reg_file[2573]), .Y(n30156) );
  NOR2X1 U27489 ( .A(n26000), .B(n30114), .Y(n22554) );
  INVX1 U27490 ( .A(reg_file[2574]), .Y(n30114) );
  NOR2X1 U27491 ( .A(n26000), .B(n30072), .Y(n22553) );
  INVX1 U27492 ( .A(reg_file[2575]), .Y(n30072) );
  NOR2X1 U27493 ( .A(n26000), .B(n30030), .Y(n22552) );
  INVX1 U27494 ( .A(reg_file[2576]), .Y(n30030) );
  NOR2X1 U27495 ( .A(n26000), .B(n29988), .Y(n22551) );
  INVX1 U27496 ( .A(reg_file[2577]), .Y(n29988) );
  NOR2X1 U27497 ( .A(n26000), .B(n29946), .Y(n22550) );
  INVX1 U27498 ( .A(reg_file[2578]), .Y(n29946) );
  NOR2X1 U27499 ( .A(n26000), .B(n29904), .Y(n22549) );
  INVX1 U27500 ( .A(reg_file[2579]), .Y(n29904) );
  NOR2X1 U27501 ( .A(n26000), .B(n29820), .Y(n22548) );
  INVX1 U27502 ( .A(reg_file[2580]), .Y(n29820) );
  NOR2X1 U27503 ( .A(n26000), .B(n29778), .Y(n22547) );
  INVX1 U27504 ( .A(reg_file[2581]), .Y(n29778) );
  NOR2X1 U27505 ( .A(n26000), .B(n29736), .Y(n22546) );
  INVX1 U27506 ( .A(reg_file[2582]), .Y(n29736) );
  NOR2X1 U27507 ( .A(n26000), .B(n29694), .Y(n22545) );
  INVX1 U27508 ( .A(reg_file[2583]), .Y(n29694) );
  NOR2X1 U27509 ( .A(n26000), .B(n29652), .Y(n22544) );
  INVX1 U27510 ( .A(reg_file[2584]), .Y(n29652) );
  NOR2X1 U27511 ( .A(n26000), .B(n29610), .Y(n22543) );
  INVX1 U27512 ( .A(reg_file[2585]), .Y(n29610) );
  NOR2X1 U27513 ( .A(n26000), .B(n29568), .Y(n22542) );
  INVX1 U27514 ( .A(reg_file[2586]), .Y(n29568) );
  NOR2X1 U27515 ( .A(n26000), .B(n29526), .Y(n22541) );
  INVX1 U27516 ( .A(reg_file[2587]), .Y(n29526) );
  NOR2X1 U27517 ( .A(n26000), .B(n29484), .Y(n22540) );
  INVX1 U27518 ( .A(reg_file[2588]), .Y(n29484) );
  NOR2X1 U27519 ( .A(n26000), .B(n29442), .Y(n22539) );
  INVX1 U27520 ( .A(reg_file[2589]), .Y(n29442) );
  NOR2X1 U27521 ( .A(n26000), .B(n29358), .Y(n22538) );
  INVX1 U27522 ( .A(reg_file[2590]), .Y(n29358) );
  NOR2X1 U27523 ( .A(n26001), .B(n29316), .Y(n22537) );
  INVX1 U27524 ( .A(reg_file[2591]), .Y(n29316) );
  NOR2X1 U27525 ( .A(n26001), .B(n29274), .Y(n22536) );
  INVX1 U27526 ( .A(reg_file[2592]), .Y(n29274) );
  NOR2X1 U27527 ( .A(n26001), .B(n29232), .Y(n22535) );
  INVX1 U27528 ( .A(reg_file[2593]), .Y(n29232) );
  NOR2X1 U27529 ( .A(n26001), .B(n29190), .Y(n22534) );
  INVX1 U27530 ( .A(reg_file[2594]), .Y(n29190) );
  NOR2X1 U27531 ( .A(n26001), .B(n29148), .Y(n22533) );
  INVX1 U27532 ( .A(reg_file[2595]), .Y(n29148) );
  NOR2X1 U27533 ( .A(n26001), .B(n29106), .Y(n22532) );
  INVX1 U27534 ( .A(reg_file[2596]), .Y(n29106) );
  NOR2X1 U27535 ( .A(n26001), .B(n29064), .Y(n22531) );
  INVX1 U27536 ( .A(reg_file[2597]), .Y(n29064) );
  NOR2X1 U27537 ( .A(n26001), .B(n29022), .Y(n22530) );
  INVX1 U27538 ( .A(reg_file[2598]), .Y(n29022) );
  NOR2X1 U27539 ( .A(n26001), .B(n28980), .Y(n22529) );
  INVX1 U27540 ( .A(reg_file[2599]), .Y(n28980) );
  NOR2X1 U27541 ( .A(n26001), .B(n28896), .Y(n22528) );
  INVX1 U27542 ( .A(reg_file[2600]), .Y(n28896) );
  NOR2X1 U27543 ( .A(n26001), .B(n28854), .Y(n22527) );
  INVX1 U27544 ( .A(reg_file[2601]), .Y(n28854) );
  NOR2X1 U27545 ( .A(n26001), .B(n28812), .Y(n22526) );
  INVX1 U27546 ( .A(reg_file[2602]), .Y(n28812) );
  NOR2X1 U27547 ( .A(n26001), .B(n28770), .Y(n22525) );
  INVX1 U27548 ( .A(reg_file[2603]), .Y(n28770) );
  NOR2X1 U27549 ( .A(n26001), .B(n28728), .Y(n22524) );
  INVX1 U27550 ( .A(reg_file[2604]), .Y(n28728) );
  NOR2X1 U27551 ( .A(n26001), .B(n28686), .Y(n22523) );
  INVX1 U27552 ( .A(reg_file[2605]), .Y(n28686) );
  NOR2X1 U27553 ( .A(n26001), .B(n28644), .Y(n22522) );
  INVX1 U27554 ( .A(reg_file[2606]), .Y(n28644) );
  NOR2X1 U27555 ( .A(n26001), .B(n28602), .Y(n22521) );
  INVX1 U27556 ( .A(reg_file[2607]), .Y(n28602) );
  NOR2X1 U27557 ( .A(n26002), .B(n28560), .Y(n22520) );
  INVX1 U27558 ( .A(reg_file[2608]), .Y(n28560) );
  NOR2X1 U27559 ( .A(n26002), .B(n28518), .Y(n22519) );
  INVX1 U27560 ( .A(reg_file[2609]), .Y(n28518) );
  NOR2X1 U27561 ( .A(n26002), .B(n28434), .Y(n22518) );
  INVX1 U27562 ( .A(reg_file[2610]), .Y(n28434) );
  NOR2X1 U27563 ( .A(n26002), .B(n28392), .Y(n22517) );
  INVX1 U27564 ( .A(reg_file[2611]), .Y(n28392) );
  NOR2X1 U27565 ( .A(n26002), .B(n28350), .Y(n22516) );
  INVX1 U27566 ( .A(reg_file[2612]), .Y(n28350) );
  NOR2X1 U27567 ( .A(n26002), .B(n28308), .Y(n22515) );
  INVX1 U27568 ( .A(reg_file[2613]), .Y(n28308) );
  NOR2X1 U27569 ( .A(n26002), .B(n28266), .Y(n22514) );
  INVX1 U27570 ( .A(reg_file[2614]), .Y(n28266) );
  NOR2X1 U27571 ( .A(n26002), .B(n28224), .Y(n22513) );
  INVX1 U27572 ( .A(reg_file[2615]), .Y(n28224) );
  NOR2X1 U27573 ( .A(n26002), .B(n28182), .Y(n22512) );
  INVX1 U27574 ( .A(reg_file[2616]), .Y(n28182) );
  NOR2X1 U27575 ( .A(n26002), .B(n28140), .Y(n22511) );
  INVX1 U27576 ( .A(reg_file[2617]), .Y(n28140) );
  NOR2X1 U27577 ( .A(n26002), .B(n28098), .Y(n22510) );
  INVX1 U27578 ( .A(reg_file[2618]), .Y(n28098) );
  NOR2X1 U27579 ( .A(n26002), .B(n28056), .Y(n22509) );
  INVX1 U27580 ( .A(reg_file[2619]), .Y(n28056) );
  NOR2X1 U27581 ( .A(n26002), .B(n27972), .Y(n22508) );
  INVX1 U27582 ( .A(reg_file[2620]), .Y(n27972) );
  NOR2X1 U27583 ( .A(n26002), .B(n27930), .Y(n22507) );
  INVX1 U27584 ( .A(reg_file[2621]), .Y(n27930) );
  NOR2X1 U27585 ( .A(n26002), .B(n27888), .Y(n22506) );
  INVX1 U27586 ( .A(reg_file[2622]), .Y(n27888) );
  NOR2X1 U27587 ( .A(n26002), .B(n27846), .Y(n22505) );
  INVX1 U27588 ( .A(reg_file[2623]), .Y(n27846) );
  NOR2X1 U27589 ( .A(n26002), .B(n27804), .Y(n22504) );
  INVX1 U27590 ( .A(reg_file[2624]), .Y(n27804) );
  NOR2X1 U27591 ( .A(n26003), .B(n27762), .Y(n22503) );
  INVX1 U27592 ( .A(reg_file[2625]), .Y(n27762) );
  NOR2X1 U27593 ( .A(n26003), .B(n27720), .Y(n22502) );
  INVX1 U27594 ( .A(reg_file[2626]), .Y(n27720) );
  NOR2X1 U27595 ( .A(n26003), .B(n27678), .Y(n22501) );
  INVX1 U27596 ( .A(reg_file[2627]), .Y(n27678) );
  NOR2X1 U27597 ( .A(n26003), .B(n27636), .Y(n22500) );
  INVX1 U27598 ( .A(reg_file[2628]), .Y(n27636) );
  NOR2X1 U27599 ( .A(n26003), .B(n27594), .Y(n22499) );
  INVX1 U27600 ( .A(reg_file[2629]), .Y(n27594) );
  NOR2X1 U27601 ( .A(n26003), .B(n27510), .Y(n22498) );
  INVX1 U27602 ( .A(reg_file[2630]), .Y(n27510) );
  NOR2X1 U27603 ( .A(n26003), .B(n27468), .Y(n22497) );
  INVX1 U27604 ( .A(reg_file[2631]), .Y(n27468) );
  NOR2X1 U27605 ( .A(n26003), .B(n27426), .Y(n22496) );
  INVX1 U27606 ( .A(reg_file[2632]), .Y(n27426) );
  NOR2X1 U27607 ( .A(n26003), .B(n27384), .Y(n22495) );
  INVX1 U27608 ( .A(reg_file[2633]), .Y(n27384) );
  NOR2X1 U27609 ( .A(n26003), .B(n27342), .Y(n22494) );
  INVX1 U27610 ( .A(reg_file[2634]), .Y(n27342) );
  NOR2X1 U27611 ( .A(n26003), .B(n27300), .Y(n22493) );
  INVX1 U27612 ( .A(reg_file[2635]), .Y(n27300) );
  NOR2X1 U27613 ( .A(n26003), .B(n27258), .Y(n22492) );
  INVX1 U27614 ( .A(reg_file[2636]), .Y(n27258) );
  NOR2X1 U27615 ( .A(n26003), .B(n27216), .Y(n22491) );
  INVX1 U27616 ( .A(reg_file[2637]), .Y(n27216) );
  NOR2X1 U27617 ( .A(n26003), .B(n27174), .Y(n22490) );
  INVX1 U27618 ( .A(reg_file[2638]), .Y(n27174) );
  NOR2X1 U27619 ( .A(n26003), .B(n27132), .Y(n22489) );
  INVX1 U27620 ( .A(reg_file[2639]), .Y(n27132) );
  NOR2X1 U27621 ( .A(n26003), .B(n27048), .Y(n22488) );
  INVX1 U27622 ( .A(reg_file[2640]), .Y(n27048) );
  NOR2X1 U27623 ( .A(n26003), .B(n27006), .Y(n22487) );
  INVX1 U27624 ( .A(reg_file[2641]), .Y(n27006) );
  NOR2X1 U27625 ( .A(n26004), .B(n26964), .Y(n22486) );
  INVX1 U27626 ( .A(reg_file[2642]), .Y(n26964) );
  NOR2X1 U27627 ( .A(n26004), .B(n26922), .Y(n22485) );
  INVX1 U27628 ( .A(reg_file[2643]), .Y(n26922) );
  NOR2X1 U27629 ( .A(n26004), .B(n26880), .Y(n22484) );
  INVX1 U27630 ( .A(reg_file[2644]), .Y(n26880) );
  NOR2X1 U27631 ( .A(n26004), .B(n26838), .Y(n22483) );
  INVX1 U27632 ( .A(reg_file[2645]), .Y(n26838) );
  NOR2X1 U27633 ( .A(n26004), .B(n26796), .Y(n22482) );
  INVX1 U27634 ( .A(reg_file[2646]), .Y(n26796) );
  NOR2X1 U27635 ( .A(n26004), .B(n26754), .Y(n22481) );
  INVX1 U27636 ( .A(reg_file[2647]), .Y(n26754) );
  NOR2X1 U27637 ( .A(n26004), .B(n26712), .Y(n22480) );
  INVX1 U27638 ( .A(reg_file[2648]), .Y(n26712) );
  NOR2X1 U27639 ( .A(n26004), .B(n26670), .Y(n22479) );
  INVX1 U27640 ( .A(reg_file[2649]), .Y(n26670) );
  NOR2X1 U27641 ( .A(n26004), .B(n26586), .Y(n22478) );
  INVX1 U27642 ( .A(reg_file[2650]), .Y(n26586) );
  NOR2X1 U27643 ( .A(n26004), .B(n26544), .Y(n22477) );
  INVX1 U27644 ( .A(reg_file[2651]), .Y(n26544) );
  NOR2X1 U27645 ( .A(n26004), .B(n26502), .Y(n22476) );
  INVX1 U27646 ( .A(reg_file[2652]), .Y(n26502) );
  NOR2X1 U27647 ( .A(n26004), .B(n26460), .Y(n22475) );
  INVX1 U27648 ( .A(reg_file[2653]), .Y(n26460) );
  NOR2X1 U27649 ( .A(n26004), .B(n26418), .Y(n22474) );
  INVX1 U27650 ( .A(reg_file[2654]), .Y(n26418) );
  NOR2X1 U27651 ( .A(n26004), .B(n26376), .Y(n22473) );
  INVX1 U27652 ( .A(reg_file[2655]), .Y(n26376) );
  NOR2X1 U27653 ( .A(n26004), .B(n26334), .Y(n22472) );
  INVX1 U27654 ( .A(reg_file[2656]), .Y(n26334) );
  NOR2X1 U27655 ( .A(n26004), .B(n26292), .Y(n22471) );
  INVX1 U27656 ( .A(reg_file[2657]), .Y(n26292) );
  NOR2X1 U27657 ( .A(n26004), .B(n26250), .Y(n22470) );
  INVX1 U27658 ( .A(reg_file[2658]), .Y(n26250) );
  NOR2X1 U27659 ( .A(n26005), .B(n26208), .Y(n22469) );
  INVX1 U27660 ( .A(reg_file[2659]), .Y(n26208) );
  NOR2X1 U27661 ( .A(n26005), .B(n31458), .Y(n22468) );
  INVX1 U27662 ( .A(reg_file[2660]), .Y(n31458) );
  NOR2X1 U27663 ( .A(n26005), .B(n31416), .Y(n22467) );
  INVX1 U27664 ( .A(reg_file[2661]), .Y(n31416) );
  NOR2X1 U27665 ( .A(n26005), .B(n31374), .Y(n22466) );
  INVX1 U27666 ( .A(reg_file[2662]), .Y(n31374) );
  NOR2X1 U27667 ( .A(n26005), .B(n31332), .Y(n22465) );
  INVX1 U27668 ( .A(reg_file[2663]), .Y(n31332) );
  NOR2X1 U27669 ( .A(n26005), .B(n31290), .Y(n22464) );
  INVX1 U27670 ( .A(reg_file[2664]), .Y(n31290) );
  NOR2X1 U27671 ( .A(n26005), .B(n31248), .Y(n22463) );
  INVX1 U27672 ( .A(reg_file[2665]), .Y(n31248) );
  NOR2X1 U27673 ( .A(n26005), .B(n31206), .Y(n22462) );
  INVX1 U27674 ( .A(reg_file[2666]), .Y(n31206) );
  NOR2X1 U27675 ( .A(n26005), .B(n31164), .Y(n22461) );
  INVX1 U27676 ( .A(reg_file[2667]), .Y(n31164) );
  NOR2X1 U27677 ( .A(n26005), .B(n31122), .Y(n22460) );
  INVX1 U27678 ( .A(reg_file[2668]), .Y(n31122) );
  NOR2X1 U27679 ( .A(n26005), .B(n31080), .Y(n22459) );
  INVX1 U27680 ( .A(reg_file[2669]), .Y(n31080) );
  NOR2X1 U27681 ( .A(n26005), .B(n30996), .Y(n22458) );
  INVX1 U27682 ( .A(reg_file[2670]), .Y(n30996) );
  NOR2X1 U27683 ( .A(n26005), .B(n30954), .Y(n22457) );
  INVX1 U27684 ( .A(reg_file[2671]), .Y(n30954) );
  NOR2X1 U27685 ( .A(n26005), .B(n30912), .Y(n22456) );
  INVX1 U27686 ( .A(reg_file[2672]), .Y(n30912) );
  NOR2X1 U27687 ( .A(n26005), .B(n30870), .Y(n22455) );
  INVX1 U27688 ( .A(reg_file[2673]), .Y(n30870) );
  NOR2X1 U27689 ( .A(n26005), .B(n30828), .Y(n22454) );
  INVX1 U27690 ( .A(reg_file[2674]), .Y(n30828) );
  NOR2X1 U27691 ( .A(n26005), .B(n30786), .Y(n22453) );
  INVX1 U27692 ( .A(reg_file[2675]), .Y(n30786) );
  NOR2X1 U27693 ( .A(n26006), .B(n30744), .Y(n22452) );
  INVX1 U27694 ( .A(reg_file[2676]), .Y(n30744) );
  NOR2X1 U27695 ( .A(n26006), .B(n30702), .Y(n22451) );
  INVX1 U27696 ( .A(reg_file[2677]), .Y(n30702) );
  NOR2X1 U27697 ( .A(n26006), .B(n30660), .Y(n22450) );
  INVX1 U27698 ( .A(reg_file[2678]), .Y(n30660) );
  NOR2X1 U27699 ( .A(n26006), .B(n30618), .Y(n22449) );
  INVX1 U27700 ( .A(reg_file[2679]), .Y(n30618) );
  NOR2X1 U27701 ( .A(n26006), .B(n30534), .Y(n22448) );
  INVX1 U27702 ( .A(reg_file[2680]), .Y(n30534) );
  NOR2X1 U27703 ( .A(n26006), .B(n30492), .Y(n22447) );
  INVX1 U27704 ( .A(reg_file[2681]), .Y(n30492) );
  NOR2X1 U27705 ( .A(n26006), .B(n30450), .Y(n22446) );
  INVX1 U27706 ( .A(reg_file[2682]), .Y(n30450) );
  NOR2X1 U27707 ( .A(n26006), .B(n30408), .Y(n22445) );
  INVX1 U27708 ( .A(reg_file[2683]), .Y(n30408) );
  NOR2X1 U27709 ( .A(n26006), .B(n30366), .Y(n22444) );
  INVX1 U27710 ( .A(reg_file[2684]), .Y(n30366) );
  NOR2X1 U27711 ( .A(n26006), .B(n30324), .Y(n22443) );
  INVX1 U27712 ( .A(reg_file[2685]), .Y(n30324) );
  NOR2X1 U27713 ( .A(n26006), .B(n30282), .Y(n22442) );
  INVX1 U27714 ( .A(reg_file[2686]), .Y(n30282) );
  NOR2X1 U27715 ( .A(n26006), .B(n30240), .Y(n22441) );
  INVX1 U27716 ( .A(reg_file[2687]), .Y(n30240) );
  NOR2X1 U27717 ( .A(n36101), .B(n35058), .Y(n36490) );
  MUX2X1 U27718 ( .B(n31520), .A(n25129), .S(n26007), .Y(n22440) );
  INVX1 U27719 ( .A(reg_file[2688]), .Y(n31520) );
  MUX2X1 U27720 ( .B(n29863), .A(n25130), .S(n26007), .Y(n22439) );
  INVX1 U27721 ( .A(reg_file[2689]), .Y(n29863) );
  MUX2X1 U27722 ( .B(n29401), .A(n25131), .S(n26007), .Y(n22438) );
  INVX1 U27723 ( .A(reg_file[2690]), .Y(n29401) );
  MUX2X1 U27724 ( .B(n28939), .A(n25132), .S(n26007), .Y(n22437) );
  INVX1 U27725 ( .A(reg_file[2691]), .Y(n28939) );
  MUX2X1 U27726 ( .B(n28477), .A(n25133), .S(n26007), .Y(n22436) );
  INVX1 U27727 ( .A(reg_file[2692]), .Y(n28477) );
  MUX2X1 U27728 ( .B(n28015), .A(n25134), .S(n26007), .Y(n22435) );
  INVX1 U27729 ( .A(reg_file[2693]), .Y(n28015) );
  MUX2X1 U27730 ( .B(n27553), .A(n25135), .S(n26007), .Y(n22434) );
  INVX1 U27731 ( .A(reg_file[2694]), .Y(n27553) );
  MUX2X1 U27732 ( .B(n27091), .A(n25136), .S(n26007), .Y(n22433) );
  INVX1 U27733 ( .A(reg_file[2695]), .Y(n27091) );
  NOR2X1 U27734 ( .A(n26007), .B(n26629), .Y(n22432) );
  INVX1 U27735 ( .A(reg_file[2696]), .Y(n26629) );
  NOR2X1 U27736 ( .A(n26007), .B(n26161), .Y(n22431) );
  INVX1 U27737 ( .A(reg_file[2697]), .Y(n26161) );
  NOR2X1 U27738 ( .A(n26007), .B(n31039), .Y(n22430) );
  INVX1 U27739 ( .A(reg_file[2698]), .Y(n31039) );
  NOR2X1 U27740 ( .A(n26007), .B(n30577), .Y(n22429) );
  INVX1 U27741 ( .A(reg_file[2699]), .Y(n30577) );
  NOR2X1 U27742 ( .A(n26007), .B(n30199), .Y(n22428) );
  INVX1 U27743 ( .A(reg_file[2700]), .Y(n30199) );
  NOR2X1 U27744 ( .A(n26007), .B(n30157), .Y(n22427) );
  INVX1 U27745 ( .A(reg_file[2701]), .Y(n30157) );
  NOR2X1 U27746 ( .A(n26008), .B(n30115), .Y(n22426) );
  INVX1 U27747 ( .A(reg_file[2702]), .Y(n30115) );
  NOR2X1 U27748 ( .A(n26008), .B(n30073), .Y(n22425) );
  INVX1 U27749 ( .A(reg_file[2703]), .Y(n30073) );
  NOR2X1 U27750 ( .A(n26008), .B(n30031), .Y(n22424) );
  INVX1 U27751 ( .A(reg_file[2704]), .Y(n30031) );
  NOR2X1 U27752 ( .A(n26008), .B(n29989), .Y(n22423) );
  INVX1 U27753 ( .A(reg_file[2705]), .Y(n29989) );
  NOR2X1 U27754 ( .A(n26008), .B(n29947), .Y(n22422) );
  INVX1 U27755 ( .A(reg_file[2706]), .Y(n29947) );
  NOR2X1 U27756 ( .A(n26008), .B(n29905), .Y(n22421) );
  INVX1 U27757 ( .A(reg_file[2707]), .Y(n29905) );
  NOR2X1 U27758 ( .A(n26008), .B(n29821), .Y(n22420) );
  INVX1 U27759 ( .A(reg_file[2708]), .Y(n29821) );
  NOR2X1 U27760 ( .A(n26008), .B(n29779), .Y(n22419) );
  INVX1 U27761 ( .A(reg_file[2709]), .Y(n29779) );
  NOR2X1 U27762 ( .A(n26008), .B(n29737), .Y(n22418) );
  INVX1 U27763 ( .A(reg_file[2710]), .Y(n29737) );
  NOR2X1 U27764 ( .A(n26008), .B(n29695), .Y(n22417) );
  INVX1 U27765 ( .A(reg_file[2711]), .Y(n29695) );
  NOR2X1 U27766 ( .A(n26008), .B(n29653), .Y(n22416) );
  INVX1 U27767 ( .A(reg_file[2712]), .Y(n29653) );
  NOR2X1 U27768 ( .A(n26008), .B(n29611), .Y(n22415) );
  INVX1 U27769 ( .A(reg_file[2713]), .Y(n29611) );
  NOR2X1 U27770 ( .A(n26008), .B(n29569), .Y(n22414) );
  INVX1 U27771 ( .A(reg_file[2714]), .Y(n29569) );
  NOR2X1 U27772 ( .A(n26008), .B(n29527), .Y(n22413) );
  INVX1 U27773 ( .A(reg_file[2715]), .Y(n29527) );
  NOR2X1 U27774 ( .A(n26008), .B(n29485), .Y(n22412) );
  INVX1 U27775 ( .A(reg_file[2716]), .Y(n29485) );
  NOR2X1 U27776 ( .A(n26008), .B(n29443), .Y(n22411) );
  INVX1 U27777 ( .A(reg_file[2717]), .Y(n29443) );
  NOR2X1 U27778 ( .A(n26008), .B(n29359), .Y(n22410) );
  INVX1 U27779 ( .A(reg_file[2718]), .Y(n29359) );
  NOR2X1 U27780 ( .A(n26009), .B(n29317), .Y(n22409) );
  INVX1 U27781 ( .A(reg_file[2719]), .Y(n29317) );
  NOR2X1 U27782 ( .A(n26009), .B(n29275), .Y(n22408) );
  INVX1 U27783 ( .A(reg_file[2720]), .Y(n29275) );
  NOR2X1 U27784 ( .A(n26009), .B(n29233), .Y(n22407) );
  INVX1 U27785 ( .A(reg_file[2721]), .Y(n29233) );
  NOR2X1 U27786 ( .A(n26009), .B(n29191), .Y(n22406) );
  INVX1 U27787 ( .A(reg_file[2722]), .Y(n29191) );
  NOR2X1 U27788 ( .A(n26009), .B(n29149), .Y(n22405) );
  INVX1 U27789 ( .A(reg_file[2723]), .Y(n29149) );
  NOR2X1 U27790 ( .A(n26009), .B(n29107), .Y(n22404) );
  INVX1 U27791 ( .A(reg_file[2724]), .Y(n29107) );
  NOR2X1 U27792 ( .A(n26009), .B(n29065), .Y(n22403) );
  INVX1 U27793 ( .A(reg_file[2725]), .Y(n29065) );
  NOR2X1 U27794 ( .A(n26009), .B(n29023), .Y(n22402) );
  INVX1 U27795 ( .A(reg_file[2726]), .Y(n29023) );
  NOR2X1 U27796 ( .A(n26009), .B(n28981), .Y(n22401) );
  INVX1 U27797 ( .A(reg_file[2727]), .Y(n28981) );
  NOR2X1 U27798 ( .A(n26009), .B(n28897), .Y(n22400) );
  INVX1 U27799 ( .A(reg_file[2728]), .Y(n28897) );
  NOR2X1 U27800 ( .A(n26009), .B(n28855), .Y(n22399) );
  INVX1 U27801 ( .A(reg_file[2729]), .Y(n28855) );
  NOR2X1 U27802 ( .A(n26009), .B(n28813), .Y(n22398) );
  INVX1 U27803 ( .A(reg_file[2730]), .Y(n28813) );
  NOR2X1 U27804 ( .A(n26009), .B(n28771), .Y(n22397) );
  INVX1 U27805 ( .A(reg_file[2731]), .Y(n28771) );
  NOR2X1 U27806 ( .A(n26009), .B(n28729), .Y(n22396) );
  INVX1 U27807 ( .A(reg_file[2732]), .Y(n28729) );
  NOR2X1 U27808 ( .A(n26009), .B(n28687), .Y(n22395) );
  INVX1 U27809 ( .A(reg_file[2733]), .Y(n28687) );
  NOR2X1 U27810 ( .A(n26009), .B(n28645), .Y(n22394) );
  INVX1 U27811 ( .A(reg_file[2734]), .Y(n28645) );
  NOR2X1 U27812 ( .A(n26009), .B(n28603), .Y(n22393) );
  INVX1 U27813 ( .A(reg_file[2735]), .Y(n28603) );
  NOR2X1 U27814 ( .A(n26010), .B(n28561), .Y(n22392) );
  INVX1 U27815 ( .A(reg_file[2736]), .Y(n28561) );
  NOR2X1 U27816 ( .A(n26010), .B(n28519), .Y(n22391) );
  INVX1 U27817 ( .A(reg_file[2737]), .Y(n28519) );
  NOR2X1 U27818 ( .A(n26010), .B(n28435), .Y(n22390) );
  INVX1 U27819 ( .A(reg_file[2738]), .Y(n28435) );
  NOR2X1 U27820 ( .A(n26010), .B(n28393), .Y(n22389) );
  INVX1 U27821 ( .A(reg_file[2739]), .Y(n28393) );
  NOR2X1 U27822 ( .A(n26010), .B(n28351), .Y(n22388) );
  INVX1 U27823 ( .A(reg_file[2740]), .Y(n28351) );
  NOR2X1 U27824 ( .A(n26010), .B(n28309), .Y(n22387) );
  INVX1 U27825 ( .A(reg_file[2741]), .Y(n28309) );
  NOR2X1 U27826 ( .A(n26010), .B(n28267), .Y(n22386) );
  INVX1 U27827 ( .A(reg_file[2742]), .Y(n28267) );
  NOR2X1 U27828 ( .A(n26010), .B(n28225), .Y(n22385) );
  INVX1 U27829 ( .A(reg_file[2743]), .Y(n28225) );
  NOR2X1 U27830 ( .A(n26010), .B(n28183), .Y(n22384) );
  INVX1 U27831 ( .A(reg_file[2744]), .Y(n28183) );
  NOR2X1 U27832 ( .A(n26010), .B(n28141), .Y(n22383) );
  INVX1 U27833 ( .A(reg_file[2745]), .Y(n28141) );
  NOR2X1 U27834 ( .A(n26010), .B(n28099), .Y(n22382) );
  INVX1 U27835 ( .A(reg_file[2746]), .Y(n28099) );
  NOR2X1 U27836 ( .A(n26010), .B(n28057), .Y(n22381) );
  INVX1 U27837 ( .A(reg_file[2747]), .Y(n28057) );
  NOR2X1 U27838 ( .A(n26010), .B(n27973), .Y(n22380) );
  INVX1 U27839 ( .A(reg_file[2748]), .Y(n27973) );
  NOR2X1 U27840 ( .A(n26010), .B(n27931), .Y(n22379) );
  INVX1 U27841 ( .A(reg_file[2749]), .Y(n27931) );
  NOR2X1 U27842 ( .A(n26010), .B(n27889), .Y(n22378) );
  INVX1 U27843 ( .A(reg_file[2750]), .Y(n27889) );
  NOR2X1 U27844 ( .A(n26010), .B(n27847), .Y(n22377) );
  INVX1 U27845 ( .A(reg_file[2751]), .Y(n27847) );
  NOR2X1 U27846 ( .A(n26010), .B(n27805), .Y(n22376) );
  INVX1 U27847 ( .A(reg_file[2752]), .Y(n27805) );
  NOR2X1 U27848 ( .A(n26011), .B(n27763), .Y(n22375) );
  INVX1 U27849 ( .A(reg_file[2753]), .Y(n27763) );
  NOR2X1 U27850 ( .A(n26011), .B(n27721), .Y(n22374) );
  INVX1 U27851 ( .A(reg_file[2754]), .Y(n27721) );
  NOR2X1 U27852 ( .A(n26011), .B(n27679), .Y(n22373) );
  INVX1 U27853 ( .A(reg_file[2755]), .Y(n27679) );
  NOR2X1 U27854 ( .A(n26011), .B(n27637), .Y(n22372) );
  INVX1 U27855 ( .A(reg_file[2756]), .Y(n27637) );
  NOR2X1 U27856 ( .A(n26011), .B(n27595), .Y(n22371) );
  INVX1 U27857 ( .A(reg_file[2757]), .Y(n27595) );
  NOR2X1 U27858 ( .A(n26011), .B(n27511), .Y(n22370) );
  INVX1 U27859 ( .A(reg_file[2758]), .Y(n27511) );
  NOR2X1 U27860 ( .A(n26011), .B(n27469), .Y(n22369) );
  INVX1 U27861 ( .A(reg_file[2759]), .Y(n27469) );
  NOR2X1 U27862 ( .A(n26011), .B(n27427), .Y(n22368) );
  INVX1 U27863 ( .A(reg_file[2760]), .Y(n27427) );
  NOR2X1 U27864 ( .A(n26011), .B(n27385), .Y(n22367) );
  INVX1 U27865 ( .A(reg_file[2761]), .Y(n27385) );
  NOR2X1 U27866 ( .A(n26011), .B(n27343), .Y(n22366) );
  INVX1 U27867 ( .A(reg_file[2762]), .Y(n27343) );
  NOR2X1 U27868 ( .A(n26011), .B(n27301), .Y(n22365) );
  INVX1 U27869 ( .A(reg_file[2763]), .Y(n27301) );
  NOR2X1 U27870 ( .A(n26011), .B(n27259), .Y(n22364) );
  INVX1 U27871 ( .A(reg_file[2764]), .Y(n27259) );
  NOR2X1 U27872 ( .A(n26011), .B(n27217), .Y(n22363) );
  INVX1 U27873 ( .A(reg_file[2765]), .Y(n27217) );
  NOR2X1 U27874 ( .A(n26011), .B(n27175), .Y(n22362) );
  INVX1 U27875 ( .A(reg_file[2766]), .Y(n27175) );
  NOR2X1 U27876 ( .A(n26011), .B(n27133), .Y(n22361) );
  INVX1 U27877 ( .A(reg_file[2767]), .Y(n27133) );
  NOR2X1 U27878 ( .A(n26011), .B(n27049), .Y(n22360) );
  INVX1 U27879 ( .A(reg_file[2768]), .Y(n27049) );
  NOR2X1 U27880 ( .A(n26011), .B(n27007), .Y(n22359) );
  INVX1 U27881 ( .A(reg_file[2769]), .Y(n27007) );
  NOR2X1 U27882 ( .A(n26012), .B(n26965), .Y(n22358) );
  INVX1 U27883 ( .A(reg_file[2770]), .Y(n26965) );
  NOR2X1 U27884 ( .A(n26012), .B(n26923), .Y(n22357) );
  INVX1 U27885 ( .A(reg_file[2771]), .Y(n26923) );
  NOR2X1 U27886 ( .A(n26012), .B(n26881), .Y(n22356) );
  INVX1 U27887 ( .A(reg_file[2772]), .Y(n26881) );
  NOR2X1 U27888 ( .A(n26012), .B(n26839), .Y(n22355) );
  INVX1 U27889 ( .A(reg_file[2773]), .Y(n26839) );
  NOR2X1 U27890 ( .A(n26012), .B(n26797), .Y(n22354) );
  INVX1 U27891 ( .A(reg_file[2774]), .Y(n26797) );
  NOR2X1 U27892 ( .A(n26012), .B(n26755), .Y(n22353) );
  INVX1 U27893 ( .A(reg_file[2775]), .Y(n26755) );
  NOR2X1 U27894 ( .A(n26012), .B(n26713), .Y(n22352) );
  INVX1 U27895 ( .A(reg_file[2776]), .Y(n26713) );
  NOR2X1 U27896 ( .A(n26012), .B(n26671), .Y(n22351) );
  INVX1 U27897 ( .A(reg_file[2777]), .Y(n26671) );
  NOR2X1 U27898 ( .A(n26012), .B(n26587), .Y(n22350) );
  INVX1 U27899 ( .A(reg_file[2778]), .Y(n26587) );
  NOR2X1 U27900 ( .A(n26012), .B(n26545), .Y(n22349) );
  INVX1 U27901 ( .A(reg_file[2779]), .Y(n26545) );
  NOR2X1 U27902 ( .A(n26012), .B(n26503), .Y(n22348) );
  INVX1 U27903 ( .A(reg_file[2780]), .Y(n26503) );
  NOR2X1 U27904 ( .A(n26012), .B(n26461), .Y(n22347) );
  INVX1 U27905 ( .A(reg_file[2781]), .Y(n26461) );
  NOR2X1 U27906 ( .A(n26012), .B(n26419), .Y(n22346) );
  INVX1 U27907 ( .A(reg_file[2782]), .Y(n26419) );
  NOR2X1 U27908 ( .A(n26012), .B(n26377), .Y(n22345) );
  INVX1 U27909 ( .A(reg_file[2783]), .Y(n26377) );
  NOR2X1 U27910 ( .A(n26012), .B(n26335), .Y(n22344) );
  INVX1 U27911 ( .A(reg_file[2784]), .Y(n26335) );
  NOR2X1 U27912 ( .A(n26012), .B(n26293), .Y(n22343) );
  INVX1 U27913 ( .A(reg_file[2785]), .Y(n26293) );
  NOR2X1 U27914 ( .A(n26012), .B(n26251), .Y(n22342) );
  INVX1 U27915 ( .A(reg_file[2786]), .Y(n26251) );
  NOR2X1 U27916 ( .A(n26013), .B(n26209), .Y(n22341) );
  INVX1 U27917 ( .A(reg_file[2787]), .Y(n26209) );
  NOR2X1 U27918 ( .A(n26013), .B(n31459), .Y(n22340) );
  INVX1 U27919 ( .A(reg_file[2788]), .Y(n31459) );
  NOR2X1 U27920 ( .A(n26013), .B(n31417), .Y(n22339) );
  INVX1 U27921 ( .A(reg_file[2789]), .Y(n31417) );
  NOR2X1 U27922 ( .A(n26013), .B(n31375), .Y(n22338) );
  INVX1 U27923 ( .A(reg_file[2790]), .Y(n31375) );
  NOR2X1 U27924 ( .A(n26013), .B(n31333), .Y(n22337) );
  INVX1 U27925 ( .A(reg_file[2791]), .Y(n31333) );
  NOR2X1 U27926 ( .A(n26013), .B(n31291), .Y(n22336) );
  INVX1 U27927 ( .A(reg_file[2792]), .Y(n31291) );
  NOR2X1 U27928 ( .A(n26013), .B(n31249), .Y(n22335) );
  INVX1 U27929 ( .A(reg_file[2793]), .Y(n31249) );
  NOR2X1 U27930 ( .A(n26013), .B(n31207), .Y(n22334) );
  INVX1 U27931 ( .A(reg_file[2794]), .Y(n31207) );
  NOR2X1 U27932 ( .A(n26013), .B(n31165), .Y(n22333) );
  INVX1 U27933 ( .A(reg_file[2795]), .Y(n31165) );
  NOR2X1 U27934 ( .A(n26013), .B(n31123), .Y(n22332) );
  INVX1 U27935 ( .A(reg_file[2796]), .Y(n31123) );
  NOR2X1 U27936 ( .A(n26013), .B(n31081), .Y(n22331) );
  INVX1 U27937 ( .A(reg_file[2797]), .Y(n31081) );
  NOR2X1 U27938 ( .A(n26013), .B(n30997), .Y(n22330) );
  INVX1 U27939 ( .A(reg_file[2798]), .Y(n30997) );
  NOR2X1 U27940 ( .A(n26013), .B(n30955), .Y(n22329) );
  INVX1 U27941 ( .A(reg_file[2799]), .Y(n30955) );
  NOR2X1 U27942 ( .A(n26013), .B(n30913), .Y(n22328) );
  INVX1 U27943 ( .A(reg_file[2800]), .Y(n30913) );
  NOR2X1 U27944 ( .A(n26013), .B(n30871), .Y(n22327) );
  INVX1 U27945 ( .A(reg_file[2801]), .Y(n30871) );
  NOR2X1 U27946 ( .A(n26013), .B(n30829), .Y(n22326) );
  INVX1 U27947 ( .A(reg_file[2802]), .Y(n30829) );
  NOR2X1 U27948 ( .A(n26013), .B(n30787), .Y(n22325) );
  INVX1 U27949 ( .A(reg_file[2803]), .Y(n30787) );
  NOR2X1 U27950 ( .A(n26014), .B(n30745), .Y(n22324) );
  INVX1 U27951 ( .A(reg_file[2804]), .Y(n30745) );
  NOR2X1 U27952 ( .A(n26014), .B(n30703), .Y(n22323) );
  INVX1 U27953 ( .A(reg_file[2805]), .Y(n30703) );
  NOR2X1 U27954 ( .A(n26014), .B(n30661), .Y(n22322) );
  INVX1 U27955 ( .A(reg_file[2806]), .Y(n30661) );
  NOR2X1 U27956 ( .A(n26014), .B(n30619), .Y(n22321) );
  INVX1 U27957 ( .A(reg_file[2807]), .Y(n30619) );
  NOR2X1 U27958 ( .A(n26014), .B(n30535), .Y(n22320) );
  INVX1 U27959 ( .A(reg_file[2808]), .Y(n30535) );
  NOR2X1 U27960 ( .A(n26014), .B(n30493), .Y(n22319) );
  INVX1 U27961 ( .A(reg_file[2809]), .Y(n30493) );
  NOR2X1 U27962 ( .A(n26014), .B(n30451), .Y(n22318) );
  INVX1 U27963 ( .A(reg_file[2810]), .Y(n30451) );
  NOR2X1 U27964 ( .A(n26014), .B(n30409), .Y(n22317) );
  INVX1 U27965 ( .A(reg_file[2811]), .Y(n30409) );
  NOR2X1 U27966 ( .A(n26014), .B(n30367), .Y(n22316) );
  INVX1 U27967 ( .A(reg_file[2812]), .Y(n30367) );
  NOR2X1 U27968 ( .A(n26014), .B(n30325), .Y(n22315) );
  INVX1 U27969 ( .A(reg_file[2813]), .Y(n30325) );
  NOR2X1 U27970 ( .A(n26014), .B(n30283), .Y(n22314) );
  INVX1 U27971 ( .A(reg_file[2814]), .Y(n30283) );
  NOR2X1 U27972 ( .A(n26014), .B(n30241), .Y(n22313) );
  INVX1 U27973 ( .A(reg_file[2815]), .Y(n30241) );
  NOR2X1 U27974 ( .A(n36231), .B(n35058), .Y(n36491) );
  MUX2X1 U27975 ( .B(n31524), .A(n25129), .S(n26015), .Y(n22312) );
  INVX1 U27976 ( .A(reg_file[2816]), .Y(n31524) );
  MUX2X1 U27977 ( .B(n29864), .A(n25130), .S(n26015), .Y(n22311) );
  INVX1 U27978 ( .A(reg_file[2817]), .Y(n29864) );
  MUX2X1 U27979 ( .B(n29402), .A(n25131), .S(n26015), .Y(n22310) );
  INVX1 U27980 ( .A(reg_file[2818]), .Y(n29402) );
  MUX2X1 U27981 ( .B(n28940), .A(n25132), .S(n26015), .Y(n22309) );
  INVX1 U27982 ( .A(reg_file[2819]), .Y(n28940) );
  MUX2X1 U27983 ( .B(n28478), .A(n25133), .S(n26015), .Y(n22308) );
  INVX1 U27984 ( .A(reg_file[2820]), .Y(n28478) );
  MUX2X1 U27985 ( .B(n28016), .A(n25134), .S(n26015), .Y(n22307) );
  INVX1 U27986 ( .A(reg_file[2821]), .Y(n28016) );
  MUX2X1 U27987 ( .B(n27554), .A(n25135), .S(n26015), .Y(n22306) );
  INVX1 U27988 ( .A(reg_file[2822]), .Y(n27554) );
  MUX2X1 U27989 ( .B(n27092), .A(n25136), .S(n26015), .Y(n22305) );
  INVX1 U27990 ( .A(reg_file[2823]), .Y(n27092) );
  NOR2X1 U27991 ( .A(n26015), .B(n26630), .Y(n22304) );
  INVX1 U27992 ( .A(reg_file[2824]), .Y(n26630) );
  NOR2X1 U27993 ( .A(n26015), .B(n26163), .Y(n22303) );
  INVX1 U27994 ( .A(reg_file[2825]), .Y(n26163) );
  NOR2X1 U27995 ( .A(n26015), .B(n31040), .Y(n22302) );
  INVX1 U27996 ( .A(reg_file[2826]), .Y(n31040) );
  NOR2X1 U27997 ( .A(n26015), .B(n30578), .Y(n22301) );
  INVX1 U27998 ( .A(reg_file[2827]), .Y(n30578) );
  NOR2X1 U27999 ( .A(n26015), .B(n30200), .Y(n22300) );
  INVX1 U28000 ( .A(reg_file[2828]), .Y(n30200) );
  NOR2X1 U28001 ( .A(n26015), .B(n30158), .Y(n22299) );
  INVX1 U28002 ( .A(reg_file[2829]), .Y(n30158) );
  NOR2X1 U28003 ( .A(n26016), .B(n30116), .Y(n22298) );
  INVX1 U28004 ( .A(reg_file[2830]), .Y(n30116) );
  NOR2X1 U28005 ( .A(n26016), .B(n30074), .Y(n22297) );
  INVX1 U28006 ( .A(reg_file[2831]), .Y(n30074) );
  NOR2X1 U28007 ( .A(n26016), .B(n30032), .Y(n22296) );
  INVX1 U28008 ( .A(reg_file[2832]), .Y(n30032) );
  NOR2X1 U28009 ( .A(n26016), .B(n29990), .Y(n22295) );
  INVX1 U28010 ( .A(reg_file[2833]), .Y(n29990) );
  NOR2X1 U28011 ( .A(n26016), .B(n29948), .Y(n22294) );
  INVX1 U28012 ( .A(reg_file[2834]), .Y(n29948) );
  NOR2X1 U28013 ( .A(n26016), .B(n29906), .Y(n22293) );
  INVX1 U28014 ( .A(reg_file[2835]), .Y(n29906) );
  NOR2X1 U28015 ( .A(n26016), .B(n29822), .Y(n22292) );
  INVX1 U28016 ( .A(reg_file[2836]), .Y(n29822) );
  NOR2X1 U28017 ( .A(n26016), .B(n29780), .Y(n22291) );
  INVX1 U28018 ( .A(reg_file[2837]), .Y(n29780) );
  NOR2X1 U28019 ( .A(n26016), .B(n29738), .Y(n22290) );
  INVX1 U28020 ( .A(reg_file[2838]), .Y(n29738) );
  NOR2X1 U28021 ( .A(n26016), .B(n29696), .Y(n22289) );
  INVX1 U28022 ( .A(reg_file[2839]), .Y(n29696) );
  NOR2X1 U28023 ( .A(n26016), .B(n29654), .Y(n22288) );
  INVX1 U28024 ( .A(reg_file[2840]), .Y(n29654) );
  NOR2X1 U28025 ( .A(n26016), .B(n29612), .Y(n22287) );
  INVX1 U28026 ( .A(reg_file[2841]), .Y(n29612) );
  NOR2X1 U28027 ( .A(n26016), .B(n29570), .Y(n22286) );
  INVX1 U28028 ( .A(reg_file[2842]), .Y(n29570) );
  NOR2X1 U28029 ( .A(n26016), .B(n29528), .Y(n22285) );
  INVX1 U28030 ( .A(reg_file[2843]), .Y(n29528) );
  NOR2X1 U28031 ( .A(n26016), .B(n29486), .Y(n22284) );
  INVX1 U28032 ( .A(reg_file[2844]), .Y(n29486) );
  NOR2X1 U28033 ( .A(n26016), .B(n29444), .Y(n22283) );
  INVX1 U28034 ( .A(reg_file[2845]), .Y(n29444) );
  NOR2X1 U28035 ( .A(n26016), .B(n29360), .Y(n22282) );
  INVX1 U28036 ( .A(reg_file[2846]), .Y(n29360) );
  NOR2X1 U28037 ( .A(n26017), .B(n29318), .Y(n22281) );
  INVX1 U28038 ( .A(reg_file[2847]), .Y(n29318) );
  NOR2X1 U28039 ( .A(n26017), .B(n29276), .Y(n22280) );
  INVX1 U28040 ( .A(reg_file[2848]), .Y(n29276) );
  NOR2X1 U28041 ( .A(n26017), .B(n29234), .Y(n22279) );
  INVX1 U28042 ( .A(reg_file[2849]), .Y(n29234) );
  NOR2X1 U28043 ( .A(n26017), .B(n29192), .Y(n22278) );
  INVX1 U28044 ( .A(reg_file[2850]), .Y(n29192) );
  NOR2X1 U28045 ( .A(n26017), .B(n29150), .Y(n22277) );
  INVX1 U28046 ( .A(reg_file[2851]), .Y(n29150) );
  NOR2X1 U28047 ( .A(n26017), .B(n29108), .Y(n22276) );
  INVX1 U28048 ( .A(reg_file[2852]), .Y(n29108) );
  NOR2X1 U28049 ( .A(n26017), .B(n29066), .Y(n22275) );
  INVX1 U28050 ( .A(reg_file[2853]), .Y(n29066) );
  NOR2X1 U28051 ( .A(n26017), .B(n29024), .Y(n22274) );
  INVX1 U28052 ( .A(reg_file[2854]), .Y(n29024) );
  NOR2X1 U28053 ( .A(n26017), .B(n28982), .Y(n22273) );
  INVX1 U28054 ( .A(reg_file[2855]), .Y(n28982) );
  NOR2X1 U28055 ( .A(n26017), .B(n28898), .Y(n22272) );
  INVX1 U28056 ( .A(reg_file[2856]), .Y(n28898) );
  NOR2X1 U28057 ( .A(n26017), .B(n28856), .Y(n22271) );
  INVX1 U28058 ( .A(reg_file[2857]), .Y(n28856) );
  NOR2X1 U28059 ( .A(n26017), .B(n28814), .Y(n22270) );
  INVX1 U28060 ( .A(reg_file[2858]), .Y(n28814) );
  NOR2X1 U28061 ( .A(n26017), .B(n28772), .Y(n22269) );
  INVX1 U28062 ( .A(reg_file[2859]), .Y(n28772) );
  NOR2X1 U28063 ( .A(n26017), .B(n28730), .Y(n22268) );
  INVX1 U28064 ( .A(reg_file[2860]), .Y(n28730) );
  NOR2X1 U28065 ( .A(n26017), .B(n28688), .Y(n22267) );
  INVX1 U28066 ( .A(reg_file[2861]), .Y(n28688) );
  NOR2X1 U28067 ( .A(n26017), .B(n28646), .Y(n22266) );
  INVX1 U28068 ( .A(reg_file[2862]), .Y(n28646) );
  NOR2X1 U28069 ( .A(n26017), .B(n28604), .Y(n22265) );
  INVX1 U28070 ( .A(reg_file[2863]), .Y(n28604) );
  NOR2X1 U28071 ( .A(n26018), .B(n28562), .Y(n22264) );
  INVX1 U28072 ( .A(reg_file[2864]), .Y(n28562) );
  NOR2X1 U28073 ( .A(n26018), .B(n28520), .Y(n22263) );
  INVX1 U28074 ( .A(reg_file[2865]), .Y(n28520) );
  NOR2X1 U28075 ( .A(n26018), .B(n28436), .Y(n22262) );
  INVX1 U28076 ( .A(reg_file[2866]), .Y(n28436) );
  NOR2X1 U28077 ( .A(n26018), .B(n28394), .Y(n22261) );
  INVX1 U28078 ( .A(reg_file[2867]), .Y(n28394) );
  NOR2X1 U28079 ( .A(n26018), .B(n28352), .Y(n22260) );
  INVX1 U28080 ( .A(reg_file[2868]), .Y(n28352) );
  NOR2X1 U28081 ( .A(n26018), .B(n28310), .Y(n22259) );
  INVX1 U28082 ( .A(reg_file[2869]), .Y(n28310) );
  NOR2X1 U28083 ( .A(n26018), .B(n28268), .Y(n22258) );
  INVX1 U28084 ( .A(reg_file[2870]), .Y(n28268) );
  NOR2X1 U28085 ( .A(n26018), .B(n28226), .Y(n22257) );
  INVX1 U28086 ( .A(reg_file[2871]), .Y(n28226) );
  NOR2X1 U28087 ( .A(n26018), .B(n28184), .Y(n22256) );
  INVX1 U28088 ( .A(reg_file[2872]), .Y(n28184) );
  NOR2X1 U28089 ( .A(n26018), .B(n28142), .Y(n22255) );
  INVX1 U28090 ( .A(reg_file[2873]), .Y(n28142) );
  NOR2X1 U28091 ( .A(n26018), .B(n28100), .Y(n22254) );
  INVX1 U28092 ( .A(reg_file[2874]), .Y(n28100) );
  NOR2X1 U28093 ( .A(n26018), .B(n28058), .Y(n22253) );
  INVX1 U28094 ( .A(reg_file[2875]), .Y(n28058) );
  NOR2X1 U28095 ( .A(n26018), .B(n27974), .Y(n22252) );
  INVX1 U28096 ( .A(reg_file[2876]), .Y(n27974) );
  NOR2X1 U28097 ( .A(n26018), .B(n27932), .Y(n22251) );
  INVX1 U28098 ( .A(reg_file[2877]), .Y(n27932) );
  NOR2X1 U28099 ( .A(n26018), .B(n27890), .Y(n22250) );
  INVX1 U28100 ( .A(reg_file[2878]), .Y(n27890) );
  NOR2X1 U28101 ( .A(n26018), .B(n27848), .Y(n22249) );
  INVX1 U28102 ( .A(reg_file[2879]), .Y(n27848) );
  NOR2X1 U28103 ( .A(n26018), .B(n27806), .Y(n22248) );
  INVX1 U28104 ( .A(reg_file[2880]), .Y(n27806) );
  NOR2X1 U28105 ( .A(n26019), .B(n27764), .Y(n22247) );
  INVX1 U28106 ( .A(reg_file[2881]), .Y(n27764) );
  NOR2X1 U28107 ( .A(n26019), .B(n27722), .Y(n22246) );
  INVX1 U28108 ( .A(reg_file[2882]), .Y(n27722) );
  NOR2X1 U28109 ( .A(n26019), .B(n27680), .Y(n22245) );
  INVX1 U28110 ( .A(reg_file[2883]), .Y(n27680) );
  NOR2X1 U28111 ( .A(n26019), .B(n27638), .Y(n22244) );
  INVX1 U28112 ( .A(reg_file[2884]), .Y(n27638) );
  NOR2X1 U28113 ( .A(n26019), .B(n27596), .Y(n22243) );
  INVX1 U28114 ( .A(reg_file[2885]), .Y(n27596) );
  NOR2X1 U28115 ( .A(n26019), .B(n27512), .Y(n22242) );
  INVX1 U28116 ( .A(reg_file[2886]), .Y(n27512) );
  NOR2X1 U28117 ( .A(n26019), .B(n27470), .Y(n22241) );
  INVX1 U28118 ( .A(reg_file[2887]), .Y(n27470) );
  NOR2X1 U28119 ( .A(n26019), .B(n27428), .Y(n22240) );
  INVX1 U28120 ( .A(reg_file[2888]), .Y(n27428) );
  NOR2X1 U28121 ( .A(n26019), .B(n27386), .Y(n22239) );
  INVX1 U28122 ( .A(reg_file[2889]), .Y(n27386) );
  NOR2X1 U28123 ( .A(n26019), .B(n27344), .Y(n22238) );
  INVX1 U28124 ( .A(reg_file[2890]), .Y(n27344) );
  NOR2X1 U28125 ( .A(n26019), .B(n27302), .Y(n22237) );
  INVX1 U28126 ( .A(reg_file[2891]), .Y(n27302) );
  NOR2X1 U28127 ( .A(n26019), .B(n27260), .Y(n22236) );
  INVX1 U28128 ( .A(reg_file[2892]), .Y(n27260) );
  NOR2X1 U28129 ( .A(n26019), .B(n27218), .Y(n22235) );
  INVX1 U28130 ( .A(reg_file[2893]), .Y(n27218) );
  NOR2X1 U28131 ( .A(n26019), .B(n27176), .Y(n22234) );
  INVX1 U28132 ( .A(reg_file[2894]), .Y(n27176) );
  NOR2X1 U28133 ( .A(n26019), .B(n27134), .Y(n22233) );
  INVX1 U28134 ( .A(reg_file[2895]), .Y(n27134) );
  NOR2X1 U28135 ( .A(n26019), .B(n27050), .Y(n22232) );
  INVX1 U28136 ( .A(reg_file[2896]), .Y(n27050) );
  NOR2X1 U28137 ( .A(n26019), .B(n27008), .Y(n22231) );
  INVX1 U28138 ( .A(reg_file[2897]), .Y(n27008) );
  NOR2X1 U28139 ( .A(n26020), .B(n26966), .Y(n22230) );
  INVX1 U28140 ( .A(reg_file[2898]), .Y(n26966) );
  NOR2X1 U28141 ( .A(n26020), .B(n26924), .Y(n22229) );
  INVX1 U28142 ( .A(reg_file[2899]), .Y(n26924) );
  NOR2X1 U28143 ( .A(n26020), .B(n26882), .Y(n22228) );
  INVX1 U28144 ( .A(reg_file[2900]), .Y(n26882) );
  NOR2X1 U28145 ( .A(n26020), .B(n26840), .Y(n22227) );
  INVX1 U28146 ( .A(reg_file[2901]), .Y(n26840) );
  NOR2X1 U28147 ( .A(n26020), .B(n26798), .Y(n22226) );
  INVX1 U28148 ( .A(reg_file[2902]), .Y(n26798) );
  NOR2X1 U28149 ( .A(n26020), .B(n26756), .Y(n22225) );
  INVX1 U28150 ( .A(reg_file[2903]), .Y(n26756) );
  NOR2X1 U28151 ( .A(n26020), .B(n26714), .Y(n22224) );
  INVX1 U28152 ( .A(reg_file[2904]), .Y(n26714) );
  NOR2X1 U28153 ( .A(n26020), .B(n26672), .Y(n22223) );
  INVX1 U28154 ( .A(reg_file[2905]), .Y(n26672) );
  NOR2X1 U28155 ( .A(n26020), .B(n26588), .Y(n22222) );
  INVX1 U28156 ( .A(reg_file[2906]), .Y(n26588) );
  NOR2X1 U28157 ( .A(n26020), .B(n26546), .Y(n22221) );
  INVX1 U28158 ( .A(reg_file[2907]), .Y(n26546) );
  NOR2X1 U28159 ( .A(n26020), .B(n26504), .Y(n22220) );
  INVX1 U28160 ( .A(reg_file[2908]), .Y(n26504) );
  NOR2X1 U28161 ( .A(n26020), .B(n26462), .Y(n22219) );
  INVX1 U28162 ( .A(reg_file[2909]), .Y(n26462) );
  NOR2X1 U28163 ( .A(n26020), .B(n26420), .Y(n22218) );
  INVX1 U28164 ( .A(reg_file[2910]), .Y(n26420) );
  NOR2X1 U28165 ( .A(n26020), .B(n26378), .Y(n22217) );
  INVX1 U28166 ( .A(reg_file[2911]), .Y(n26378) );
  NOR2X1 U28167 ( .A(n26020), .B(n26336), .Y(n22216) );
  INVX1 U28168 ( .A(reg_file[2912]), .Y(n26336) );
  NOR2X1 U28169 ( .A(n26020), .B(n26294), .Y(n22215) );
  INVX1 U28170 ( .A(reg_file[2913]), .Y(n26294) );
  NOR2X1 U28171 ( .A(n26020), .B(n26252), .Y(n22214) );
  INVX1 U28172 ( .A(reg_file[2914]), .Y(n26252) );
  NOR2X1 U28173 ( .A(n26021), .B(n26210), .Y(n22213) );
  INVX1 U28174 ( .A(reg_file[2915]), .Y(n26210) );
  NOR2X1 U28175 ( .A(n26021), .B(n31460), .Y(n22212) );
  INVX1 U28176 ( .A(reg_file[2916]), .Y(n31460) );
  NOR2X1 U28177 ( .A(n26021), .B(n31418), .Y(n22211) );
  INVX1 U28178 ( .A(reg_file[2917]), .Y(n31418) );
  NOR2X1 U28179 ( .A(n26021), .B(n31376), .Y(n22210) );
  INVX1 U28180 ( .A(reg_file[2918]), .Y(n31376) );
  NOR2X1 U28181 ( .A(n26021), .B(n31334), .Y(n22209) );
  INVX1 U28182 ( .A(reg_file[2919]), .Y(n31334) );
  NOR2X1 U28183 ( .A(n26021), .B(n31292), .Y(n22208) );
  INVX1 U28184 ( .A(reg_file[2920]), .Y(n31292) );
  NOR2X1 U28185 ( .A(n26021), .B(n31250), .Y(n22207) );
  INVX1 U28186 ( .A(reg_file[2921]), .Y(n31250) );
  NOR2X1 U28187 ( .A(n26021), .B(n31208), .Y(n22206) );
  INVX1 U28188 ( .A(reg_file[2922]), .Y(n31208) );
  NOR2X1 U28189 ( .A(n26021), .B(n31166), .Y(n22205) );
  INVX1 U28190 ( .A(reg_file[2923]), .Y(n31166) );
  NOR2X1 U28191 ( .A(n26021), .B(n31124), .Y(n22204) );
  INVX1 U28192 ( .A(reg_file[2924]), .Y(n31124) );
  NOR2X1 U28193 ( .A(n26021), .B(n31082), .Y(n22203) );
  INVX1 U28194 ( .A(reg_file[2925]), .Y(n31082) );
  NOR2X1 U28195 ( .A(n26021), .B(n30998), .Y(n22202) );
  INVX1 U28196 ( .A(reg_file[2926]), .Y(n30998) );
  NOR2X1 U28197 ( .A(n26021), .B(n30956), .Y(n22201) );
  INVX1 U28198 ( .A(reg_file[2927]), .Y(n30956) );
  NOR2X1 U28199 ( .A(n26021), .B(n30914), .Y(n22200) );
  INVX1 U28200 ( .A(reg_file[2928]), .Y(n30914) );
  NOR2X1 U28201 ( .A(n26021), .B(n30872), .Y(n22199) );
  INVX1 U28202 ( .A(reg_file[2929]), .Y(n30872) );
  NOR2X1 U28203 ( .A(n26021), .B(n30830), .Y(n22198) );
  INVX1 U28204 ( .A(reg_file[2930]), .Y(n30830) );
  NOR2X1 U28205 ( .A(n26021), .B(n30788), .Y(n22197) );
  INVX1 U28206 ( .A(reg_file[2931]), .Y(n30788) );
  NOR2X1 U28207 ( .A(n26022), .B(n30746), .Y(n22196) );
  INVX1 U28208 ( .A(reg_file[2932]), .Y(n30746) );
  NOR2X1 U28209 ( .A(n26022), .B(n30704), .Y(n22195) );
  INVX1 U28210 ( .A(reg_file[2933]), .Y(n30704) );
  NOR2X1 U28211 ( .A(n26022), .B(n30662), .Y(n22194) );
  INVX1 U28212 ( .A(reg_file[2934]), .Y(n30662) );
  NOR2X1 U28213 ( .A(n26022), .B(n30620), .Y(n22193) );
  INVX1 U28214 ( .A(reg_file[2935]), .Y(n30620) );
  NOR2X1 U28215 ( .A(n26022), .B(n30536), .Y(n22192) );
  INVX1 U28216 ( .A(reg_file[2936]), .Y(n30536) );
  NOR2X1 U28217 ( .A(n26022), .B(n30494), .Y(n22191) );
  INVX1 U28218 ( .A(reg_file[2937]), .Y(n30494) );
  NOR2X1 U28219 ( .A(n26022), .B(n30452), .Y(n22190) );
  INVX1 U28220 ( .A(reg_file[2938]), .Y(n30452) );
  NOR2X1 U28221 ( .A(n26022), .B(n30410), .Y(n22189) );
  INVX1 U28222 ( .A(reg_file[2939]), .Y(n30410) );
  NOR2X1 U28223 ( .A(n26022), .B(n30368), .Y(n22188) );
  INVX1 U28224 ( .A(reg_file[2940]), .Y(n30368) );
  NOR2X1 U28225 ( .A(n26022), .B(n30326), .Y(n22187) );
  INVX1 U28226 ( .A(reg_file[2941]), .Y(n30326) );
  NOR2X1 U28227 ( .A(n26022), .B(n30284), .Y(n22186) );
  INVX1 U28228 ( .A(reg_file[2942]), .Y(n30284) );
  NOR2X1 U28229 ( .A(n26022), .B(n30242), .Y(n22185) );
  INVX1 U28230 ( .A(reg_file[2943]), .Y(n30242) );
  NOR2X1 U28231 ( .A(n36101), .B(n35317), .Y(n36492) );
  NAND3X1 U28232 ( .A(n35320), .B(n35318), .C(wraddr[4]), .Y(n36101) );
  MUX2X1 U28233 ( .B(n31525), .A(n25129), .S(n26023), .Y(n22184) );
  INVX1 U28234 ( .A(reg_file[2944]), .Y(n31525) );
  MUX2X1 U28235 ( .B(n29865), .A(n25130), .S(n26023), .Y(n22183) );
  INVX1 U28236 ( .A(reg_file[2945]), .Y(n29865) );
  MUX2X1 U28237 ( .B(n29403), .A(n25131), .S(n26023), .Y(n22182) );
  INVX1 U28238 ( .A(reg_file[2946]), .Y(n29403) );
  MUX2X1 U28239 ( .B(n28941), .A(n25132), .S(n26023), .Y(n22181) );
  INVX1 U28240 ( .A(reg_file[2947]), .Y(n28941) );
  MUX2X1 U28241 ( .B(n28479), .A(n25133), .S(n26023), .Y(n22180) );
  INVX1 U28242 ( .A(reg_file[2948]), .Y(n28479) );
  MUX2X1 U28243 ( .B(n28017), .A(n25134), .S(n26023), .Y(n22179) );
  INVX1 U28244 ( .A(reg_file[2949]), .Y(n28017) );
  MUX2X1 U28245 ( .B(n27555), .A(n25135), .S(n26023), .Y(n22178) );
  INVX1 U28246 ( .A(reg_file[2950]), .Y(n27555) );
  MUX2X1 U28247 ( .B(n27093), .A(n25136), .S(n26023), .Y(n22177) );
  INVX1 U28248 ( .A(reg_file[2951]), .Y(n27093) );
  NOR2X1 U28249 ( .A(n26023), .B(n26631), .Y(n22176) );
  INVX1 U28250 ( .A(reg_file[2952]), .Y(n26631) );
  NOR2X1 U28251 ( .A(n26023), .B(n26165), .Y(n22175) );
  INVX1 U28252 ( .A(reg_file[2953]), .Y(n26165) );
  NOR2X1 U28253 ( .A(n26023), .B(n31041), .Y(n22174) );
  INVX1 U28254 ( .A(reg_file[2954]), .Y(n31041) );
  NOR2X1 U28255 ( .A(n26023), .B(n30579), .Y(n22173) );
  INVX1 U28256 ( .A(reg_file[2955]), .Y(n30579) );
  NOR2X1 U28257 ( .A(n26023), .B(n30201), .Y(n22172) );
  INVX1 U28258 ( .A(reg_file[2956]), .Y(n30201) );
  NOR2X1 U28259 ( .A(n26023), .B(n30159), .Y(n22171) );
  INVX1 U28260 ( .A(reg_file[2957]), .Y(n30159) );
  NOR2X1 U28261 ( .A(n26024), .B(n30117), .Y(n22170) );
  INVX1 U28262 ( .A(reg_file[2958]), .Y(n30117) );
  NOR2X1 U28263 ( .A(n26024), .B(n30075), .Y(n22169) );
  INVX1 U28264 ( .A(reg_file[2959]), .Y(n30075) );
  NOR2X1 U28265 ( .A(n26024), .B(n30033), .Y(n22168) );
  INVX1 U28266 ( .A(reg_file[2960]), .Y(n30033) );
  NOR2X1 U28267 ( .A(n26024), .B(n29991), .Y(n22167) );
  INVX1 U28268 ( .A(reg_file[2961]), .Y(n29991) );
  NOR2X1 U28269 ( .A(n26024), .B(n29949), .Y(n22166) );
  INVX1 U28270 ( .A(reg_file[2962]), .Y(n29949) );
  NOR2X1 U28271 ( .A(n26024), .B(n29907), .Y(n22165) );
  INVX1 U28272 ( .A(reg_file[2963]), .Y(n29907) );
  NOR2X1 U28273 ( .A(n26024), .B(n29823), .Y(n22164) );
  INVX1 U28274 ( .A(reg_file[2964]), .Y(n29823) );
  NOR2X1 U28275 ( .A(n26024), .B(n29781), .Y(n22163) );
  INVX1 U28276 ( .A(reg_file[2965]), .Y(n29781) );
  NOR2X1 U28277 ( .A(n26024), .B(n29739), .Y(n22162) );
  INVX1 U28278 ( .A(reg_file[2966]), .Y(n29739) );
  NOR2X1 U28279 ( .A(n26024), .B(n29697), .Y(n22161) );
  INVX1 U28280 ( .A(reg_file[2967]), .Y(n29697) );
  NOR2X1 U28281 ( .A(n26024), .B(n29655), .Y(n22160) );
  INVX1 U28282 ( .A(reg_file[2968]), .Y(n29655) );
  NOR2X1 U28283 ( .A(n26024), .B(n29613), .Y(n22159) );
  INVX1 U28284 ( .A(reg_file[2969]), .Y(n29613) );
  NOR2X1 U28285 ( .A(n26024), .B(n29571), .Y(n22158) );
  INVX1 U28286 ( .A(reg_file[2970]), .Y(n29571) );
  NOR2X1 U28287 ( .A(n26024), .B(n29529), .Y(n22157) );
  INVX1 U28288 ( .A(reg_file[2971]), .Y(n29529) );
  NOR2X1 U28289 ( .A(n26024), .B(n29487), .Y(n22156) );
  INVX1 U28290 ( .A(reg_file[2972]), .Y(n29487) );
  NOR2X1 U28291 ( .A(n26024), .B(n29445), .Y(n22155) );
  INVX1 U28292 ( .A(reg_file[2973]), .Y(n29445) );
  NOR2X1 U28293 ( .A(n26024), .B(n29361), .Y(n22154) );
  INVX1 U28294 ( .A(reg_file[2974]), .Y(n29361) );
  NOR2X1 U28295 ( .A(n26025), .B(n29319), .Y(n22153) );
  INVX1 U28296 ( .A(reg_file[2975]), .Y(n29319) );
  NOR2X1 U28297 ( .A(n26025), .B(n29277), .Y(n22152) );
  INVX1 U28298 ( .A(reg_file[2976]), .Y(n29277) );
  NOR2X1 U28299 ( .A(n26025), .B(n29235), .Y(n22151) );
  INVX1 U28300 ( .A(reg_file[2977]), .Y(n29235) );
  NOR2X1 U28301 ( .A(n26025), .B(n29193), .Y(n22150) );
  INVX1 U28302 ( .A(reg_file[2978]), .Y(n29193) );
  NOR2X1 U28303 ( .A(n26025), .B(n29151), .Y(n22149) );
  INVX1 U28304 ( .A(reg_file[2979]), .Y(n29151) );
  NOR2X1 U28305 ( .A(n26025), .B(n29109), .Y(n22148) );
  INVX1 U28306 ( .A(reg_file[2980]), .Y(n29109) );
  NOR2X1 U28307 ( .A(n26025), .B(n29067), .Y(n22147) );
  INVX1 U28308 ( .A(reg_file[2981]), .Y(n29067) );
  NOR2X1 U28309 ( .A(n26025), .B(n29025), .Y(n22146) );
  INVX1 U28310 ( .A(reg_file[2982]), .Y(n29025) );
  NOR2X1 U28311 ( .A(n26025), .B(n28983), .Y(n22145) );
  INVX1 U28312 ( .A(reg_file[2983]), .Y(n28983) );
  NOR2X1 U28313 ( .A(n26025), .B(n28899), .Y(n22144) );
  INVX1 U28314 ( .A(reg_file[2984]), .Y(n28899) );
  NOR2X1 U28315 ( .A(n26025), .B(n28857), .Y(n22143) );
  INVX1 U28316 ( .A(reg_file[2985]), .Y(n28857) );
  NOR2X1 U28317 ( .A(n26025), .B(n28815), .Y(n22142) );
  INVX1 U28318 ( .A(reg_file[2986]), .Y(n28815) );
  NOR2X1 U28319 ( .A(n26025), .B(n28773), .Y(n22141) );
  INVX1 U28320 ( .A(reg_file[2987]), .Y(n28773) );
  NOR2X1 U28321 ( .A(n26025), .B(n28731), .Y(n22140) );
  INVX1 U28322 ( .A(reg_file[2988]), .Y(n28731) );
  NOR2X1 U28323 ( .A(n26025), .B(n28689), .Y(n22139) );
  INVX1 U28324 ( .A(reg_file[2989]), .Y(n28689) );
  NOR2X1 U28325 ( .A(n26025), .B(n28647), .Y(n22138) );
  INVX1 U28326 ( .A(reg_file[2990]), .Y(n28647) );
  NOR2X1 U28327 ( .A(n26025), .B(n28605), .Y(n22137) );
  INVX1 U28328 ( .A(reg_file[2991]), .Y(n28605) );
  NOR2X1 U28329 ( .A(n26026), .B(n28563), .Y(n22136) );
  INVX1 U28330 ( .A(reg_file[2992]), .Y(n28563) );
  NOR2X1 U28331 ( .A(n26026), .B(n28521), .Y(n22135) );
  INVX1 U28332 ( .A(reg_file[2993]), .Y(n28521) );
  NOR2X1 U28333 ( .A(n26026), .B(n28437), .Y(n22134) );
  INVX1 U28334 ( .A(reg_file[2994]), .Y(n28437) );
  NOR2X1 U28335 ( .A(n26026), .B(n28395), .Y(n22133) );
  INVX1 U28336 ( .A(reg_file[2995]), .Y(n28395) );
  NOR2X1 U28337 ( .A(n26026), .B(n28353), .Y(n22132) );
  INVX1 U28338 ( .A(reg_file[2996]), .Y(n28353) );
  NOR2X1 U28339 ( .A(n26026), .B(n28311), .Y(n22131) );
  INVX1 U28340 ( .A(reg_file[2997]), .Y(n28311) );
  NOR2X1 U28341 ( .A(n26026), .B(n28269), .Y(n22130) );
  INVX1 U28342 ( .A(reg_file[2998]), .Y(n28269) );
  NOR2X1 U28343 ( .A(n26026), .B(n28227), .Y(n22129) );
  INVX1 U28344 ( .A(reg_file[2999]), .Y(n28227) );
  NOR2X1 U28345 ( .A(n26026), .B(n28185), .Y(n22128) );
  INVX1 U28346 ( .A(reg_file[3000]), .Y(n28185) );
  NOR2X1 U28347 ( .A(n26026), .B(n28143), .Y(n22127) );
  INVX1 U28348 ( .A(reg_file[3001]), .Y(n28143) );
  NOR2X1 U28349 ( .A(n26026), .B(n28101), .Y(n22126) );
  INVX1 U28350 ( .A(reg_file[3002]), .Y(n28101) );
  NOR2X1 U28351 ( .A(n26026), .B(n28059), .Y(n22125) );
  INVX1 U28352 ( .A(reg_file[3003]), .Y(n28059) );
  NOR2X1 U28353 ( .A(n26026), .B(n27975), .Y(n22124) );
  INVX1 U28354 ( .A(reg_file[3004]), .Y(n27975) );
  NOR2X1 U28355 ( .A(n26026), .B(n27933), .Y(n22123) );
  INVX1 U28356 ( .A(reg_file[3005]), .Y(n27933) );
  NOR2X1 U28357 ( .A(n26026), .B(n27891), .Y(n22122) );
  INVX1 U28358 ( .A(reg_file[3006]), .Y(n27891) );
  NOR2X1 U28359 ( .A(n26026), .B(n27849), .Y(n22121) );
  INVX1 U28360 ( .A(reg_file[3007]), .Y(n27849) );
  NOR2X1 U28361 ( .A(n26026), .B(n27807), .Y(n22120) );
  INVX1 U28362 ( .A(reg_file[3008]), .Y(n27807) );
  NOR2X1 U28363 ( .A(n26027), .B(n27765), .Y(n22119) );
  INVX1 U28364 ( .A(reg_file[3009]), .Y(n27765) );
  NOR2X1 U28365 ( .A(n26027), .B(n27723), .Y(n22118) );
  INVX1 U28366 ( .A(reg_file[3010]), .Y(n27723) );
  NOR2X1 U28367 ( .A(n26027), .B(n27681), .Y(n22117) );
  INVX1 U28368 ( .A(reg_file[3011]), .Y(n27681) );
  NOR2X1 U28369 ( .A(n26027), .B(n27639), .Y(n22116) );
  INVX1 U28370 ( .A(reg_file[3012]), .Y(n27639) );
  NOR2X1 U28371 ( .A(n26027), .B(n27597), .Y(n22115) );
  INVX1 U28372 ( .A(reg_file[3013]), .Y(n27597) );
  NOR2X1 U28373 ( .A(n26027), .B(n27513), .Y(n22114) );
  INVX1 U28374 ( .A(reg_file[3014]), .Y(n27513) );
  NOR2X1 U28375 ( .A(n26027), .B(n27471), .Y(n22113) );
  INVX1 U28376 ( .A(reg_file[3015]), .Y(n27471) );
  NOR2X1 U28377 ( .A(n26027), .B(n27429), .Y(n22112) );
  INVX1 U28378 ( .A(reg_file[3016]), .Y(n27429) );
  NOR2X1 U28379 ( .A(n26027), .B(n27387), .Y(n22111) );
  INVX1 U28380 ( .A(reg_file[3017]), .Y(n27387) );
  NOR2X1 U28381 ( .A(n26027), .B(n27345), .Y(n22110) );
  INVX1 U28382 ( .A(reg_file[3018]), .Y(n27345) );
  NOR2X1 U28383 ( .A(n26027), .B(n27303), .Y(n22109) );
  INVX1 U28384 ( .A(reg_file[3019]), .Y(n27303) );
  NOR2X1 U28385 ( .A(n26027), .B(n27261), .Y(n22108) );
  INVX1 U28386 ( .A(reg_file[3020]), .Y(n27261) );
  NOR2X1 U28387 ( .A(n26027), .B(n27219), .Y(n22107) );
  INVX1 U28388 ( .A(reg_file[3021]), .Y(n27219) );
  NOR2X1 U28389 ( .A(n26027), .B(n27177), .Y(n22106) );
  INVX1 U28390 ( .A(reg_file[3022]), .Y(n27177) );
  NOR2X1 U28391 ( .A(n26027), .B(n27135), .Y(n22105) );
  INVX1 U28392 ( .A(reg_file[3023]), .Y(n27135) );
  NOR2X1 U28393 ( .A(n26027), .B(n27051), .Y(n22104) );
  INVX1 U28394 ( .A(reg_file[3024]), .Y(n27051) );
  NOR2X1 U28395 ( .A(n26027), .B(n27009), .Y(n22103) );
  INVX1 U28396 ( .A(reg_file[3025]), .Y(n27009) );
  NOR2X1 U28397 ( .A(n26028), .B(n26967), .Y(n22102) );
  INVX1 U28398 ( .A(reg_file[3026]), .Y(n26967) );
  NOR2X1 U28399 ( .A(n26028), .B(n26925), .Y(n22101) );
  INVX1 U28400 ( .A(reg_file[3027]), .Y(n26925) );
  NOR2X1 U28401 ( .A(n26028), .B(n26883), .Y(n22100) );
  INVX1 U28402 ( .A(reg_file[3028]), .Y(n26883) );
  NOR2X1 U28403 ( .A(n26028), .B(n26841), .Y(n22099) );
  INVX1 U28404 ( .A(reg_file[3029]), .Y(n26841) );
  NOR2X1 U28405 ( .A(n26028), .B(n26799), .Y(n22098) );
  INVX1 U28406 ( .A(reg_file[3030]), .Y(n26799) );
  NOR2X1 U28407 ( .A(n26028), .B(n26757), .Y(n22097) );
  INVX1 U28408 ( .A(reg_file[3031]), .Y(n26757) );
  NOR2X1 U28409 ( .A(n26028), .B(n26715), .Y(n22096) );
  INVX1 U28410 ( .A(reg_file[3032]), .Y(n26715) );
  NOR2X1 U28411 ( .A(n26028), .B(n26673), .Y(n22095) );
  INVX1 U28412 ( .A(reg_file[3033]), .Y(n26673) );
  NOR2X1 U28413 ( .A(n26028), .B(n26589), .Y(n22094) );
  INVX1 U28414 ( .A(reg_file[3034]), .Y(n26589) );
  NOR2X1 U28415 ( .A(n26028), .B(n26547), .Y(n22093) );
  INVX1 U28416 ( .A(reg_file[3035]), .Y(n26547) );
  NOR2X1 U28417 ( .A(n26028), .B(n26505), .Y(n22092) );
  INVX1 U28418 ( .A(reg_file[3036]), .Y(n26505) );
  NOR2X1 U28419 ( .A(n26028), .B(n26463), .Y(n22091) );
  INVX1 U28420 ( .A(reg_file[3037]), .Y(n26463) );
  NOR2X1 U28421 ( .A(n26028), .B(n26421), .Y(n22090) );
  INVX1 U28422 ( .A(reg_file[3038]), .Y(n26421) );
  NOR2X1 U28423 ( .A(n26028), .B(n26379), .Y(n22089) );
  INVX1 U28424 ( .A(reg_file[3039]), .Y(n26379) );
  NOR2X1 U28425 ( .A(n26028), .B(n26337), .Y(n22088) );
  INVX1 U28426 ( .A(reg_file[3040]), .Y(n26337) );
  NOR2X1 U28427 ( .A(n26028), .B(n26295), .Y(n22087) );
  INVX1 U28428 ( .A(reg_file[3041]), .Y(n26295) );
  NOR2X1 U28429 ( .A(n26028), .B(n26253), .Y(n22086) );
  INVX1 U28430 ( .A(reg_file[3042]), .Y(n26253) );
  NOR2X1 U28431 ( .A(n26029), .B(n26211), .Y(n22085) );
  INVX1 U28432 ( .A(reg_file[3043]), .Y(n26211) );
  NOR2X1 U28433 ( .A(n26029), .B(n31461), .Y(n22084) );
  INVX1 U28434 ( .A(reg_file[3044]), .Y(n31461) );
  NOR2X1 U28435 ( .A(n26029), .B(n31419), .Y(n22083) );
  INVX1 U28436 ( .A(reg_file[3045]), .Y(n31419) );
  NOR2X1 U28437 ( .A(n26029), .B(n31377), .Y(n22082) );
  INVX1 U28438 ( .A(reg_file[3046]), .Y(n31377) );
  NOR2X1 U28439 ( .A(n26029), .B(n31335), .Y(n22081) );
  INVX1 U28440 ( .A(reg_file[3047]), .Y(n31335) );
  NOR2X1 U28441 ( .A(n26029), .B(n31293), .Y(n22080) );
  INVX1 U28442 ( .A(reg_file[3048]), .Y(n31293) );
  NOR2X1 U28443 ( .A(n26029), .B(n31251), .Y(n22079) );
  INVX1 U28444 ( .A(reg_file[3049]), .Y(n31251) );
  NOR2X1 U28445 ( .A(n26029), .B(n31209), .Y(n22078) );
  INVX1 U28446 ( .A(reg_file[3050]), .Y(n31209) );
  NOR2X1 U28447 ( .A(n26029), .B(n31167), .Y(n22077) );
  INVX1 U28448 ( .A(reg_file[3051]), .Y(n31167) );
  NOR2X1 U28449 ( .A(n26029), .B(n31125), .Y(n22076) );
  INVX1 U28450 ( .A(reg_file[3052]), .Y(n31125) );
  NOR2X1 U28451 ( .A(n26029), .B(n31083), .Y(n22075) );
  INVX1 U28452 ( .A(reg_file[3053]), .Y(n31083) );
  NOR2X1 U28453 ( .A(n26029), .B(n30999), .Y(n22074) );
  INVX1 U28454 ( .A(reg_file[3054]), .Y(n30999) );
  NOR2X1 U28455 ( .A(n26029), .B(n30957), .Y(n22073) );
  INVX1 U28456 ( .A(reg_file[3055]), .Y(n30957) );
  NOR2X1 U28457 ( .A(n26029), .B(n30915), .Y(n22072) );
  INVX1 U28458 ( .A(reg_file[3056]), .Y(n30915) );
  NOR2X1 U28459 ( .A(n26029), .B(n30873), .Y(n22071) );
  INVX1 U28460 ( .A(reg_file[3057]), .Y(n30873) );
  NOR2X1 U28461 ( .A(n26029), .B(n30831), .Y(n22070) );
  INVX1 U28462 ( .A(reg_file[3058]), .Y(n30831) );
  NOR2X1 U28463 ( .A(n26029), .B(n30789), .Y(n22069) );
  INVX1 U28464 ( .A(reg_file[3059]), .Y(n30789) );
  NOR2X1 U28465 ( .A(n26030), .B(n30747), .Y(n22068) );
  INVX1 U28466 ( .A(reg_file[3060]), .Y(n30747) );
  NOR2X1 U28467 ( .A(n26030), .B(n30705), .Y(n22067) );
  INVX1 U28468 ( .A(reg_file[3061]), .Y(n30705) );
  NOR2X1 U28469 ( .A(n26030), .B(n30663), .Y(n22066) );
  INVX1 U28470 ( .A(reg_file[3062]), .Y(n30663) );
  NOR2X1 U28471 ( .A(n26030), .B(n30621), .Y(n22065) );
  INVX1 U28472 ( .A(reg_file[3063]), .Y(n30621) );
  NOR2X1 U28473 ( .A(n26030), .B(n30537), .Y(n22064) );
  INVX1 U28474 ( .A(reg_file[3064]), .Y(n30537) );
  NOR2X1 U28475 ( .A(n26030), .B(n30495), .Y(n22063) );
  INVX1 U28476 ( .A(reg_file[3065]), .Y(n30495) );
  NOR2X1 U28477 ( .A(n26030), .B(n30453), .Y(n22062) );
  INVX1 U28478 ( .A(reg_file[3066]), .Y(n30453) );
  NOR2X1 U28479 ( .A(n26030), .B(n30411), .Y(n22061) );
  INVX1 U28480 ( .A(reg_file[3067]), .Y(n30411) );
  NOR2X1 U28481 ( .A(n26030), .B(n30369), .Y(n22060) );
  INVX1 U28482 ( .A(reg_file[3068]), .Y(n30369) );
  NOR2X1 U28483 ( .A(n26030), .B(n30327), .Y(n22059) );
  INVX1 U28484 ( .A(reg_file[3069]), .Y(n30327) );
  NOR2X1 U28485 ( .A(n26030), .B(n30285), .Y(n22058) );
  INVX1 U28486 ( .A(reg_file[3070]), .Y(n30285) );
  NOR2X1 U28487 ( .A(n26030), .B(n30243), .Y(n22057) );
  INVX1 U28488 ( .A(reg_file[3071]), .Y(n30243) );
  NOR2X1 U28489 ( .A(n36231), .B(n35317), .Y(n36493) );
  NAND3X1 U28490 ( .A(wraddr[0]), .B(n35318), .C(wraddr[4]), .Y(n36231) );
  INVX1 U28491 ( .A(wraddr[3]), .Y(n35318) );
  MUX2X1 U28492 ( .B(n36494), .A(n25129), .S(n26031), .Y(n22056) );
  INVX1 U28493 ( .A(reg_file[3072]), .Y(n36494) );
  MUX2X1 U28494 ( .B(n36496), .A(n25130), .S(n26031), .Y(n22055) );
  INVX1 U28495 ( .A(reg_file[3073]), .Y(n36496) );
  MUX2X1 U28496 ( .B(n36497), .A(n25131), .S(n26031), .Y(n22054) );
  INVX1 U28497 ( .A(reg_file[3074]), .Y(n36497) );
  MUX2X1 U28498 ( .B(n36498), .A(n25132), .S(n26031), .Y(n22053) );
  INVX1 U28499 ( .A(reg_file[3075]), .Y(n36498) );
  MUX2X1 U28500 ( .B(n36499), .A(n25133), .S(n26031), .Y(n22052) );
  INVX1 U28501 ( .A(reg_file[3076]), .Y(n36499) );
  MUX2X1 U28502 ( .B(n36500), .A(n25134), .S(n26031), .Y(n22051) );
  INVX1 U28503 ( .A(reg_file[3077]), .Y(n36500) );
  MUX2X1 U28504 ( .B(n36501), .A(n25135), .S(n26031), .Y(n22050) );
  INVX1 U28505 ( .A(reg_file[3078]), .Y(n36501) );
  MUX2X1 U28506 ( .B(n36502), .A(n25136), .S(n26031), .Y(n22049) );
  INVX1 U28507 ( .A(reg_file[3079]), .Y(n36502) );
  NOR2X1 U28508 ( .A(n26031), .B(n36503), .Y(n22048) );
  INVX1 U28509 ( .A(reg_file[3080]), .Y(n36503) );
  NOR2X1 U28510 ( .A(n26031), .B(n36504), .Y(n22047) );
  INVX1 U28511 ( .A(reg_file[3081]), .Y(n36504) );
  NOR2X1 U28512 ( .A(n26031), .B(n36505), .Y(n22046) );
  INVX1 U28513 ( .A(reg_file[3082]), .Y(n36505) );
  NOR2X1 U28514 ( .A(n26031), .B(n36506), .Y(n22045) );
  INVX1 U28515 ( .A(reg_file[3083]), .Y(n36506) );
  NOR2X1 U28516 ( .A(n26031), .B(n36507), .Y(n22044) );
  INVX1 U28517 ( .A(reg_file[3084]), .Y(n36507) );
  NOR2X1 U28518 ( .A(n26031), .B(n36508), .Y(n22043) );
  INVX1 U28519 ( .A(reg_file[3085]), .Y(n36508) );
  NOR2X1 U28520 ( .A(n26032), .B(n36509), .Y(n22042) );
  INVX1 U28521 ( .A(reg_file[3086]), .Y(n36509) );
  NOR2X1 U28522 ( .A(n26032), .B(n36510), .Y(n22041) );
  INVX1 U28523 ( .A(reg_file[3087]), .Y(n36510) );
  NOR2X1 U28524 ( .A(n26032), .B(n36511), .Y(n22040) );
  INVX1 U28525 ( .A(reg_file[3088]), .Y(n36511) );
  NOR2X1 U28526 ( .A(n26032), .B(n36512), .Y(n22039) );
  INVX1 U28527 ( .A(reg_file[3089]), .Y(n36512) );
  NOR2X1 U28528 ( .A(n26032), .B(n36513), .Y(n22038) );
  INVX1 U28529 ( .A(reg_file[3090]), .Y(n36513) );
  NOR2X1 U28530 ( .A(n26032), .B(n36514), .Y(n22037) );
  INVX1 U28531 ( .A(reg_file[3091]), .Y(n36514) );
  NOR2X1 U28532 ( .A(n26032), .B(n36515), .Y(n22036) );
  INVX1 U28533 ( .A(reg_file[3092]), .Y(n36515) );
  NOR2X1 U28534 ( .A(n26032), .B(n36516), .Y(n22035) );
  INVX1 U28535 ( .A(reg_file[3093]), .Y(n36516) );
  NOR2X1 U28536 ( .A(n26032), .B(n36517), .Y(n22034) );
  INVX1 U28537 ( .A(reg_file[3094]), .Y(n36517) );
  NOR2X1 U28538 ( .A(n26032), .B(n36518), .Y(n22033) );
  INVX1 U28539 ( .A(reg_file[3095]), .Y(n36518) );
  NOR2X1 U28540 ( .A(n26032), .B(n36519), .Y(n22032) );
  INVX1 U28541 ( .A(reg_file[3096]), .Y(n36519) );
  NOR2X1 U28542 ( .A(n26032), .B(n36520), .Y(n22031) );
  INVX1 U28543 ( .A(reg_file[3097]), .Y(n36520) );
  NOR2X1 U28544 ( .A(n26032), .B(n36521), .Y(n22030) );
  INVX1 U28545 ( .A(reg_file[3098]), .Y(n36521) );
  NOR2X1 U28546 ( .A(n26032), .B(n36522), .Y(n22029) );
  INVX1 U28547 ( .A(reg_file[3099]), .Y(n36522) );
  NOR2X1 U28548 ( .A(n26032), .B(n36523), .Y(n22028) );
  INVX1 U28549 ( .A(reg_file[3100]), .Y(n36523) );
  NOR2X1 U28550 ( .A(n26032), .B(n36524), .Y(n22027) );
  INVX1 U28551 ( .A(reg_file[3101]), .Y(n36524) );
  NOR2X1 U28552 ( .A(n26032), .B(n36525), .Y(n22026) );
  INVX1 U28553 ( .A(reg_file[3102]), .Y(n36525) );
  NOR2X1 U28554 ( .A(n26033), .B(n36526), .Y(n22025) );
  INVX1 U28555 ( .A(reg_file[3103]), .Y(n36526) );
  NOR2X1 U28556 ( .A(n26033), .B(n36527), .Y(n22024) );
  INVX1 U28557 ( .A(reg_file[3104]), .Y(n36527) );
  NOR2X1 U28558 ( .A(n26033), .B(n36528), .Y(n22023) );
  INVX1 U28559 ( .A(reg_file[3105]), .Y(n36528) );
  NOR2X1 U28560 ( .A(n26033), .B(n36529), .Y(n22022) );
  INVX1 U28561 ( .A(reg_file[3106]), .Y(n36529) );
  NOR2X1 U28562 ( .A(n26033), .B(n36530), .Y(n22021) );
  INVX1 U28563 ( .A(reg_file[3107]), .Y(n36530) );
  NOR2X1 U28564 ( .A(n26033), .B(n36531), .Y(n22020) );
  INVX1 U28565 ( .A(reg_file[3108]), .Y(n36531) );
  NOR2X1 U28566 ( .A(n26033), .B(n36532), .Y(n22019) );
  INVX1 U28567 ( .A(reg_file[3109]), .Y(n36532) );
  NOR2X1 U28568 ( .A(n26033), .B(n36533), .Y(n22018) );
  INVX1 U28569 ( .A(reg_file[3110]), .Y(n36533) );
  NOR2X1 U28570 ( .A(n26033), .B(n36534), .Y(n22017) );
  INVX1 U28571 ( .A(reg_file[3111]), .Y(n36534) );
  NOR2X1 U28572 ( .A(n26033), .B(n36535), .Y(n22016) );
  INVX1 U28573 ( .A(reg_file[3112]), .Y(n36535) );
  NOR2X1 U28574 ( .A(n26033), .B(n36536), .Y(n22015) );
  INVX1 U28575 ( .A(reg_file[3113]), .Y(n36536) );
  NOR2X1 U28576 ( .A(n26033), .B(n36537), .Y(n22014) );
  INVX1 U28577 ( .A(reg_file[3114]), .Y(n36537) );
  NOR2X1 U28578 ( .A(n26033), .B(n36538), .Y(n22013) );
  INVX1 U28579 ( .A(reg_file[3115]), .Y(n36538) );
  NOR2X1 U28580 ( .A(n26033), .B(n36539), .Y(n22012) );
  INVX1 U28581 ( .A(reg_file[3116]), .Y(n36539) );
  NOR2X1 U28582 ( .A(n26033), .B(n36540), .Y(n22011) );
  INVX1 U28583 ( .A(reg_file[3117]), .Y(n36540) );
  NOR2X1 U28584 ( .A(n26033), .B(n36541), .Y(n22010) );
  INVX1 U28585 ( .A(reg_file[3118]), .Y(n36541) );
  NOR2X1 U28586 ( .A(n26033), .B(n36542), .Y(n22009) );
  INVX1 U28587 ( .A(reg_file[3119]), .Y(n36542) );
  NOR2X1 U28588 ( .A(n26034), .B(n36543), .Y(n22008) );
  INVX1 U28589 ( .A(reg_file[3120]), .Y(n36543) );
  NOR2X1 U28590 ( .A(n26034), .B(n36544), .Y(n22007) );
  INVX1 U28591 ( .A(reg_file[3121]), .Y(n36544) );
  NOR2X1 U28592 ( .A(n26034), .B(n36545), .Y(n22006) );
  INVX1 U28593 ( .A(reg_file[3122]), .Y(n36545) );
  NOR2X1 U28594 ( .A(n26034), .B(n36546), .Y(n22005) );
  INVX1 U28595 ( .A(reg_file[3123]), .Y(n36546) );
  NOR2X1 U28596 ( .A(n26034), .B(n36547), .Y(n22004) );
  INVX1 U28597 ( .A(reg_file[3124]), .Y(n36547) );
  NOR2X1 U28598 ( .A(n26034), .B(n36548), .Y(n22003) );
  INVX1 U28599 ( .A(reg_file[3125]), .Y(n36548) );
  NOR2X1 U28600 ( .A(n26034), .B(n36549), .Y(n22002) );
  INVX1 U28601 ( .A(reg_file[3126]), .Y(n36549) );
  NOR2X1 U28602 ( .A(n26034), .B(n36550), .Y(n22001) );
  INVX1 U28603 ( .A(reg_file[3127]), .Y(n36550) );
  NOR2X1 U28604 ( .A(n26034), .B(n36551), .Y(n22000) );
  INVX1 U28605 ( .A(reg_file[3128]), .Y(n36551) );
  NOR2X1 U28606 ( .A(n26034), .B(n36552), .Y(n21999) );
  INVX1 U28607 ( .A(reg_file[3129]), .Y(n36552) );
  NOR2X1 U28608 ( .A(n26034), .B(n36553), .Y(n21998) );
  INVX1 U28609 ( .A(reg_file[3130]), .Y(n36553) );
  NOR2X1 U28610 ( .A(n26034), .B(n36554), .Y(n21997) );
  INVX1 U28611 ( .A(reg_file[3131]), .Y(n36554) );
  NOR2X1 U28612 ( .A(n26034), .B(n36555), .Y(n21996) );
  INVX1 U28613 ( .A(reg_file[3132]), .Y(n36555) );
  NOR2X1 U28614 ( .A(n26034), .B(n36556), .Y(n21995) );
  INVX1 U28615 ( .A(reg_file[3133]), .Y(n36556) );
  NOR2X1 U28616 ( .A(n26034), .B(n36557), .Y(n21994) );
  INVX1 U28617 ( .A(reg_file[3134]), .Y(n36557) );
  NOR2X1 U28618 ( .A(n26034), .B(n36558), .Y(n21993) );
  INVX1 U28619 ( .A(reg_file[3135]), .Y(n36558) );
  NOR2X1 U28620 ( .A(n26034), .B(n36559), .Y(n21992) );
  INVX1 U28621 ( .A(reg_file[3136]), .Y(n36559) );
  NOR2X1 U28622 ( .A(n26035), .B(n36560), .Y(n21991) );
  INVX1 U28623 ( .A(reg_file[3137]), .Y(n36560) );
  NOR2X1 U28624 ( .A(n26035), .B(n36561), .Y(n21990) );
  INVX1 U28625 ( .A(reg_file[3138]), .Y(n36561) );
  NOR2X1 U28626 ( .A(n26035), .B(n36562), .Y(n21989) );
  INVX1 U28627 ( .A(reg_file[3139]), .Y(n36562) );
  NOR2X1 U28628 ( .A(n26035), .B(n36563), .Y(n21988) );
  INVX1 U28629 ( .A(reg_file[3140]), .Y(n36563) );
  NOR2X1 U28630 ( .A(n26035), .B(n36564), .Y(n21987) );
  INVX1 U28631 ( .A(reg_file[3141]), .Y(n36564) );
  NOR2X1 U28632 ( .A(n26035), .B(n36565), .Y(n21986) );
  INVX1 U28633 ( .A(reg_file[3142]), .Y(n36565) );
  NOR2X1 U28634 ( .A(n26035), .B(n36566), .Y(n21985) );
  INVX1 U28635 ( .A(reg_file[3143]), .Y(n36566) );
  NOR2X1 U28636 ( .A(n26035), .B(n36567), .Y(n21984) );
  INVX1 U28637 ( .A(reg_file[3144]), .Y(n36567) );
  NOR2X1 U28638 ( .A(n26035), .B(n36568), .Y(n21983) );
  INVX1 U28639 ( .A(reg_file[3145]), .Y(n36568) );
  NOR2X1 U28640 ( .A(n26035), .B(n36569), .Y(n21982) );
  INVX1 U28641 ( .A(reg_file[3146]), .Y(n36569) );
  NOR2X1 U28642 ( .A(n26035), .B(n36570), .Y(n21981) );
  INVX1 U28643 ( .A(reg_file[3147]), .Y(n36570) );
  NOR2X1 U28644 ( .A(n26035), .B(n36571), .Y(n21980) );
  INVX1 U28645 ( .A(reg_file[3148]), .Y(n36571) );
  NOR2X1 U28646 ( .A(n26035), .B(n36572), .Y(n21979) );
  INVX1 U28647 ( .A(reg_file[3149]), .Y(n36572) );
  NOR2X1 U28648 ( .A(n26035), .B(n36573), .Y(n21978) );
  INVX1 U28649 ( .A(reg_file[3150]), .Y(n36573) );
  NOR2X1 U28650 ( .A(n26035), .B(n36574), .Y(n21977) );
  INVX1 U28651 ( .A(reg_file[3151]), .Y(n36574) );
  NOR2X1 U28652 ( .A(n26035), .B(n36575), .Y(n21976) );
  INVX1 U28653 ( .A(reg_file[3152]), .Y(n36575) );
  NOR2X1 U28654 ( .A(n26035), .B(n36576), .Y(n21975) );
  INVX1 U28655 ( .A(reg_file[3153]), .Y(n36576) );
  NOR2X1 U28656 ( .A(n26036), .B(n36577), .Y(n21974) );
  INVX1 U28657 ( .A(reg_file[3154]), .Y(n36577) );
  NOR2X1 U28658 ( .A(n26036), .B(n36578), .Y(n21973) );
  INVX1 U28659 ( .A(reg_file[3155]), .Y(n36578) );
  NOR2X1 U28660 ( .A(n26036), .B(n36579), .Y(n21972) );
  INVX1 U28661 ( .A(reg_file[3156]), .Y(n36579) );
  NOR2X1 U28662 ( .A(n26036), .B(n36580), .Y(n21971) );
  INVX1 U28663 ( .A(reg_file[3157]), .Y(n36580) );
  NOR2X1 U28664 ( .A(n26036), .B(n36581), .Y(n21970) );
  INVX1 U28665 ( .A(reg_file[3158]), .Y(n36581) );
  NOR2X1 U28666 ( .A(n26036), .B(n36582), .Y(n21969) );
  INVX1 U28667 ( .A(reg_file[3159]), .Y(n36582) );
  NOR2X1 U28668 ( .A(n26036), .B(n36583), .Y(n21968) );
  INVX1 U28669 ( .A(reg_file[3160]), .Y(n36583) );
  NOR2X1 U28670 ( .A(n26036), .B(n36584), .Y(n21967) );
  INVX1 U28671 ( .A(reg_file[3161]), .Y(n36584) );
  NOR2X1 U28672 ( .A(n26036), .B(n36585), .Y(n21966) );
  INVX1 U28673 ( .A(reg_file[3162]), .Y(n36585) );
  NOR2X1 U28674 ( .A(n26036), .B(n36586), .Y(n21965) );
  INVX1 U28675 ( .A(reg_file[3163]), .Y(n36586) );
  NOR2X1 U28676 ( .A(n26036), .B(n36587), .Y(n21964) );
  INVX1 U28677 ( .A(reg_file[3164]), .Y(n36587) );
  NOR2X1 U28678 ( .A(n26036), .B(n36588), .Y(n21963) );
  INVX1 U28679 ( .A(reg_file[3165]), .Y(n36588) );
  NOR2X1 U28680 ( .A(n26036), .B(n36589), .Y(n21962) );
  INVX1 U28681 ( .A(reg_file[3166]), .Y(n36589) );
  NOR2X1 U28682 ( .A(n26036), .B(n36590), .Y(n21961) );
  INVX1 U28683 ( .A(reg_file[3167]), .Y(n36590) );
  NOR2X1 U28684 ( .A(n26036), .B(n36591), .Y(n21960) );
  INVX1 U28685 ( .A(reg_file[3168]), .Y(n36591) );
  NOR2X1 U28686 ( .A(n26036), .B(n36592), .Y(n21959) );
  INVX1 U28687 ( .A(reg_file[3169]), .Y(n36592) );
  NOR2X1 U28688 ( .A(n26036), .B(n36593), .Y(n21958) );
  INVX1 U28689 ( .A(reg_file[3170]), .Y(n36593) );
  NOR2X1 U28690 ( .A(n26037), .B(n36594), .Y(n21957) );
  INVX1 U28691 ( .A(reg_file[3171]), .Y(n36594) );
  NOR2X1 U28692 ( .A(n26037), .B(n36595), .Y(n21956) );
  INVX1 U28693 ( .A(reg_file[3172]), .Y(n36595) );
  NOR2X1 U28694 ( .A(n26037), .B(n36596), .Y(n21955) );
  INVX1 U28695 ( .A(reg_file[3173]), .Y(n36596) );
  NOR2X1 U28696 ( .A(n26037), .B(n36597), .Y(n21954) );
  INVX1 U28697 ( .A(reg_file[3174]), .Y(n36597) );
  NOR2X1 U28698 ( .A(n26037), .B(n36598), .Y(n21953) );
  INVX1 U28699 ( .A(reg_file[3175]), .Y(n36598) );
  NOR2X1 U28700 ( .A(n26037), .B(n36599), .Y(n21952) );
  INVX1 U28701 ( .A(reg_file[3176]), .Y(n36599) );
  NOR2X1 U28702 ( .A(n26037), .B(n36600), .Y(n21951) );
  INVX1 U28703 ( .A(reg_file[3177]), .Y(n36600) );
  NOR2X1 U28704 ( .A(n26037), .B(n36601), .Y(n21950) );
  INVX1 U28705 ( .A(reg_file[3178]), .Y(n36601) );
  NOR2X1 U28706 ( .A(n26037), .B(n36602), .Y(n21949) );
  INVX1 U28707 ( .A(reg_file[3179]), .Y(n36602) );
  NOR2X1 U28708 ( .A(n26037), .B(n36603), .Y(n21948) );
  INVX1 U28709 ( .A(reg_file[3180]), .Y(n36603) );
  NOR2X1 U28710 ( .A(n26037), .B(n36604), .Y(n21947) );
  INVX1 U28711 ( .A(reg_file[3181]), .Y(n36604) );
  NOR2X1 U28712 ( .A(n26037), .B(n36605), .Y(n21946) );
  INVX1 U28713 ( .A(reg_file[3182]), .Y(n36605) );
  NOR2X1 U28714 ( .A(n26037), .B(n36606), .Y(n21945) );
  INVX1 U28715 ( .A(reg_file[3183]), .Y(n36606) );
  NOR2X1 U28716 ( .A(n26037), .B(n36607), .Y(n21944) );
  INVX1 U28717 ( .A(reg_file[3184]), .Y(n36607) );
  NOR2X1 U28718 ( .A(n26037), .B(n36608), .Y(n21943) );
  INVX1 U28719 ( .A(reg_file[3185]), .Y(n36608) );
  NOR2X1 U28720 ( .A(n26037), .B(n36609), .Y(n21942) );
  INVX1 U28721 ( .A(reg_file[3186]), .Y(n36609) );
  NOR2X1 U28722 ( .A(n26037), .B(n36610), .Y(n21941) );
  INVX1 U28723 ( .A(reg_file[3187]), .Y(n36610) );
  NOR2X1 U28724 ( .A(n26038), .B(n36611), .Y(n21940) );
  INVX1 U28725 ( .A(reg_file[3188]), .Y(n36611) );
  NOR2X1 U28726 ( .A(n26038), .B(n36612), .Y(n21939) );
  INVX1 U28727 ( .A(reg_file[3189]), .Y(n36612) );
  NOR2X1 U28728 ( .A(n26038), .B(n36613), .Y(n21938) );
  INVX1 U28729 ( .A(reg_file[3190]), .Y(n36613) );
  NOR2X1 U28730 ( .A(n26038), .B(n36614), .Y(n21937) );
  INVX1 U28731 ( .A(reg_file[3191]), .Y(n36614) );
  NOR2X1 U28732 ( .A(n26038), .B(n36615), .Y(n21936) );
  INVX1 U28733 ( .A(reg_file[3192]), .Y(n36615) );
  NOR2X1 U28734 ( .A(n26038), .B(n36616), .Y(n21935) );
  INVX1 U28735 ( .A(reg_file[3193]), .Y(n36616) );
  NOR2X1 U28736 ( .A(n26038), .B(n36617), .Y(n21934) );
  INVX1 U28737 ( .A(reg_file[3194]), .Y(n36617) );
  NOR2X1 U28738 ( .A(n26038), .B(n36618), .Y(n21933) );
  INVX1 U28739 ( .A(reg_file[3195]), .Y(n36618) );
  NOR2X1 U28740 ( .A(n26038), .B(n36619), .Y(n21932) );
  INVX1 U28741 ( .A(reg_file[3196]), .Y(n36619) );
  NOR2X1 U28742 ( .A(n26038), .B(n36620), .Y(n21931) );
  INVX1 U28743 ( .A(reg_file[3197]), .Y(n36620) );
  NOR2X1 U28744 ( .A(n26038), .B(n36621), .Y(n21930) );
  INVX1 U28745 ( .A(reg_file[3198]), .Y(n36621) );
  NOR2X1 U28746 ( .A(n26038), .B(n36622), .Y(n21929) );
  INVX1 U28747 ( .A(reg_file[3199]), .Y(n36622) );
  NOR2X1 U28748 ( .A(n36623), .B(n34923), .Y(n36495) );
  MUX2X1 U28749 ( .B(n36624), .A(n25129), .S(n26039), .Y(n21928) );
  INVX1 U28750 ( .A(reg_file[3200]), .Y(n36624) );
  MUX2X1 U28751 ( .B(n36626), .A(n25130), .S(n26039), .Y(n21927) );
  INVX1 U28752 ( .A(reg_file[3201]), .Y(n36626) );
  MUX2X1 U28753 ( .B(n36627), .A(n25131), .S(n26039), .Y(n21926) );
  INVX1 U28754 ( .A(reg_file[3202]), .Y(n36627) );
  MUX2X1 U28755 ( .B(n36628), .A(n25132), .S(n26039), .Y(n21925) );
  INVX1 U28756 ( .A(reg_file[3203]), .Y(n36628) );
  MUX2X1 U28757 ( .B(n36629), .A(n25133), .S(n26039), .Y(n21924) );
  INVX1 U28758 ( .A(reg_file[3204]), .Y(n36629) );
  MUX2X1 U28759 ( .B(n36630), .A(n25134), .S(n26039), .Y(n21923) );
  INVX1 U28760 ( .A(reg_file[3205]), .Y(n36630) );
  MUX2X1 U28761 ( .B(n36631), .A(n25135), .S(n26039), .Y(n21922) );
  INVX1 U28762 ( .A(reg_file[3206]), .Y(n36631) );
  MUX2X1 U28763 ( .B(n36632), .A(n25136), .S(n26039), .Y(n21921) );
  INVX1 U28764 ( .A(reg_file[3207]), .Y(n36632) );
  NOR2X1 U28765 ( .A(n26039), .B(n36633), .Y(n21920) );
  INVX1 U28766 ( .A(reg_file[3208]), .Y(n36633) );
  NOR2X1 U28767 ( .A(n26039), .B(n36634), .Y(n21919) );
  INVX1 U28768 ( .A(reg_file[3209]), .Y(n36634) );
  NOR2X1 U28769 ( .A(n26039), .B(n36635), .Y(n21918) );
  INVX1 U28770 ( .A(reg_file[3210]), .Y(n36635) );
  NOR2X1 U28771 ( .A(n26039), .B(n36636), .Y(n21917) );
  INVX1 U28772 ( .A(reg_file[3211]), .Y(n36636) );
  NOR2X1 U28773 ( .A(n26039), .B(n36637), .Y(n21916) );
  INVX1 U28774 ( .A(reg_file[3212]), .Y(n36637) );
  NOR2X1 U28775 ( .A(n26039), .B(n36638), .Y(n21915) );
  INVX1 U28776 ( .A(reg_file[3213]), .Y(n36638) );
  NOR2X1 U28777 ( .A(n26040), .B(n36639), .Y(n21914) );
  INVX1 U28778 ( .A(reg_file[3214]), .Y(n36639) );
  NOR2X1 U28779 ( .A(n26040), .B(n36640), .Y(n21913) );
  INVX1 U28780 ( .A(reg_file[3215]), .Y(n36640) );
  NOR2X1 U28781 ( .A(n26040), .B(n36641), .Y(n21912) );
  INVX1 U28782 ( .A(reg_file[3216]), .Y(n36641) );
  NOR2X1 U28783 ( .A(n26040), .B(n36642), .Y(n21911) );
  INVX1 U28784 ( .A(reg_file[3217]), .Y(n36642) );
  NOR2X1 U28785 ( .A(n26040), .B(n36643), .Y(n21910) );
  INVX1 U28786 ( .A(reg_file[3218]), .Y(n36643) );
  NOR2X1 U28787 ( .A(n26040), .B(n36644), .Y(n21909) );
  INVX1 U28788 ( .A(reg_file[3219]), .Y(n36644) );
  NOR2X1 U28789 ( .A(n26040), .B(n36645), .Y(n21908) );
  INVX1 U28790 ( .A(reg_file[3220]), .Y(n36645) );
  NOR2X1 U28791 ( .A(n26040), .B(n36646), .Y(n21907) );
  INVX1 U28792 ( .A(reg_file[3221]), .Y(n36646) );
  NOR2X1 U28793 ( .A(n26040), .B(n36647), .Y(n21906) );
  INVX1 U28794 ( .A(reg_file[3222]), .Y(n36647) );
  NOR2X1 U28795 ( .A(n26040), .B(n36648), .Y(n21905) );
  INVX1 U28796 ( .A(reg_file[3223]), .Y(n36648) );
  NOR2X1 U28797 ( .A(n26040), .B(n36649), .Y(n21904) );
  INVX1 U28798 ( .A(reg_file[3224]), .Y(n36649) );
  NOR2X1 U28799 ( .A(n26040), .B(n36650), .Y(n21903) );
  INVX1 U28800 ( .A(reg_file[3225]), .Y(n36650) );
  NOR2X1 U28801 ( .A(n26040), .B(n36651), .Y(n21902) );
  INVX1 U28802 ( .A(reg_file[3226]), .Y(n36651) );
  NOR2X1 U28803 ( .A(n26040), .B(n36652), .Y(n21901) );
  INVX1 U28804 ( .A(reg_file[3227]), .Y(n36652) );
  NOR2X1 U28805 ( .A(n26040), .B(n36653), .Y(n21900) );
  INVX1 U28806 ( .A(reg_file[3228]), .Y(n36653) );
  NOR2X1 U28807 ( .A(n26040), .B(n36654), .Y(n21899) );
  INVX1 U28808 ( .A(reg_file[3229]), .Y(n36654) );
  NOR2X1 U28809 ( .A(n26040), .B(n36655), .Y(n21898) );
  INVX1 U28810 ( .A(reg_file[3230]), .Y(n36655) );
  NOR2X1 U28811 ( .A(n26041), .B(n36656), .Y(n21897) );
  INVX1 U28812 ( .A(reg_file[3231]), .Y(n36656) );
  NOR2X1 U28813 ( .A(n26041), .B(n36657), .Y(n21896) );
  INVX1 U28814 ( .A(reg_file[3232]), .Y(n36657) );
  NOR2X1 U28815 ( .A(n26041), .B(n36658), .Y(n21895) );
  INVX1 U28816 ( .A(reg_file[3233]), .Y(n36658) );
  NOR2X1 U28817 ( .A(n26041), .B(n36659), .Y(n21894) );
  INVX1 U28818 ( .A(reg_file[3234]), .Y(n36659) );
  NOR2X1 U28819 ( .A(n26041), .B(n36660), .Y(n21893) );
  INVX1 U28820 ( .A(reg_file[3235]), .Y(n36660) );
  NOR2X1 U28821 ( .A(n26041), .B(n36661), .Y(n21892) );
  INVX1 U28822 ( .A(reg_file[3236]), .Y(n36661) );
  NOR2X1 U28823 ( .A(n26041), .B(n36662), .Y(n21891) );
  INVX1 U28824 ( .A(reg_file[3237]), .Y(n36662) );
  NOR2X1 U28825 ( .A(n26041), .B(n36663), .Y(n21890) );
  INVX1 U28826 ( .A(reg_file[3238]), .Y(n36663) );
  NOR2X1 U28827 ( .A(n26041), .B(n36664), .Y(n21889) );
  INVX1 U28828 ( .A(reg_file[3239]), .Y(n36664) );
  NOR2X1 U28829 ( .A(n26041), .B(n36665), .Y(n21888) );
  INVX1 U28830 ( .A(reg_file[3240]), .Y(n36665) );
  NOR2X1 U28831 ( .A(n26041), .B(n36666), .Y(n21887) );
  INVX1 U28832 ( .A(reg_file[3241]), .Y(n36666) );
  NOR2X1 U28833 ( .A(n26041), .B(n36667), .Y(n21886) );
  INVX1 U28834 ( .A(reg_file[3242]), .Y(n36667) );
  NOR2X1 U28835 ( .A(n26041), .B(n36668), .Y(n21885) );
  INVX1 U28836 ( .A(reg_file[3243]), .Y(n36668) );
  NOR2X1 U28837 ( .A(n26041), .B(n36669), .Y(n21884) );
  INVX1 U28838 ( .A(reg_file[3244]), .Y(n36669) );
  NOR2X1 U28839 ( .A(n26041), .B(n36670), .Y(n21883) );
  INVX1 U28840 ( .A(reg_file[3245]), .Y(n36670) );
  NOR2X1 U28841 ( .A(n26041), .B(n36671), .Y(n21882) );
  INVX1 U28842 ( .A(reg_file[3246]), .Y(n36671) );
  NOR2X1 U28843 ( .A(n26041), .B(n36672), .Y(n21881) );
  INVX1 U28844 ( .A(reg_file[3247]), .Y(n36672) );
  NOR2X1 U28845 ( .A(n26042), .B(n36673), .Y(n21880) );
  INVX1 U28846 ( .A(reg_file[3248]), .Y(n36673) );
  NOR2X1 U28847 ( .A(n26042), .B(n36674), .Y(n21879) );
  INVX1 U28848 ( .A(reg_file[3249]), .Y(n36674) );
  NOR2X1 U28849 ( .A(n26042), .B(n36675), .Y(n21878) );
  INVX1 U28850 ( .A(reg_file[3250]), .Y(n36675) );
  NOR2X1 U28851 ( .A(n26042), .B(n36676), .Y(n21877) );
  INVX1 U28852 ( .A(reg_file[3251]), .Y(n36676) );
  NOR2X1 U28853 ( .A(n26042), .B(n36677), .Y(n21876) );
  INVX1 U28854 ( .A(reg_file[3252]), .Y(n36677) );
  NOR2X1 U28855 ( .A(n26042), .B(n36678), .Y(n21875) );
  INVX1 U28856 ( .A(reg_file[3253]), .Y(n36678) );
  NOR2X1 U28857 ( .A(n26042), .B(n36679), .Y(n21874) );
  INVX1 U28858 ( .A(reg_file[3254]), .Y(n36679) );
  NOR2X1 U28859 ( .A(n26042), .B(n36680), .Y(n21873) );
  INVX1 U28860 ( .A(reg_file[3255]), .Y(n36680) );
  NOR2X1 U28861 ( .A(n26042), .B(n36681), .Y(n21872) );
  INVX1 U28862 ( .A(reg_file[3256]), .Y(n36681) );
  NOR2X1 U28863 ( .A(n26042), .B(n36682), .Y(n21871) );
  INVX1 U28864 ( .A(reg_file[3257]), .Y(n36682) );
  NOR2X1 U28865 ( .A(n26042), .B(n36683), .Y(n21870) );
  INVX1 U28866 ( .A(reg_file[3258]), .Y(n36683) );
  NOR2X1 U28867 ( .A(n26042), .B(n36684), .Y(n21869) );
  INVX1 U28868 ( .A(reg_file[3259]), .Y(n36684) );
  NOR2X1 U28869 ( .A(n26042), .B(n36685), .Y(n21868) );
  INVX1 U28870 ( .A(reg_file[3260]), .Y(n36685) );
  NOR2X1 U28871 ( .A(n26042), .B(n36686), .Y(n21867) );
  INVX1 U28872 ( .A(reg_file[3261]), .Y(n36686) );
  NOR2X1 U28873 ( .A(n26042), .B(n36687), .Y(n21866) );
  INVX1 U28874 ( .A(reg_file[3262]), .Y(n36687) );
  NOR2X1 U28875 ( .A(n26042), .B(n36688), .Y(n21865) );
  INVX1 U28876 ( .A(reg_file[3263]), .Y(n36688) );
  NOR2X1 U28877 ( .A(n26042), .B(n36689), .Y(n21864) );
  INVX1 U28878 ( .A(reg_file[3264]), .Y(n36689) );
  NOR2X1 U28879 ( .A(n26043), .B(n36690), .Y(n21863) );
  INVX1 U28880 ( .A(reg_file[3265]), .Y(n36690) );
  NOR2X1 U28881 ( .A(n26043), .B(n36691), .Y(n21862) );
  INVX1 U28882 ( .A(reg_file[3266]), .Y(n36691) );
  NOR2X1 U28883 ( .A(n26043), .B(n36692), .Y(n21861) );
  INVX1 U28884 ( .A(reg_file[3267]), .Y(n36692) );
  NOR2X1 U28885 ( .A(n26043), .B(n36693), .Y(n21860) );
  INVX1 U28886 ( .A(reg_file[3268]), .Y(n36693) );
  NOR2X1 U28887 ( .A(n26043), .B(n36694), .Y(n21859) );
  INVX1 U28888 ( .A(reg_file[3269]), .Y(n36694) );
  NOR2X1 U28889 ( .A(n26043), .B(n36695), .Y(n21858) );
  INVX1 U28890 ( .A(reg_file[3270]), .Y(n36695) );
  NOR2X1 U28891 ( .A(n26043), .B(n36696), .Y(n21857) );
  INVX1 U28892 ( .A(reg_file[3271]), .Y(n36696) );
  NOR2X1 U28893 ( .A(n26043), .B(n36697), .Y(n21856) );
  INVX1 U28894 ( .A(reg_file[3272]), .Y(n36697) );
  NOR2X1 U28895 ( .A(n26043), .B(n36698), .Y(n21855) );
  INVX1 U28896 ( .A(reg_file[3273]), .Y(n36698) );
  NOR2X1 U28897 ( .A(n26043), .B(n36699), .Y(n21854) );
  INVX1 U28898 ( .A(reg_file[3274]), .Y(n36699) );
  NOR2X1 U28899 ( .A(n26043), .B(n36700), .Y(n21853) );
  INVX1 U28900 ( .A(reg_file[3275]), .Y(n36700) );
  NOR2X1 U28901 ( .A(n26043), .B(n36701), .Y(n21852) );
  INVX1 U28902 ( .A(reg_file[3276]), .Y(n36701) );
  NOR2X1 U28903 ( .A(n26043), .B(n36702), .Y(n21851) );
  INVX1 U28904 ( .A(reg_file[3277]), .Y(n36702) );
  NOR2X1 U28905 ( .A(n26043), .B(n36703), .Y(n21850) );
  INVX1 U28906 ( .A(reg_file[3278]), .Y(n36703) );
  NOR2X1 U28907 ( .A(n26043), .B(n36704), .Y(n21849) );
  INVX1 U28908 ( .A(reg_file[3279]), .Y(n36704) );
  NOR2X1 U28909 ( .A(n26043), .B(n36705), .Y(n21848) );
  INVX1 U28910 ( .A(reg_file[3280]), .Y(n36705) );
  NOR2X1 U28911 ( .A(n26043), .B(n36706), .Y(n21847) );
  INVX1 U28912 ( .A(reg_file[3281]), .Y(n36706) );
  NOR2X1 U28913 ( .A(n26044), .B(n36707), .Y(n21846) );
  INVX1 U28914 ( .A(reg_file[3282]), .Y(n36707) );
  NOR2X1 U28915 ( .A(n26044), .B(n36708), .Y(n21845) );
  INVX1 U28916 ( .A(reg_file[3283]), .Y(n36708) );
  NOR2X1 U28917 ( .A(n26044), .B(n36709), .Y(n21844) );
  INVX1 U28918 ( .A(reg_file[3284]), .Y(n36709) );
  NOR2X1 U28919 ( .A(n26044), .B(n36710), .Y(n21843) );
  INVX1 U28920 ( .A(reg_file[3285]), .Y(n36710) );
  NOR2X1 U28921 ( .A(n26044), .B(n36711), .Y(n21842) );
  INVX1 U28922 ( .A(reg_file[3286]), .Y(n36711) );
  NOR2X1 U28923 ( .A(n26044), .B(n36712), .Y(n21841) );
  INVX1 U28924 ( .A(reg_file[3287]), .Y(n36712) );
  NOR2X1 U28925 ( .A(n26044), .B(n36713), .Y(n21840) );
  INVX1 U28926 ( .A(reg_file[3288]), .Y(n36713) );
  NOR2X1 U28927 ( .A(n26044), .B(n36714), .Y(n21839) );
  INVX1 U28928 ( .A(reg_file[3289]), .Y(n36714) );
  NOR2X1 U28929 ( .A(n26044), .B(n36715), .Y(n21838) );
  INVX1 U28930 ( .A(reg_file[3290]), .Y(n36715) );
  NOR2X1 U28931 ( .A(n26044), .B(n36716), .Y(n21837) );
  INVX1 U28932 ( .A(reg_file[3291]), .Y(n36716) );
  NOR2X1 U28933 ( .A(n26044), .B(n36717), .Y(n21836) );
  INVX1 U28934 ( .A(reg_file[3292]), .Y(n36717) );
  NOR2X1 U28935 ( .A(n26044), .B(n36718), .Y(n21835) );
  INVX1 U28936 ( .A(reg_file[3293]), .Y(n36718) );
  NOR2X1 U28937 ( .A(n26044), .B(n36719), .Y(n21834) );
  INVX1 U28938 ( .A(reg_file[3294]), .Y(n36719) );
  NOR2X1 U28939 ( .A(n26044), .B(n36720), .Y(n21833) );
  INVX1 U28940 ( .A(reg_file[3295]), .Y(n36720) );
  NOR2X1 U28941 ( .A(n26044), .B(n36721), .Y(n21832) );
  INVX1 U28942 ( .A(reg_file[3296]), .Y(n36721) );
  NOR2X1 U28943 ( .A(n26044), .B(n36722), .Y(n21831) );
  INVX1 U28944 ( .A(reg_file[3297]), .Y(n36722) );
  NOR2X1 U28945 ( .A(n26044), .B(n36723), .Y(n21830) );
  INVX1 U28946 ( .A(reg_file[3298]), .Y(n36723) );
  NOR2X1 U28947 ( .A(n26045), .B(n36724), .Y(n21829) );
  INVX1 U28948 ( .A(reg_file[3299]), .Y(n36724) );
  NOR2X1 U28949 ( .A(n26045), .B(n36725), .Y(n21828) );
  INVX1 U28950 ( .A(reg_file[3300]), .Y(n36725) );
  NOR2X1 U28951 ( .A(n26045), .B(n36726), .Y(n21827) );
  INVX1 U28952 ( .A(reg_file[3301]), .Y(n36726) );
  NOR2X1 U28953 ( .A(n26045), .B(n36727), .Y(n21826) );
  INVX1 U28954 ( .A(reg_file[3302]), .Y(n36727) );
  NOR2X1 U28955 ( .A(n26045), .B(n36728), .Y(n21825) );
  INVX1 U28956 ( .A(reg_file[3303]), .Y(n36728) );
  NOR2X1 U28957 ( .A(n26045), .B(n36729), .Y(n21824) );
  INVX1 U28958 ( .A(reg_file[3304]), .Y(n36729) );
  NOR2X1 U28959 ( .A(n26045), .B(n36730), .Y(n21823) );
  INVX1 U28960 ( .A(reg_file[3305]), .Y(n36730) );
  NOR2X1 U28961 ( .A(n26045), .B(n36731), .Y(n21822) );
  INVX1 U28962 ( .A(reg_file[3306]), .Y(n36731) );
  NOR2X1 U28963 ( .A(n26045), .B(n36732), .Y(n21821) );
  INVX1 U28964 ( .A(reg_file[3307]), .Y(n36732) );
  NOR2X1 U28965 ( .A(n26045), .B(n36733), .Y(n21820) );
  INVX1 U28966 ( .A(reg_file[3308]), .Y(n36733) );
  NOR2X1 U28967 ( .A(n26045), .B(n36734), .Y(n21819) );
  INVX1 U28968 ( .A(reg_file[3309]), .Y(n36734) );
  NOR2X1 U28969 ( .A(n26045), .B(n36735), .Y(n21818) );
  INVX1 U28970 ( .A(reg_file[3310]), .Y(n36735) );
  NOR2X1 U28971 ( .A(n26045), .B(n36736), .Y(n21817) );
  INVX1 U28972 ( .A(reg_file[3311]), .Y(n36736) );
  NOR2X1 U28973 ( .A(n26045), .B(n36737), .Y(n21816) );
  INVX1 U28974 ( .A(reg_file[3312]), .Y(n36737) );
  NOR2X1 U28975 ( .A(n26045), .B(n36738), .Y(n21815) );
  INVX1 U28976 ( .A(reg_file[3313]), .Y(n36738) );
  NOR2X1 U28977 ( .A(n26045), .B(n36739), .Y(n21814) );
  INVX1 U28978 ( .A(reg_file[3314]), .Y(n36739) );
  NOR2X1 U28979 ( .A(n26045), .B(n36740), .Y(n21813) );
  INVX1 U28980 ( .A(reg_file[3315]), .Y(n36740) );
  NOR2X1 U28981 ( .A(n26046), .B(n36741), .Y(n21812) );
  INVX1 U28982 ( .A(reg_file[3316]), .Y(n36741) );
  NOR2X1 U28983 ( .A(n26046), .B(n36742), .Y(n21811) );
  INVX1 U28984 ( .A(reg_file[3317]), .Y(n36742) );
  NOR2X1 U28985 ( .A(n26046), .B(n36743), .Y(n21810) );
  INVX1 U28986 ( .A(reg_file[3318]), .Y(n36743) );
  NOR2X1 U28987 ( .A(n26046), .B(n36744), .Y(n21809) );
  INVX1 U28988 ( .A(reg_file[3319]), .Y(n36744) );
  NOR2X1 U28989 ( .A(n26046), .B(n36745), .Y(n21808) );
  INVX1 U28990 ( .A(reg_file[3320]), .Y(n36745) );
  NOR2X1 U28991 ( .A(n26046), .B(n36746), .Y(n21807) );
  INVX1 U28992 ( .A(reg_file[3321]), .Y(n36746) );
  NOR2X1 U28993 ( .A(n26046), .B(n36747), .Y(n21806) );
  INVX1 U28994 ( .A(reg_file[3322]), .Y(n36747) );
  NOR2X1 U28995 ( .A(n26046), .B(n36748), .Y(n21805) );
  INVX1 U28996 ( .A(reg_file[3323]), .Y(n36748) );
  NOR2X1 U28997 ( .A(n26046), .B(n36749), .Y(n21804) );
  INVX1 U28998 ( .A(reg_file[3324]), .Y(n36749) );
  NOR2X1 U28999 ( .A(n26046), .B(n36750), .Y(n21803) );
  INVX1 U29000 ( .A(reg_file[3325]), .Y(n36750) );
  NOR2X1 U29001 ( .A(n26046), .B(n36751), .Y(n21802) );
  INVX1 U29002 ( .A(reg_file[3326]), .Y(n36751) );
  NOR2X1 U29003 ( .A(n26046), .B(n36752), .Y(n21801) );
  INVX1 U29004 ( .A(reg_file[3327]), .Y(n36752) );
  NOR2X1 U29005 ( .A(n36753), .B(n34923), .Y(n36625) );
  NAND3X1 U29006 ( .A(n36754), .B(n36755), .C(n36756), .Y(n34923) );
  MUX2X1 U29007 ( .B(n36757), .A(n25129), .S(n26047), .Y(n21800) );
  INVX1 U29008 ( .A(reg_file[3328]), .Y(n36757) );
  MUX2X1 U29009 ( .B(n36759), .A(n25130), .S(n26047), .Y(n21799) );
  INVX1 U29010 ( .A(reg_file[3329]), .Y(n36759) );
  MUX2X1 U29011 ( .B(n36760), .A(n25131), .S(n26047), .Y(n21798) );
  INVX1 U29012 ( .A(reg_file[3330]), .Y(n36760) );
  MUX2X1 U29013 ( .B(n36761), .A(n25132), .S(n26047), .Y(n21797) );
  INVX1 U29014 ( .A(reg_file[3331]), .Y(n36761) );
  MUX2X1 U29015 ( .B(n36762), .A(n25133), .S(n26047), .Y(n21796) );
  INVX1 U29016 ( .A(reg_file[3332]), .Y(n36762) );
  MUX2X1 U29017 ( .B(n36763), .A(n25134), .S(n26047), .Y(n21795) );
  INVX1 U29018 ( .A(reg_file[3333]), .Y(n36763) );
  MUX2X1 U29019 ( .B(n36764), .A(n25135), .S(n26047), .Y(n21794) );
  INVX1 U29020 ( .A(reg_file[3334]), .Y(n36764) );
  MUX2X1 U29021 ( .B(n36765), .A(n25136), .S(n26047), .Y(n21793) );
  INVX1 U29022 ( .A(reg_file[3335]), .Y(n36765) );
  NOR2X1 U29023 ( .A(n26047), .B(n36766), .Y(n21792) );
  INVX1 U29024 ( .A(reg_file[3336]), .Y(n36766) );
  NOR2X1 U29025 ( .A(n26047), .B(n36767), .Y(n21791) );
  INVX1 U29026 ( .A(reg_file[3337]), .Y(n36767) );
  NOR2X1 U29027 ( .A(n26047), .B(n36768), .Y(n21790) );
  INVX1 U29028 ( .A(reg_file[3338]), .Y(n36768) );
  NOR2X1 U29029 ( .A(n26047), .B(n36769), .Y(n21789) );
  INVX1 U29030 ( .A(reg_file[3339]), .Y(n36769) );
  NOR2X1 U29031 ( .A(n26047), .B(n36770), .Y(n21788) );
  INVX1 U29032 ( .A(reg_file[3340]), .Y(n36770) );
  NOR2X1 U29033 ( .A(n26047), .B(n36771), .Y(n21787) );
  INVX1 U29034 ( .A(reg_file[3341]), .Y(n36771) );
  NOR2X1 U29035 ( .A(n26048), .B(n36772), .Y(n21786) );
  INVX1 U29036 ( .A(reg_file[3342]), .Y(n36772) );
  NOR2X1 U29037 ( .A(n26048), .B(n36773), .Y(n21785) );
  INVX1 U29038 ( .A(reg_file[3343]), .Y(n36773) );
  NOR2X1 U29039 ( .A(n26048), .B(n36774), .Y(n21784) );
  INVX1 U29040 ( .A(reg_file[3344]), .Y(n36774) );
  NOR2X1 U29041 ( .A(n26048), .B(n36775), .Y(n21783) );
  INVX1 U29042 ( .A(reg_file[3345]), .Y(n36775) );
  NOR2X1 U29043 ( .A(n26048), .B(n36776), .Y(n21782) );
  INVX1 U29044 ( .A(reg_file[3346]), .Y(n36776) );
  NOR2X1 U29045 ( .A(n26048), .B(n36777), .Y(n21781) );
  INVX1 U29046 ( .A(reg_file[3347]), .Y(n36777) );
  NOR2X1 U29047 ( .A(n26048), .B(n36778), .Y(n21780) );
  INVX1 U29048 ( .A(reg_file[3348]), .Y(n36778) );
  NOR2X1 U29049 ( .A(n26048), .B(n36779), .Y(n21779) );
  INVX1 U29050 ( .A(reg_file[3349]), .Y(n36779) );
  NOR2X1 U29051 ( .A(n26048), .B(n36780), .Y(n21778) );
  INVX1 U29052 ( .A(reg_file[3350]), .Y(n36780) );
  NOR2X1 U29053 ( .A(n26048), .B(n36781), .Y(n21777) );
  INVX1 U29054 ( .A(reg_file[3351]), .Y(n36781) );
  NOR2X1 U29055 ( .A(n26048), .B(n36782), .Y(n21776) );
  INVX1 U29056 ( .A(reg_file[3352]), .Y(n36782) );
  NOR2X1 U29057 ( .A(n26048), .B(n36783), .Y(n21775) );
  INVX1 U29058 ( .A(reg_file[3353]), .Y(n36783) );
  NOR2X1 U29059 ( .A(n26048), .B(n36784), .Y(n21774) );
  INVX1 U29060 ( .A(reg_file[3354]), .Y(n36784) );
  NOR2X1 U29061 ( .A(n26048), .B(n36785), .Y(n21773) );
  INVX1 U29062 ( .A(reg_file[3355]), .Y(n36785) );
  NOR2X1 U29063 ( .A(n26048), .B(n36786), .Y(n21772) );
  INVX1 U29064 ( .A(reg_file[3356]), .Y(n36786) );
  NOR2X1 U29065 ( .A(n26048), .B(n36787), .Y(n21771) );
  INVX1 U29066 ( .A(reg_file[3357]), .Y(n36787) );
  NOR2X1 U29067 ( .A(n26048), .B(n36788), .Y(n21770) );
  INVX1 U29068 ( .A(reg_file[3358]), .Y(n36788) );
  NOR2X1 U29069 ( .A(n26049), .B(n36789), .Y(n21769) );
  INVX1 U29070 ( .A(reg_file[3359]), .Y(n36789) );
  NOR2X1 U29071 ( .A(n26049), .B(n36790), .Y(n21768) );
  INVX1 U29072 ( .A(reg_file[3360]), .Y(n36790) );
  NOR2X1 U29073 ( .A(n26049), .B(n36791), .Y(n21767) );
  INVX1 U29074 ( .A(reg_file[3361]), .Y(n36791) );
  NOR2X1 U29075 ( .A(n26049), .B(n36792), .Y(n21766) );
  INVX1 U29076 ( .A(reg_file[3362]), .Y(n36792) );
  NOR2X1 U29077 ( .A(n26049), .B(n36793), .Y(n21765) );
  INVX1 U29078 ( .A(reg_file[3363]), .Y(n36793) );
  NOR2X1 U29079 ( .A(n26049), .B(n36794), .Y(n21764) );
  INVX1 U29080 ( .A(reg_file[3364]), .Y(n36794) );
  NOR2X1 U29081 ( .A(n26049), .B(n36795), .Y(n21763) );
  INVX1 U29082 ( .A(reg_file[3365]), .Y(n36795) );
  NOR2X1 U29083 ( .A(n26049), .B(n36796), .Y(n21762) );
  INVX1 U29084 ( .A(reg_file[3366]), .Y(n36796) );
  NOR2X1 U29085 ( .A(n26049), .B(n36797), .Y(n21761) );
  INVX1 U29086 ( .A(reg_file[3367]), .Y(n36797) );
  NOR2X1 U29087 ( .A(n26049), .B(n36798), .Y(n21760) );
  INVX1 U29088 ( .A(reg_file[3368]), .Y(n36798) );
  NOR2X1 U29089 ( .A(n26049), .B(n36799), .Y(n21759) );
  INVX1 U29090 ( .A(reg_file[3369]), .Y(n36799) );
  NOR2X1 U29091 ( .A(n26049), .B(n36800), .Y(n21758) );
  INVX1 U29092 ( .A(reg_file[3370]), .Y(n36800) );
  NOR2X1 U29093 ( .A(n26049), .B(n36801), .Y(n21757) );
  INVX1 U29094 ( .A(reg_file[3371]), .Y(n36801) );
  NOR2X1 U29095 ( .A(n26049), .B(n36802), .Y(n21756) );
  INVX1 U29096 ( .A(reg_file[3372]), .Y(n36802) );
  NOR2X1 U29097 ( .A(n26049), .B(n36803), .Y(n21755) );
  INVX1 U29098 ( .A(reg_file[3373]), .Y(n36803) );
  NOR2X1 U29099 ( .A(n26049), .B(n36804), .Y(n21754) );
  INVX1 U29100 ( .A(reg_file[3374]), .Y(n36804) );
  NOR2X1 U29101 ( .A(n26049), .B(n36805), .Y(n21753) );
  INVX1 U29102 ( .A(reg_file[3375]), .Y(n36805) );
  NOR2X1 U29103 ( .A(n26050), .B(n36806), .Y(n21752) );
  INVX1 U29104 ( .A(reg_file[3376]), .Y(n36806) );
  NOR2X1 U29105 ( .A(n26050), .B(n36807), .Y(n21751) );
  INVX1 U29106 ( .A(reg_file[3377]), .Y(n36807) );
  NOR2X1 U29107 ( .A(n26050), .B(n36808), .Y(n21750) );
  INVX1 U29108 ( .A(reg_file[3378]), .Y(n36808) );
  NOR2X1 U29109 ( .A(n26050), .B(n36809), .Y(n21749) );
  INVX1 U29110 ( .A(reg_file[3379]), .Y(n36809) );
  NOR2X1 U29111 ( .A(n26050), .B(n36810), .Y(n21748) );
  INVX1 U29112 ( .A(reg_file[3380]), .Y(n36810) );
  NOR2X1 U29113 ( .A(n26050), .B(n36811), .Y(n21747) );
  INVX1 U29114 ( .A(reg_file[3381]), .Y(n36811) );
  NOR2X1 U29115 ( .A(n26050), .B(n36812), .Y(n21746) );
  INVX1 U29116 ( .A(reg_file[3382]), .Y(n36812) );
  NOR2X1 U29117 ( .A(n26050), .B(n36813), .Y(n21745) );
  INVX1 U29118 ( .A(reg_file[3383]), .Y(n36813) );
  NOR2X1 U29119 ( .A(n26050), .B(n36814), .Y(n21744) );
  INVX1 U29120 ( .A(reg_file[3384]), .Y(n36814) );
  NOR2X1 U29121 ( .A(n26050), .B(n36815), .Y(n21743) );
  INVX1 U29122 ( .A(reg_file[3385]), .Y(n36815) );
  NOR2X1 U29123 ( .A(n26050), .B(n36816), .Y(n21742) );
  INVX1 U29124 ( .A(reg_file[3386]), .Y(n36816) );
  NOR2X1 U29125 ( .A(n26050), .B(n36817), .Y(n21741) );
  INVX1 U29126 ( .A(reg_file[3387]), .Y(n36817) );
  NOR2X1 U29127 ( .A(n26050), .B(n36818), .Y(n21740) );
  INVX1 U29128 ( .A(reg_file[3388]), .Y(n36818) );
  NOR2X1 U29129 ( .A(n26050), .B(n36819), .Y(n21739) );
  INVX1 U29130 ( .A(reg_file[3389]), .Y(n36819) );
  NOR2X1 U29131 ( .A(n26050), .B(n36820), .Y(n21738) );
  INVX1 U29132 ( .A(reg_file[3390]), .Y(n36820) );
  NOR2X1 U29133 ( .A(n26050), .B(n36821), .Y(n21737) );
  INVX1 U29134 ( .A(reg_file[3391]), .Y(n36821) );
  NOR2X1 U29135 ( .A(n26050), .B(n36822), .Y(n21736) );
  INVX1 U29136 ( .A(reg_file[3392]), .Y(n36822) );
  NOR2X1 U29137 ( .A(n26051), .B(n36823), .Y(n21735) );
  INVX1 U29138 ( .A(reg_file[3393]), .Y(n36823) );
  NOR2X1 U29139 ( .A(n26051), .B(n36824), .Y(n21734) );
  INVX1 U29140 ( .A(reg_file[3394]), .Y(n36824) );
  NOR2X1 U29141 ( .A(n26051), .B(n36825), .Y(n21733) );
  INVX1 U29142 ( .A(reg_file[3395]), .Y(n36825) );
  NOR2X1 U29143 ( .A(n26051), .B(n36826), .Y(n21732) );
  INVX1 U29144 ( .A(reg_file[3396]), .Y(n36826) );
  NOR2X1 U29145 ( .A(n26051), .B(n36827), .Y(n21731) );
  INVX1 U29146 ( .A(reg_file[3397]), .Y(n36827) );
  NOR2X1 U29147 ( .A(n26051), .B(n36828), .Y(n21730) );
  INVX1 U29148 ( .A(reg_file[3398]), .Y(n36828) );
  NOR2X1 U29149 ( .A(n26051), .B(n36829), .Y(n21729) );
  INVX1 U29150 ( .A(reg_file[3399]), .Y(n36829) );
  NOR2X1 U29151 ( .A(n26051), .B(n36830), .Y(n21728) );
  INVX1 U29152 ( .A(reg_file[3400]), .Y(n36830) );
  NOR2X1 U29153 ( .A(n26051), .B(n36831), .Y(n21727) );
  INVX1 U29154 ( .A(reg_file[3401]), .Y(n36831) );
  NOR2X1 U29155 ( .A(n26051), .B(n36832), .Y(n21726) );
  INVX1 U29156 ( .A(reg_file[3402]), .Y(n36832) );
  NOR2X1 U29157 ( .A(n26051), .B(n36833), .Y(n21725) );
  INVX1 U29158 ( .A(reg_file[3403]), .Y(n36833) );
  NOR2X1 U29159 ( .A(n26051), .B(n36834), .Y(n21724) );
  INVX1 U29160 ( .A(reg_file[3404]), .Y(n36834) );
  NOR2X1 U29161 ( .A(n26051), .B(n36835), .Y(n21723) );
  INVX1 U29162 ( .A(reg_file[3405]), .Y(n36835) );
  NOR2X1 U29163 ( .A(n26051), .B(n36836), .Y(n21722) );
  INVX1 U29164 ( .A(reg_file[3406]), .Y(n36836) );
  NOR2X1 U29165 ( .A(n26051), .B(n36837), .Y(n21721) );
  INVX1 U29166 ( .A(reg_file[3407]), .Y(n36837) );
  NOR2X1 U29167 ( .A(n26051), .B(n36838), .Y(n21720) );
  INVX1 U29168 ( .A(reg_file[3408]), .Y(n36838) );
  NOR2X1 U29169 ( .A(n26051), .B(n36839), .Y(n21719) );
  INVX1 U29170 ( .A(reg_file[3409]), .Y(n36839) );
  NOR2X1 U29171 ( .A(n26052), .B(n36840), .Y(n21718) );
  INVX1 U29172 ( .A(reg_file[3410]), .Y(n36840) );
  NOR2X1 U29173 ( .A(n26052), .B(n36841), .Y(n21717) );
  INVX1 U29174 ( .A(reg_file[3411]), .Y(n36841) );
  NOR2X1 U29175 ( .A(n26052), .B(n36842), .Y(n21716) );
  INVX1 U29176 ( .A(reg_file[3412]), .Y(n36842) );
  NOR2X1 U29177 ( .A(n26052), .B(n36843), .Y(n21715) );
  INVX1 U29178 ( .A(reg_file[3413]), .Y(n36843) );
  NOR2X1 U29179 ( .A(n26052), .B(n36844), .Y(n21714) );
  INVX1 U29180 ( .A(reg_file[3414]), .Y(n36844) );
  NOR2X1 U29181 ( .A(n26052), .B(n36845), .Y(n21713) );
  INVX1 U29182 ( .A(reg_file[3415]), .Y(n36845) );
  NOR2X1 U29183 ( .A(n26052), .B(n36846), .Y(n21712) );
  INVX1 U29184 ( .A(reg_file[3416]), .Y(n36846) );
  NOR2X1 U29185 ( .A(n26052), .B(n36847), .Y(n21711) );
  INVX1 U29186 ( .A(reg_file[3417]), .Y(n36847) );
  NOR2X1 U29187 ( .A(n26052), .B(n36848), .Y(n21710) );
  INVX1 U29188 ( .A(reg_file[3418]), .Y(n36848) );
  NOR2X1 U29189 ( .A(n26052), .B(n36849), .Y(n21709) );
  INVX1 U29190 ( .A(reg_file[3419]), .Y(n36849) );
  NOR2X1 U29191 ( .A(n26052), .B(n36850), .Y(n21708) );
  INVX1 U29192 ( .A(reg_file[3420]), .Y(n36850) );
  NOR2X1 U29193 ( .A(n26052), .B(n36851), .Y(n21707) );
  INVX1 U29194 ( .A(reg_file[3421]), .Y(n36851) );
  NOR2X1 U29195 ( .A(n26052), .B(n36852), .Y(n21706) );
  INVX1 U29196 ( .A(reg_file[3422]), .Y(n36852) );
  NOR2X1 U29197 ( .A(n26052), .B(n36853), .Y(n21705) );
  INVX1 U29198 ( .A(reg_file[3423]), .Y(n36853) );
  NOR2X1 U29199 ( .A(n26052), .B(n36854), .Y(n21704) );
  INVX1 U29200 ( .A(reg_file[3424]), .Y(n36854) );
  NOR2X1 U29201 ( .A(n26052), .B(n36855), .Y(n21703) );
  INVX1 U29202 ( .A(reg_file[3425]), .Y(n36855) );
  NOR2X1 U29203 ( .A(n26052), .B(n36856), .Y(n21702) );
  INVX1 U29204 ( .A(reg_file[3426]), .Y(n36856) );
  NOR2X1 U29205 ( .A(n26053), .B(n36857), .Y(n21701) );
  INVX1 U29206 ( .A(reg_file[3427]), .Y(n36857) );
  NOR2X1 U29207 ( .A(n26053), .B(n36858), .Y(n21700) );
  INVX1 U29208 ( .A(reg_file[3428]), .Y(n36858) );
  NOR2X1 U29209 ( .A(n26053), .B(n36859), .Y(n21699) );
  INVX1 U29210 ( .A(reg_file[3429]), .Y(n36859) );
  NOR2X1 U29211 ( .A(n26053), .B(n36860), .Y(n21698) );
  INVX1 U29212 ( .A(reg_file[3430]), .Y(n36860) );
  NOR2X1 U29213 ( .A(n26053), .B(n36861), .Y(n21697) );
  INVX1 U29214 ( .A(reg_file[3431]), .Y(n36861) );
  NOR2X1 U29215 ( .A(n26053), .B(n36862), .Y(n21696) );
  INVX1 U29216 ( .A(reg_file[3432]), .Y(n36862) );
  NOR2X1 U29217 ( .A(n26053), .B(n36863), .Y(n21695) );
  INVX1 U29218 ( .A(reg_file[3433]), .Y(n36863) );
  NOR2X1 U29219 ( .A(n26053), .B(n36864), .Y(n21694) );
  INVX1 U29220 ( .A(reg_file[3434]), .Y(n36864) );
  NOR2X1 U29221 ( .A(n26053), .B(n36865), .Y(n21693) );
  INVX1 U29222 ( .A(reg_file[3435]), .Y(n36865) );
  NOR2X1 U29223 ( .A(n26053), .B(n36866), .Y(n21692) );
  INVX1 U29224 ( .A(reg_file[3436]), .Y(n36866) );
  NOR2X1 U29225 ( .A(n26053), .B(n36867), .Y(n21691) );
  INVX1 U29226 ( .A(reg_file[3437]), .Y(n36867) );
  NOR2X1 U29227 ( .A(n26053), .B(n36868), .Y(n21690) );
  INVX1 U29228 ( .A(reg_file[3438]), .Y(n36868) );
  NOR2X1 U29229 ( .A(n26053), .B(n36869), .Y(n21689) );
  INVX1 U29230 ( .A(reg_file[3439]), .Y(n36869) );
  NOR2X1 U29231 ( .A(n26053), .B(n36870), .Y(n21688) );
  INVX1 U29232 ( .A(reg_file[3440]), .Y(n36870) );
  NOR2X1 U29233 ( .A(n26053), .B(n36871), .Y(n21687) );
  INVX1 U29234 ( .A(reg_file[3441]), .Y(n36871) );
  NOR2X1 U29235 ( .A(n26053), .B(n36872), .Y(n21686) );
  INVX1 U29236 ( .A(reg_file[3442]), .Y(n36872) );
  NOR2X1 U29237 ( .A(n26053), .B(n36873), .Y(n21685) );
  INVX1 U29238 ( .A(reg_file[3443]), .Y(n36873) );
  NOR2X1 U29239 ( .A(n26054), .B(n36874), .Y(n21684) );
  INVX1 U29240 ( .A(reg_file[3444]), .Y(n36874) );
  NOR2X1 U29241 ( .A(n26054), .B(n36875), .Y(n21683) );
  INVX1 U29242 ( .A(reg_file[3445]), .Y(n36875) );
  NOR2X1 U29243 ( .A(n26054), .B(n36876), .Y(n21682) );
  INVX1 U29244 ( .A(reg_file[3446]), .Y(n36876) );
  NOR2X1 U29245 ( .A(n26054), .B(n36877), .Y(n21681) );
  INVX1 U29246 ( .A(reg_file[3447]), .Y(n36877) );
  NOR2X1 U29247 ( .A(n26054), .B(n36878), .Y(n21680) );
  INVX1 U29248 ( .A(reg_file[3448]), .Y(n36878) );
  NOR2X1 U29249 ( .A(n26054), .B(n36879), .Y(n21679) );
  INVX1 U29250 ( .A(reg_file[3449]), .Y(n36879) );
  NOR2X1 U29251 ( .A(n26054), .B(n36880), .Y(n21678) );
  INVX1 U29252 ( .A(reg_file[3450]), .Y(n36880) );
  NOR2X1 U29253 ( .A(n26054), .B(n36881), .Y(n21677) );
  INVX1 U29254 ( .A(reg_file[3451]), .Y(n36881) );
  NOR2X1 U29255 ( .A(n26054), .B(n36882), .Y(n21676) );
  INVX1 U29256 ( .A(reg_file[3452]), .Y(n36882) );
  NOR2X1 U29257 ( .A(n26054), .B(n36883), .Y(n21675) );
  INVX1 U29258 ( .A(reg_file[3453]), .Y(n36883) );
  NOR2X1 U29259 ( .A(n26054), .B(n36884), .Y(n21674) );
  INVX1 U29260 ( .A(reg_file[3454]), .Y(n36884) );
  NOR2X1 U29261 ( .A(n26054), .B(n36885), .Y(n21673) );
  INVX1 U29262 ( .A(reg_file[3455]), .Y(n36885) );
  NOR2X1 U29263 ( .A(n36623), .B(n34927), .Y(n36758) );
  MUX2X1 U29264 ( .B(n36886), .A(n25129), .S(n26055), .Y(n21672) );
  INVX1 U29265 ( .A(reg_file[3456]), .Y(n36886) );
  MUX2X1 U29266 ( .B(n36888), .A(n25130), .S(n26055), .Y(n21671) );
  INVX1 U29267 ( .A(reg_file[3457]), .Y(n36888) );
  MUX2X1 U29268 ( .B(n36889), .A(n25131), .S(n26055), .Y(n21670) );
  INVX1 U29269 ( .A(reg_file[3458]), .Y(n36889) );
  MUX2X1 U29270 ( .B(n36890), .A(n25132), .S(n26055), .Y(n21669) );
  INVX1 U29271 ( .A(reg_file[3459]), .Y(n36890) );
  MUX2X1 U29272 ( .B(n36891), .A(n25133), .S(n26055), .Y(n21668) );
  INVX1 U29273 ( .A(reg_file[3460]), .Y(n36891) );
  MUX2X1 U29274 ( .B(n36892), .A(n25134), .S(n26055), .Y(n21667) );
  INVX1 U29275 ( .A(reg_file[3461]), .Y(n36892) );
  MUX2X1 U29276 ( .B(n36893), .A(n25135), .S(n26055), .Y(n21666) );
  INVX1 U29277 ( .A(reg_file[3462]), .Y(n36893) );
  MUX2X1 U29278 ( .B(n36894), .A(n25136), .S(n26055), .Y(n21665) );
  INVX1 U29279 ( .A(reg_file[3463]), .Y(n36894) );
  NOR2X1 U29280 ( .A(n26055), .B(n36895), .Y(n21664) );
  INVX1 U29281 ( .A(reg_file[3464]), .Y(n36895) );
  NOR2X1 U29282 ( .A(n26055), .B(n36896), .Y(n21663) );
  INVX1 U29283 ( .A(reg_file[3465]), .Y(n36896) );
  NOR2X1 U29284 ( .A(n26055), .B(n36897), .Y(n21662) );
  INVX1 U29285 ( .A(reg_file[3466]), .Y(n36897) );
  NOR2X1 U29286 ( .A(n26055), .B(n36898), .Y(n21661) );
  INVX1 U29287 ( .A(reg_file[3467]), .Y(n36898) );
  NOR2X1 U29288 ( .A(n26055), .B(n36899), .Y(n21660) );
  INVX1 U29289 ( .A(reg_file[3468]), .Y(n36899) );
  NOR2X1 U29290 ( .A(n26055), .B(n36900), .Y(n21659) );
  INVX1 U29291 ( .A(reg_file[3469]), .Y(n36900) );
  NOR2X1 U29292 ( .A(n26056), .B(n36901), .Y(n21658) );
  INVX1 U29293 ( .A(reg_file[3470]), .Y(n36901) );
  NOR2X1 U29294 ( .A(n26056), .B(n36902), .Y(n21657) );
  INVX1 U29295 ( .A(reg_file[3471]), .Y(n36902) );
  NOR2X1 U29296 ( .A(n26056), .B(n36903), .Y(n21656) );
  INVX1 U29297 ( .A(reg_file[3472]), .Y(n36903) );
  NOR2X1 U29298 ( .A(n26056), .B(n36904), .Y(n21655) );
  INVX1 U29299 ( .A(reg_file[3473]), .Y(n36904) );
  NOR2X1 U29300 ( .A(n26056), .B(n36905), .Y(n21654) );
  INVX1 U29301 ( .A(reg_file[3474]), .Y(n36905) );
  NOR2X1 U29302 ( .A(n26056), .B(n36906), .Y(n21653) );
  INVX1 U29303 ( .A(reg_file[3475]), .Y(n36906) );
  NOR2X1 U29304 ( .A(n26056), .B(n36907), .Y(n21652) );
  INVX1 U29305 ( .A(reg_file[3476]), .Y(n36907) );
  NOR2X1 U29306 ( .A(n26056), .B(n36908), .Y(n21651) );
  INVX1 U29307 ( .A(reg_file[3477]), .Y(n36908) );
  NOR2X1 U29308 ( .A(n26056), .B(n36909), .Y(n21650) );
  INVX1 U29309 ( .A(reg_file[3478]), .Y(n36909) );
  NOR2X1 U29310 ( .A(n26056), .B(n36910), .Y(n21649) );
  INVX1 U29311 ( .A(reg_file[3479]), .Y(n36910) );
  NOR2X1 U29312 ( .A(n26056), .B(n36911), .Y(n21648) );
  INVX1 U29313 ( .A(reg_file[3480]), .Y(n36911) );
  NOR2X1 U29314 ( .A(n26056), .B(n36912), .Y(n21647) );
  INVX1 U29315 ( .A(reg_file[3481]), .Y(n36912) );
  NOR2X1 U29316 ( .A(n26056), .B(n36913), .Y(n21646) );
  INVX1 U29317 ( .A(reg_file[3482]), .Y(n36913) );
  NOR2X1 U29318 ( .A(n26056), .B(n36914), .Y(n21645) );
  INVX1 U29319 ( .A(reg_file[3483]), .Y(n36914) );
  NOR2X1 U29320 ( .A(n26056), .B(n36915), .Y(n21644) );
  INVX1 U29321 ( .A(reg_file[3484]), .Y(n36915) );
  NOR2X1 U29322 ( .A(n26056), .B(n36916), .Y(n21643) );
  INVX1 U29323 ( .A(reg_file[3485]), .Y(n36916) );
  NOR2X1 U29324 ( .A(n26056), .B(n36917), .Y(n21642) );
  INVX1 U29325 ( .A(reg_file[3486]), .Y(n36917) );
  NOR2X1 U29326 ( .A(n26057), .B(n36918), .Y(n21641) );
  INVX1 U29327 ( .A(reg_file[3487]), .Y(n36918) );
  NOR2X1 U29328 ( .A(n26057), .B(n36919), .Y(n21640) );
  INVX1 U29329 ( .A(reg_file[3488]), .Y(n36919) );
  NOR2X1 U29330 ( .A(n26057), .B(n36920), .Y(n21639) );
  INVX1 U29331 ( .A(reg_file[3489]), .Y(n36920) );
  NOR2X1 U29332 ( .A(n26057), .B(n36921), .Y(n21638) );
  INVX1 U29333 ( .A(reg_file[3490]), .Y(n36921) );
  NOR2X1 U29334 ( .A(n26057), .B(n36922), .Y(n21637) );
  INVX1 U29335 ( .A(reg_file[3491]), .Y(n36922) );
  NOR2X1 U29336 ( .A(n26057), .B(n36923), .Y(n21636) );
  INVX1 U29337 ( .A(reg_file[3492]), .Y(n36923) );
  NOR2X1 U29338 ( .A(n26057), .B(n36924), .Y(n21635) );
  INVX1 U29339 ( .A(reg_file[3493]), .Y(n36924) );
  NOR2X1 U29340 ( .A(n26057), .B(n36925), .Y(n21634) );
  INVX1 U29341 ( .A(reg_file[3494]), .Y(n36925) );
  NOR2X1 U29342 ( .A(n26057), .B(n36926), .Y(n21633) );
  INVX1 U29343 ( .A(reg_file[3495]), .Y(n36926) );
  NOR2X1 U29344 ( .A(n26057), .B(n36927), .Y(n21632) );
  INVX1 U29345 ( .A(reg_file[3496]), .Y(n36927) );
  NOR2X1 U29346 ( .A(n26057), .B(n36928), .Y(n21631) );
  INVX1 U29347 ( .A(reg_file[3497]), .Y(n36928) );
  NOR2X1 U29348 ( .A(n26057), .B(n36929), .Y(n21630) );
  INVX1 U29349 ( .A(reg_file[3498]), .Y(n36929) );
  NOR2X1 U29350 ( .A(n26057), .B(n36930), .Y(n21629) );
  INVX1 U29351 ( .A(reg_file[3499]), .Y(n36930) );
  NOR2X1 U29352 ( .A(n26057), .B(n36931), .Y(n21628) );
  INVX1 U29353 ( .A(reg_file[3500]), .Y(n36931) );
  NOR2X1 U29354 ( .A(n26057), .B(n36932), .Y(n21627) );
  INVX1 U29355 ( .A(reg_file[3501]), .Y(n36932) );
  NOR2X1 U29356 ( .A(n26057), .B(n36933), .Y(n21626) );
  INVX1 U29357 ( .A(reg_file[3502]), .Y(n36933) );
  NOR2X1 U29358 ( .A(n26057), .B(n36934), .Y(n21625) );
  INVX1 U29359 ( .A(reg_file[3503]), .Y(n36934) );
  NOR2X1 U29360 ( .A(n26058), .B(n36935), .Y(n21624) );
  INVX1 U29361 ( .A(reg_file[3504]), .Y(n36935) );
  NOR2X1 U29362 ( .A(n26058), .B(n36936), .Y(n21623) );
  INVX1 U29363 ( .A(reg_file[3505]), .Y(n36936) );
  NOR2X1 U29364 ( .A(n26058), .B(n36937), .Y(n21622) );
  INVX1 U29365 ( .A(reg_file[3506]), .Y(n36937) );
  NOR2X1 U29366 ( .A(n26058), .B(n36938), .Y(n21621) );
  INVX1 U29367 ( .A(reg_file[3507]), .Y(n36938) );
  NOR2X1 U29368 ( .A(n26058), .B(n36939), .Y(n21620) );
  INVX1 U29369 ( .A(reg_file[3508]), .Y(n36939) );
  NOR2X1 U29370 ( .A(n26058), .B(n36940), .Y(n21619) );
  INVX1 U29371 ( .A(reg_file[3509]), .Y(n36940) );
  NOR2X1 U29372 ( .A(n26058), .B(n36941), .Y(n21618) );
  INVX1 U29373 ( .A(reg_file[3510]), .Y(n36941) );
  NOR2X1 U29374 ( .A(n26058), .B(n36942), .Y(n21617) );
  INVX1 U29375 ( .A(reg_file[3511]), .Y(n36942) );
  NOR2X1 U29376 ( .A(n26058), .B(n36943), .Y(n21616) );
  INVX1 U29377 ( .A(reg_file[3512]), .Y(n36943) );
  NOR2X1 U29378 ( .A(n26058), .B(n36944), .Y(n21615) );
  INVX1 U29379 ( .A(reg_file[3513]), .Y(n36944) );
  NOR2X1 U29380 ( .A(n26058), .B(n36945), .Y(n21614) );
  INVX1 U29381 ( .A(reg_file[3514]), .Y(n36945) );
  NOR2X1 U29382 ( .A(n26058), .B(n36946), .Y(n21613) );
  INVX1 U29383 ( .A(reg_file[3515]), .Y(n36946) );
  NOR2X1 U29384 ( .A(n26058), .B(n36947), .Y(n21612) );
  INVX1 U29385 ( .A(reg_file[3516]), .Y(n36947) );
  NOR2X1 U29386 ( .A(n26058), .B(n36948), .Y(n21611) );
  INVX1 U29387 ( .A(reg_file[3517]), .Y(n36948) );
  NOR2X1 U29388 ( .A(n26058), .B(n36949), .Y(n21610) );
  INVX1 U29389 ( .A(reg_file[3518]), .Y(n36949) );
  NOR2X1 U29390 ( .A(n26058), .B(n36950), .Y(n21609) );
  INVX1 U29391 ( .A(reg_file[3519]), .Y(n36950) );
  NOR2X1 U29392 ( .A(n26058), .B(n36951), .Y(n21608) );
  INVX1 U29393 ( .A(reg_file[3520]), .Y(n36951) );
  NOR2X1 U29394 ( .A(n26059), .B(n36952), .Y(n21607) );
  INVX1 U29395 ( .A(reg_file[3521]), .Y(n36952) );
  NOR2X1 U29396 ( .A(n26059), .B(n36953), .Y(n21606) );
  INVX1 U29397 ( .A(reg_file[3522]), .Y(n36953) );
  NOR2X1 U29398 ( .A(n26059), .B(n36954), .Y(n21605) );
  INVX1 U29399 ( .A(reg_file[3523]), .Y(n36954) );
  NOR2X1 U29400 ( .A(n26059), .B(n36955), .Y(n21604) );
  INVX1 U29401 ( .A(reg_file[3524]), .Y(n36955) );
  NOR2X1 U29402 ( .A(n26059), .B(n36956), .Y(n21603) );
  INVX1 U29403 ( .A(reg_file[3525]), .Y(n36956) );
  NOR2X1 U29404 ( .A(n26059), .B(n36957), .Y(n21602) );
  INVX1 U29405 ( .A(reg_file[3526]), .Y(n36957) );
  NOR2X1 U29406 ( .A(n26059), .B(n36958), .Y(n21601) );
  INVX1 U29407 ( .A(reg_file[3527]), .Y(n36958) );
  NOR2X1 U29408 ( .A(n26059), .B(n36959), .Y(n21600) );
  INVX1 U29409 ( .A(reg_file[3528]), .Y(n36959) );
  NOR2X1 U29410 ( .A(n26059), .B(n36960), .Y(n21599) );
  INVX1 U29411 ( .A(reg_file[3529]), .Y(n36960) );
  NOR2X1 U29412 ( .A(n26059), .B(n36961), .Y(n21598) );
  INVX1 U29413 ( .A(reg_file[3530]), .Y(n36961) );
  NOR2X1 U29414 ( .A(n26059), .B(n36962), .Y(n21597) );
  INVX1 U29415 ( .A(reg_file[3531]), .Y(n36962) );
  NOR2X1 U29416 ( .A(n26059), .B(n36963), .Y(n21596) );
  INVX1 U29417 ( .A(reg_file[3532]), .Y(n36963) );
  NOR2X1 U29418 ( .A(n26059), .B(n36964), .Y(n21595) );
  INVX1 U29419 ( .A(reg_file[3533]), .Y(n36964) );
  NOR2X1 U29420 ( .A(n26059), .B(n36965), .Y(n21594) );
  INVX1 U29421 ( .A(reg_file[3534]), .Y(n36965) );
  NOR2X1 U29422 ( .A(n26059), .B(n36966), .Y(n21593) );
  INVX1 U29423 ( .A(reg_file[3535]), .Y(n36966) );
  NOR2X1 U29424 ( .A(n26059), .B(n36967), .Y(n21592) );
  INVX1 U29425 ( .A(reg_file[3536]), .Y(n36967) );
  NOR2X1 U29426 ( .A(n26059), .B(n36968), .Y(n21591) );
  INVX1 U29427 ( .A(reg_file[3537]), .Y(n36968) );
  NOR2X1 U29428 ( .A(n26060), .B(n36969), .Y(n21590) );
  INVX1 U29429 ( .A(reg_file[3538]), .Y(n36969) );
  NOR2X1 U29430 ( .A(n26060), .B(n36970), .Y(n21589) );
  INVX1 U29431 ( .A(reg_file[3539]), .Y(n36970) );
  NOR2X1 U29432 ( .A(n26060), .B(n36971), .Y(n21588) );
  INVX1 U29433 ( .A(reg_file[3540]), .Y(n36971) );
  NOR2X1 U29434 ( .A(n26060), .B(n36972), .Y(n21587) );
  INVX1 U29435 ( .A(reg_file[3541]), .Y(n36972) );
  NOR2X1 U29436 ( .A(n26060), .B(n36973), .Y(n21586) );
  INVX1 U29437 ( .A(reg_file[3542]), .Y(n36973) );
  NOR2X1 U29438 ( .A(n26060), .B(n36974), .Y(n21585) );
  INVX1 U29439 ( .A(reg_file[3543]), .Y(n36974) );
  NOR2X1 U29440 ( .A(n26060), .B(n36975), .Y(n21584) );
  INVX1 U29441 ( .A(reg_file[3544]), .Y(n36975) );
  NOR2X1 U29442 ( .A(n26060), .B(n36976), .Y(n21583) );
  INVX1 U29443 ( .A(reg_file[3545]), .Y(n36976) );
  NOR2X1 U29444 ( .A(n26060), .B(n36977), .Y(n21582) );
  INVX1 U29445 ( .A(reg_file[3546]), .Y(n36977) );
  NOR2X1 U29446 ( .A(n26060), .B(n36978), .Y(n21581) );
  INVX1 U29447 ( .A(reg_file[3547]), .Y(n36978) );
  NOR2X1 U29448 ( .A(n26060), .B(n36979), .Y(n21580) );
  INVX1 U29449 ( .A(reg_file[3548]), .Y(n36979) );
  NOR2X1 U29450 ( .A(n26060), .B(n36980), .Y(n21579) );
  INVX1 U29451 ( .A(reg_file[3549]), .Y(n36980) );
  NOR2X1 U29452 ( .A(n26060), .B(n36981), .Y(n21578) );
  INVX1 U29453 ( .A(reg_file[3550]), .Y(n36981) );
  NOR2X1 U29454 ( .A(n26060), .B(n36982), .Y(n21577) );
  INVX1 U29455 ( .A(reg_file[3551]), .Y(n36982) );
  NOR2X1 U29456 ( .A(n26060), .B(n36983), .Y(n21576) );
  INVX1 U29457 ( .A(reg_file[3552]), .Y(n36983) );
  NOR2X1 U29458 ( .A(n26060), .B(n36984), .Y(n21575) );
  INVX1 U29459 ( .A(reg_file[3553]), .Y(n36984) );
  NOR2X1 U29460 ( .A(n26060), .B(n36985), .Y(n21574) );
  INVX1 U29461 ( .A(reg_file[3554]), .Y(n36985) );
  NOR2X1 U29462 ( .A(n26061), .B(n36986), .Y(n21573) );
  INVX1 U29463 ( .A(reg_file[3555]), .Y(n36986) );
  NOR2X1 U29464 ( .A(n26061), .B(n36987), .Y(n21572) );
  INVX1 U29465 ( .A(reg_file[3556]), .Y(n36987) );
  NOR2X1 U29466 ( .A(n26061), .B(n36988), .Y(n21571) );
  INVX1 U29467 ( .A(reg_file[3557]), .Y(n36988) );
  NOR2X1 U29468 ( .A(n26061), .B(n36989), .Y(n21570) );
  INVX1 U29469 ( .A(reg_file[3558]), .Y(n36989) );
  NOR2X1 U29470 ( .A(n26061), .B(n36990), .Y(n21569) );
  INVX1 U29471 ( .A(reg_file[3559]), .Y(n36990) );
  NOR2X1 U29472 ( .A(n26061), .B(n36991), .Y(n21568) );
  INVX1 U29473 ( .A(reg_file[3560]), .Y(n36991) );
  NOR2X1 U29474 ( .A(n26061), .B(n36992), .Y(n21567) );
  INVX1 U29475 ( .A(reg_file[3561]), .Y(n36992) );
  NOR2X1 U29476 ( .A(n26061), .B(n36993), .Y(n21566) );
  INVX1 U29477 ( .A(reg_file[3562]), .Y(n36993) );
  NOR2X1 U29478 ( .A(n26061), .B(n36994), .Y(n21565) );
  INVX1 U29479 ( .A(reg_file[3563]), .Y(n36994) );
  NOR2X1 U29480 ( .A(n26061), .B(n36995), .Y(n21564) );
  INVX1 U29481 ( .A(reg_file[3564]), .Y(n36995) );
  NOR2X1 U29482 ( .A(n26061), .B(n36996), .Y(n21563) );
  INVX1 U29483 ( .A(reg_file[3565]), .Y(n36996) );
  NOR2X1 U29484 ( .A(n26061), .B(n36997), .Y(n21562) );
  INVX1 U29485 ( .A(reg_file[3566]), .Y(n36997) );
  NOR2X1 U29486 ( .A(n26061), .B(n36998), .Y(n21561) );
  INVX1 U29487 ( .A(reg_file[3567]), .Y(n36998) );
  NOR2X1 U29488 ( .A(n26061), .B(n36999), .Y(n21560) );
  INVX1 U29489 ( .A(reg_file[3568]), .Y(n36999) );
  NOR2X1 U29490 ( .A(n26061), .B(n37000), .Y(n21559) );
  INVX1 U29491 ( .A(reg_file[3569]), .Y(n37000) );
  NOR2X1 U29492 ( .A(n26061), .B(n37001), .Y(n21558) );
  INVX1 U29493 ( .A(reg_file[3570]), .Y(n37001) );
  NOR2X1 U29494 ( .A(n26061), .B(n37002), .Y(n21557) );
  INVX1 U29495 ( .A(reg_file[3571]), .Y(n37002) );
  NOR2X1 U29496 ( .A(n26062), .B(n37003), .Y(n21556) );
  INVX1 U29497 ( .A(reg_file[3572]), .Y(n37003) );
  NOR2X1 U29498 ( .A(n26062), .B(n37004), .Y(n21555) );
  INVX1 U29499 ( .A(reg_file[3573]), .Y(n37004) );
  NOR2X1 U29500 ( .A(n26062), .B(n37005), .Y(n21554) );
  INVX1 U29501 ( .A(reg_file[3574]), .Y(n37005) );
  NOR2X1 U29502 ( .A(n26062), .B(n37006), .Y(n21553) );
  INVX1 U29503 ( .A(reg_file[3575]), .Y(n37006) );
  NOR2X1 U29504 ( .A(n26062), .B(n37007), .Y(n21552) );
  INVX1 U29505 ( .A(reg_file[3576]), .Y(n37007) );
  NOR2X1 U29506 ( .A(n26062), .B(n37008), .Y(n21551) );
  INVX1 U29507 ( .A(reg_file[3577]), .Y(n37008) );
  NOR2X1 U29508 ( .A(n26062), .B(n37009), .Y(n21550) );
  INVX1 U29509 ( .A(reg_file[3578]), .Y(n37009) );
  NOR2X1 U29510 ( .A(n26062), .B(n37010), .Y(n21549) );
  INVX1 U29511 ( .A(reg_file[3579]), .Y(n37010) );
  NOR2X1 U29512 ( .A(n26062), .B(n37011), .Y(n21548) );
  INVX1 U29513 ( .A(reg_file[3580]), .Y(n37011) );
  NOR2X1 U29514 ( .A(n26062), .B(n37012), .Y(n21547) );
  INVX1 U29515 ( .A(reg_file[3581]), .Y(n37012) );
  NOR2X1 U29516 ( .A(n26062), .B(n37013), .Y(n21546) );
  INVX1 U29517 ( .A(reg_file[3582]), .Y(n37013) );
  NOR2X1 U29518 ( .A(n26062), .B(n37014), .Y(n21545) );
  INVX1 U29519 ( .A(reg_file[3583]), .Y(n37014) );
  NOR2X1 U29520 ( .A(n36753), .B(n34927), .Y(n36887) );
  NAND3X1 U29521 ( .A(n36756), .B(n36755), .C(wraddr[1]), .Y(n34927) );
  INVX1 U29522 ( .A(wraddr[2]), .Y(n36755) );
  MUX2X1 U29523 ( .B(n31506), .A(n25129), .S(n26063), .Y(n21544) );
  INVX1 U29524 ( .A(reg_file[3584]), .Y(n31506) );
  MUX2X1 U29525 ( .B(n29853), .A(n25130), .S(n26063), .Y(n21543) );
  INVX1 U29526 ( .A(reg_file[3585]), .Y(n29853) );
  MUX2X1 U29527 ( .B(n29391), .A(n25131), .S(n26063), .Y(n21542) );
  INVX1 U29528 ( .A(reg_file[3586]), .Y(n29391) );
  MUX2X1 U29529 ( .B(n28929), .A(n25132), .S(n26063), .Y(n21541) );
  INVX1 U29530 ( .A(reg_file[3587]), .Y(n28929) );
  MUX2X1 U29531 ( .B(n28467), .A(n25133), .S(n26063), .Y(n21540) );
  INVX1 U29532 ( .A(reg_file[3588]), .Y(n28467) );
  MUX2X1 U29533 ( .B(n28005), .A(n25134), .S(n26063), .Y(n21539) );
  INVX1 U29534 ( .A(reg_file[3589]), .Y(n28005) );
  MUX2X1 U29535 ( .B(n27543), .A(n25135), .S(n26063), .Y(n21538) );
  INVX1 U29536 ( .A(reg_file[3590]), .Y(n27543) );
  MUX2X1 U29537 ( .B(n27081), .A(n25136), .S(n26063), .Y(n21537) );
  INVX1 U29538 ( .A(reg_file[3591]), .Y(n27081) );
  NOR2X1 U29539 ( .A(n26063), .B(n26619), .Y(n21536) );
  INVX1 U29540 ( .A(reg_file[3592]), .Y(n26619) );
  NOR2X1 U29541 ( .A(n26063), .B(n26142), .Y(n21535) );
  INVX1 U29542 ( .A(reg_file[3593]), .Y(n26142) );
  NOR2X1 U29543 ( .A(n26063), .B(n31029), .Y(n21534) );
  INVX1 U29544 ( .A(reg_file[3594]), .Y(n31029) );
  NOR2X1 U29545 ( .A(n26063), .B(n30567), .Y(n21533) );
  INVX1 U29546 ( .A(reg_file[3595]), .Y(n30567) );
  NOR2X1 U29547 ( .A(n26063), .B(n30189), .Y(n21532) );
  INVX1 U29548 ( .A(reg_file[3596]), .Y(n30189) );
  NOR2X1 U29549 ( .A(n26063), .B(n30147), .Y(n21531) );
  INVX1 U29550 ( .A(reg_file[3597]), .Y(n30147) );
  NOR2X1 U29551 ( .A(n26064), .B(n30105), .Y(n21530) );
  INVX1 U29552 ( .A(reg_file[3598]), .Y(n30105) );
  NOR2X1 U29553 ( .A(n26064), .B(n30063), .Y(n21529) );
  INVX1 U29554 ( .A(reg_file[3599]), .Y(n30063) );
  NOR2X1 U29555 ( .A(n26064), .B(n30021), .Y(n21528) );
  INVX1 U29556 ( .A(reg_file[3600]), .Y(n30021) );
  NOR2X1 U29557 ( .A(n26064), .B(n29979), .Y(n21527) );
  INVX1 U29558 ( .A(reg_file[3601]), .Y(n29979) );
  NOR2X1 U29559 ( .A(n26064), .B(n29937), .Y(n21526) );
  INVX1 U29560 ( .A(reg_file[3602]), .Y(n29937) );
  NOR2X1 U29561 ( .A(n26064), .B(n29895), .Y(n21525) );
  INVX1 U29562 ( .A(reg_file[3603]), .Y(n29895) );
  NOR2X1 U29563 ( .A(n26064), .B(n29811), .Y(n21524) );
  INVX1 U29564 ( .A(reg_file[3604]), .Y(n29811) );
  NOR2X1 U29565 ( .A(n26064), .B(n29769), .Y(n21523) );
  INVX1 U29566 ( .A(reg_file[3605]), .Y(n29769) );
  NOR2X1 U29567 ( .A(n26064), .B(n29727), .Y(n21522) );
  INVX1 U29568 ( .A(reg_file[3606]), .Y(n29727) );
  NOR2X1 U29569 ( .A(n26064), .B(n29685), .Y(n21521) );
  INVX1 U29570 ( .A(reg_file[3607]), .Y(n29685) );
  NOR2X1 U29571 ( .A(n26064), .B(n29643), .Y(n21520) );
  INVX1 U29572 ( .A(reg_file[3608]), .Y(n29643) );
  NOR2X1 U29573 ( .A(n26064), .B(n29601), .Y(n21519) );
  INVX1 U29574 ( .A(reg_file[3609]), .Y(n29601) );
  NOR2X1 U29575 ( .A(n26064), .B(n29559), .Y(n21518) );
  INVX1 U29576 ( .A(reg_file[3610]), .Y(n29559) );
  NOR2X1 U29577 ( .A(n26064), .B(n29517), .Y(n21517) );
  INVX1 U29578 ( .A(reg_file[3611]), .Y(n29517) );
  NOR2X1 U29579 ( .A(n26064), .B(n29475), .Y(n21516) );
  INVX1 U29580 ( .A(reg_file[3612]), .Y(n29475) );
  NOR2X1 U29581 ( .A(n26064), .B(n29433), .Y(n21515) );
  INVX1 U29582 ( .A(reg_file[3613]), .Y(n29433) );
  NOR2X1 U29583 ( .A(n26064), .B(n29349), .Y(n21514) );
  INVX1 U29584 ( .A(reg_file[3614]), .Y(n29349) );
  NOR2X1 U29585 ( .A(n26065), .B(n29307), .Y(n21513) );
  INVX1 U29586 ( .A(reg_file[3615]), .Y(n29307) );
  NOR2X1 U29587 ( .A(n26065), .B(n29265), .Y(n21512) );
  INVX1 U29588 ( .A(reg_file[3616]), .Y(n29265) );
  NOR2X1 U29589 ( .A(n26065), .B(n29223), .Y(n21511) );
  INVX1 U29590 ( .A(reg_file[3617]), .Y(n29223) );
  NOR2X1 U29591 ( .A(n26065), .B(n29181), .Y(n21510) );
  INVX1 U29592 ( .A(reg_file[3618]), .Y(n29181) );
  NOR2X1 U29593 ( .A(n26065), .B(n29139), .Y(n21509) );
  INVX1 U29594 ( .A(reg_file[3619]), .Y(n29139) );
  NOR2X1 U29595 ( .A(n26065), .B(n29097), .Y(n21508) );
  INVX1 U29596 ( .A(reg_file[3620]), .Y(n29097) );
  NOR2X1 U29597 ( .A(n26065), .B(n29055), .Y(n21507) );
  INVX1 U29598 ( .A(reg_file[3621]), .Y(n29055) );
  NOR2X1 U29599 ( .A(n26065), .B(n29013), .Y(n21506) );
  INVX1 U29600 ( .A(reg_file[3622]), .Y(n29013) );
  NOR2X1 U29601 ( .A(n26065), .B(n28971), .Y(n21505) );
  INVX1 U29602 ( .A(reg_file[3623]), .Y(n28971) );
  NOR2X1 U29603 ( .A(n26065), .B(n28887), .Y(n21504) );
  INVX1 U29604 ( .A(reg_file[3624]), .Y(n28887) );
  NOR2X1 U29605 ( .A(n26065), .B(n28845), .Y(n21503) );
  INVX1 U29606 ( .A(reg_file[3625]), .Y(n28845) );
  NOR2X1 U29607 ( .A(n26065), .B(n28803), .Y(n21502) );
  INVX1 U29608 ( .A(reg_file[3626]), .Y(n28803) );
  NOR2X1 U29609 ( .A(n26065), .B(n28761), .Y(n21501) );
  INVX1 U29610 ( .A(reg_file[3627]), .Y(n28761) );
  NOR2X1 U29611 ( .A(n26065), .B(n28719), .Y(n21500) );
  INVX1 U29612 ( .A(reg_file[3628]), .Y(n28719) );
  NOR2X1 U29613 ( .A(n26065), .B(n28677), .Y(n21499) );
  INVX1 U29614 ( .A(reg_file[3629]), .Y(n28677) );
  NOR2X1 U29615 ( .A(n26065), .B(n28635), .Y(n21498) );
  INVX1 U29616 ( .A(reg_file[3630]), .Y(n28635) );
  NOR2X1 U29617 ( .A(n26065), .B(n28593), .Y(n21497) );
  INVX1 U29618 ( .A(reg_file[3631]), .Y(n28593) );
  NOR2X1 U29619 ( .A(n26066), .B(n28551), .Y(n21496) );
  INVX1 U29620 ( .A(reg_file[3632]), .Y(n28551) );
  NOR2X1 U29621 ( .A(n26066), .B(n28509), .Y(n21495) );
  INVX1 U29622 ( .A(reg_file[3633]), .Y(n28509) );
  NOR2X1 U29623 ( .A(n26066), .B(n28425), .Y(n21494) );
  INVX1 U29624 ( .A(reg_file[3634]), .Y(n28425) );
  NOR2X1 U29625 ( .A(n26066), .B(n28383), .Y(n21493) );
  INVX1 U29626 ( .A(reg_file[3635]), .Y(n28383) );
  NOR2X1 U29627 ( .A(n26066), .B(n28341), .Y(n21492) );
  INVX1 U29628 ( .A(reg_file[3636]), .Y(n28341) );
  NOR2X1 U29629 ( .A(n26066), .B(n28299), .Y(n21491) );
  INVX1 U29630 ( .A(reg_file[3637]), .Y(n28299) );
  NOR2X1 U29631 ( .A(n26066), .B(n28257), .Y(n21490) );
  INVX1 U29632 ( .A(reg_file[3638]), .Y(n28257) );
  NOR2X1 U29633 ( .A(n26066), .B(n28215), .Y(n21489) );
  INVX1 U29634 ( .A(reg_file[3639]), .Y(n28215) );
  NOR2X1 U29635 ( .A(n26066), .B(n28173), .Y(n21488) );
  INVX1 U29636 ( .A(reg_file[3640]), .Y(n28173) );
  NOR2X1 U29637 ( .A(n26066), .B(n28131), .Y(n21487) );
  INVX1 U29638 ( .A(reg_file[3641]), .Y(n28131) );
  NOR2X1 U29639 ( .A(n26066), .B(n28089), .Y(n21486) );
  INVX1 U29640 ( .A(reg_file[3642]), .Y(n28089) );
  NOR2X1 U29641 ( .A(n26066), .B(n28047), .Y(n21485) );
  INVX1 U29642 ( .A(reg_file[3643]), .Y(n28047) );
  NOR2X1 U29643 ( .A(n26066), .B(n27963), .Y(n21484) );
  INVX1 U29644 ( .A(reg_file[3644]), .Y(n27963) );
  NOR2X1 U29645 ( .A(n26066), .B(n27921), .Y(n21483) );
  INVX1 U29646 ( .A(reg_file[3645]), .Y(n27921) );
  NOR2X1 U29647 ( .A(n26066), .B(n27879), .Y(n21482) );
  INVX1 U29648 ( .A(reg_file[3646]), .Y(n27879) );
  NOR2X1 U29649 ( .A(n26066), .B(n27837), .Y(n21481) );
  INVX1 U29650 ( .A(reg_file[3647]), .Y(n27837) );
  NOR2X1 U29651 ( .A(n26066), .B(n27795), .Y(n21480) );
  INVX1 U29652 ( .A(reg_file[3648]), .Y(n27795) );
  NOR2X1 U29653 ( .A(n26067), .B(n27753), .Y(n21479) );
  INVX1 U29654 ( .A(reg_file[3649]), .Y(n27753) );
  NOR2X1 U29655 ( .A(n26067), .B(n27711), .Y(n21478) );
  INVX1 U29656 ( .A(reg_file[3650]), .Y(n27711) );
  NOR2X1 U29657 ( .A(n26067), .B(n27669), .Y(n21477) );
  INVX1 U29658 ( .A(reg_file[3651]), .Y(n27669) );
  NOR2X1 U29659 ( .A(n26067), .B(n27627), .Y(n21476) );
  INVX1 U29660 ( .A(reg_file[3652]), .Y(n27627) );
  NOR2X1 U29661 ( .A(n26067), .B(n27585), .Y(n21475) );
  INVX1 U29662 ( .A(reg_file[3653]), .Y(n27585) );
  NOR2X1 U29663 ( .A(n26067), .B(n27501), .Y(n21474) );
  INVX1 U29664 ( .A(reg_file[3654]), .Y(n27501) );
  NOR2X1 U29665 ( .A(n26067), .B(n27459), .Y(n21473) );
  INVX1 U29666 ( .A(reg_file[3655]), .Y(n27459) );
  NOR2X1 U29667 ( .A(n26067), .B(n27417), .Y(n21472) );
  INVX1 U29668 ( .A(reg_file[3656]), .Y(n27417) );
  NOR2X1 U29669 ( .A(n26067), .B(n27375), .Y(n21471) );
  INVX1 U29670 ( .A(reg_file[3657]), .Y(n27375) );
  NOR2X1 U29671 ( .A(n26067), .B(n27333), .Y(n21470) );
  INVX1 U29672 ( .A(reg_file[3658]), .Y(n27333) );
  NOR2X1 U29673 ( .A(n26067), .B(n27291), .Y(n21469) );
  INVX1 U29674 ( .A(reg_file[3659]), .Y(n27291) );
  NOR2X1 U29675 ( .A(n26067), .B(n27249), .Y(n21468) );
  INVX1 U29676 ( .A(reg_file[3660]), .Y(n27249) );
  NOR2X1 U29677 ( .A(n26067), .B(n27207), .Y(n21467) );
  INVX1 U29678 ( .A(reg_file[3661]), .Y(n27207) );
  NOR2X1 U29679 ( .A(n26067), .B(n27165), .Y(n21466) );
  INVX1 U29680 ( .A(reg_file[3662]), .Y(n27165) );
  NOR2X1 U29681 ( .A(n26067), .B(n27123), .Y(n21465) );
  INVX1 U29682 ( .A(reg_file[3663]), .Y(n27123) );
  NOR2X1 U29683 ( .A(n26067), .B(n27039), .Y(n21464) );
  INVX1 U29684 ( .A(reg_file[3664]), .Y(n27039) );
  NOR2X1 U29685 ( .A(n26067), .B(n26997), .Y(n21463) );
  INVX1 U29686 ( .A(reg_file[3665]), .Y(n26997) );
  NOR2X1 U29687 ( .A(n26068), .B(n26955), .Y(n21462) );
  INVX1 U29688 ( .A(reg_file[3666]), .Y(n26955) );
  NOR2X1 U29689 ( .A(n26068), .B(n26913), .Y(n21461) );
  INVX1 U29690 ( .A(reg_file[3667]), .Y(n26913) );
  NOR2X1 U29691 ( .A(n26068), .B(n26871), .Y(n21460) );
  INVX1 U29692 ( .A(reg_file[3668]), .Y(n26871) );
  NOR2X1 U29693 ( .A(n26068), .B(n26829), .Y(n21459) );
  INVX1 U29694 ( .A(reg_file[3669]), .Y(n26829) );
  NOR2X1 U29695 ( .A(n26068), .B(n26787), .Y(n21458) );
  INVX1 U29696 ( .A(reg_file[3670]), .Y(n26787) );
  NOR2X1 U29697 ( .A(n26068), .B(n26745), .Y(n21457) );
  INVX1 U29698 ( .A(reg_file[3671]), .Y(n26745) );
  NOR2X1 U29699 ( .A(n26068), .B(n26703), .Y(n21456) );
  INVX1 U29700 ( .A(reg_file[3672]), .Y(n26703) );
  NOR2X1 U29701 ( .A(n26068), .B(n26661), .Y(n21455) );
  INVX1 U29702 ( .A(reg_file[3673]), .Y(n26661) );
  NOR2X1 U29703 ( .A(n26068), .B(n26577), .Y(n21454) );
  INVX1 U29704 ( .A(reg_file[3674]), .Y(n26577) );
  NOR2X1 U29705 ( .A(n26068), .B(n26535), .Y(n21453) );
  INVX1 U29706 ( .A(reg_file[3675]), .Y(n26535) );
  NOR2X1 U29707 ( .A(n26068), .B(n26493), .Y(n21452) );
  INVX1 U29708 ( .A(reg_file[3676]), .Y(n26493) );
  NOR2X1 U29709 ( .A(n26068), .B(n26451), .Y(n21451) );
  INVX1 U29710 ( .A(reg_file[3677]), .Y(n26451) );
  NOR2X1 U29711 ( .A(n26068), .B(n26409), .Y(n21450) );
  INVX1 U29712 ( .A(reg_file[3678]), .Y(n26409) );
  NOR2X1 U29713 ( .A(n26068), .B(n26367), .Y(n21449) );
  INVX1 U29714 ( .A(reg_file[3679]), .Y(n26367) );
  NOR2X1 U29715 ( .A(n26068), .B(n26325), .Y(n21448) );
  INVX1 U29716 ( .A(reg_file[3680]), .Y(n26325) );
  NOR2X1 U29717 ( .A(n26068), .B(n26283), .Y(n21447) );
  INVX1 U29718 ( .A(reg_file[3681]), .Y(n26283) );
  NOR2X1 U29719 ( .A(n26068), .B(n26241), .Y(n21446) );
  INVX1 U29720 ( .A(reg_file[3682]), .Y(n26241) );
  NOR2X1 U29721 ( .A(n26069), .B(n26199), .Y(n21445) );
  INVX1 U29722 ( .A(reg_file[3683]), .Y(n26199) );
  NOR2X1 U29723 ( .A(n26069), .B(n31449), .Y(n21444) );
  INVX1 U29724 ( .A(reg_file[3684]), .Y(n31449) );
  NOR2X1 U29725 ( .A(n26069), .B(n31407), .Y(n21443) );
  INVX1 U29726 ( .A(reg_file[3685]), .Y(n31407) );
  NOR2X1 U29727 ( .A(n26069), .B(n31365), .Y(n21442) );
  INVX1 U29728 ( .A(reg_file[3686]), .Y(n31365) );
  NOR2X1 U29729 ( .A(n26069), .B(n31323), .Y(n21441) );
  INVX1 U29730 ( .A(reg_file[3687]), .Y(n31323) );
  NOR2X1 U29731 ( .A(n26069), .B(n31281), .Y(n21440) );
  INVX1 U29732 ( .A(reg_file[3688]), .Y(n31281) );
  NOR2X1 U29733 ( .A(n26069), .B(n31239), .Y(n21439) );
  INVX1 U29734 ( .A(reg_file[3689]), .Y(n31239) );
  NOR2X1 U29735 ( .A(n26069), .B(n31197), .Y(n21438) );
  INVX1 U29736 ( .A(reg_file[3690]), .Y(n31197) );
  NOR2X1 U29737 ( .A(n26069), .B(n31155), .Y(n21437) );
  INVX1 U29738 ( .A(reg_file[3691]), .Y(n31155) );
  NOR2X1 U29739 ( .A(n26069), .B(n31113), .Y(n21436) );
  INVX1 U29740 ( .A(reg_file[3692]), .Y(n31113) );
  NOR2X1 U29741 ( .A(n26069), .B(n31071), .Y(n21435) );
  INVX1 U29742 ( .A(reg_file[3693]), .Y(n31071) );
  NOR2X1 U29743 ( .A(n26069), .B(n30987), .Y(n21434) );
  INVX1 U29744 ( .A(reg_file[3694]), .Y(n30987) );
  NOR2X1 U29745 ( .A(n26069), .B(n30945), .Y(n21433) );
  INVX1 U29746 ( .A(reg_file[3695]), .Y(n30945) );
  NOR2X1 U29747 ( .A(n26069), .B(n30903), .Y(n21432) );
  INVX1 U29748 ( .A(reg_file[3696]), .Y(n30903) );
  NOR2X1 U29749 ( .A(n26069), .B(n30861), .Y(n21431) );
  INVX1 U29750 ( .A(reg_file[3697]), .Y(n30861) );
  NOR2X1 U29751 ( .A(n26069), .B(n30819), .Y(n21430) );
  INVX1 U29752 ( .A(reg_file[3698]), .Y(n30819) );
  NOR2X1 U29753 ( .A(n26069), .B(n30777), .Y(n21429) );
  INVX1 U29754 ( .A(reg_file[3699]), .Y(n30777) );
  NOR2X1 U29755 ( .A(n26070), .B(n30735), .Y(n21428) );
  INVX1 U29756 ( .A(reg_file[3700]), .Y(n30735) );
  NOR2X1 U29757 ( .A(n26070), .B(n30693), .Y(n21427) );
  INVX1 U29758 ( .A(reg_file[3701]), .Y(n30693) );
  NOR2X1 U29759 ( .A(n26070), .B(n30651), .Y(n21426) );
  INVX1 U29760 ( .A(reg_file[3702]), .Y(n30651) );
  NOR2X1 U29761 ( .A(n26070), .B(n30609), .Y(n21425) );
  INVX1 U29762 ( .A(reg_file[3703]), .Y(n30609) );
  NOR2X1 U29763 ( .A(n26070), .B(n30525), .Y(n21424) );
  INVX1 U29764 ( .A(reg_file[3704]), .Y(n30525) );
  NOR2X1 U29765 ( .A(n26070), .B(n30483), .Y(n21423) );
  INVX1 U29766 ( .A(reg_file[3705]), .Y(n30483) );
  NOR2X1 U29767 ( .A(n26070), .B(n30441), .Y(n21422) );
  INVX1 U29768 ( .A(reg_file[3706]), .Y(n30441) );
  NOR2X1 U29769 ( .A(n26070), .B(n30399), .Y(n21421) );
  INVX1 U29770 ( .A(reg_file[3707]), .Y(n30399) );
  NOR2X1 U29771 ( .A(n26070), .B(n30357), .Y(n21420) );
  INVX1 U29772 ( .A(reg_file[3708]), .Y(n30357) );
  NOR2X1 U29773 ( .A(n26070), .B(n30315), .Y(n21419) );
  INVX1 U29774 ( .A(reg_file[3709]), .Y(n30315) );
  NOR2X1 U29775 ( .A(n26070), .B(n30273), .Y(n21418) );
  INVX1 U29776 ( .A(reg_file[3710]), .Y(n30273) );
  NOR2X1 U29777 ( .A(n26070), .B(n30231), .Y(n21417) );
  INVX1 U29778 ( .A(reg_file[3711]), .Y(n30231) );
  NOR2X1 U29779 ( .A(n36623), .B(n35058), .Y(n37015) );
  MUX2X1 U29780 ( .B(n31507), .A(n25129), .S(n26071), .Y(n21416) );
  INVX1 U29781 ( .A(reg_file[3712]), .Y(n31507) );
  MUX2X1 U29782 ( .B(n29854), .A(n25130), .S(n26071), .Y(n21415) );
  INVX1 U29783 ( .A(reg_file[3713]), .Y(n29854) );
  MUX2X1 U29784 ( .B(n29392), .A(n25131), .S(n26071), .Y(n21414) );
  INVX1 U29785 ( .A(reg_file[3714]), .Y(n29392) );
  MUX2X1 U29786 ( .B(n28930), .A(n25132), .S(n26071), .Y(n21413) );
  INVX1 U29787 ( .A(reg_file[3715]), .Y(n28930) );
  MUX2X1 U29788 ( .B(n28468), .A(n25133), .S(n26071), .Y(n21412) );
  INVX1 U29789 ( .A(reg_file[3716]), .Y(n28468) );
  MUX2X1 U29790 ( .B(n28006), .A(n25134), .S(n26071), .Y(n21411) );
  INVX1 U29791 ( .A(reg_file[3717]), .Y(n28006) );
  MUX2X1 U29792 ( .B(n27544), .A(n25135), .S(n26071), .Y(n21410) );
  INVX1 U29793 ( .A(reg_file[3718]), .Y(n27544) );
  MUX2X1 U29794 ( .B(n27082), .A(n25136), .S(n26071), .Y(n21409) );
  INVX1 U29795 ( .A(reg_file[3719]), .Y(n27082) );
  NOR2X1 U29796 ( .A(n26071), .B(n26620), .Y(n21408) );
  INVX1 U29797 ( .A(reg_file[3720]), .Y(n26620) );
  NOR2X1 U29798 ( .A(n26071), .B(n26144), .Y(n21407) );
  INVX1 U29799 ( .A(reg_file[3721]), .Y(n26144) );
  NOR2X1 U29800 ( .A(n26071), .B(n31030), .Y(n21406) );
  INVX1 U29801 ( .A(reg_file[3722]), .Y(n31030) );
  NOR2X1 U29802 ( .A(n26071), .B(n30568), .Y(n21405) );
  INVX1 U29803 ( .A(reg_file[3723]), .Y(n30568) );
  NOR2X1 U29804 ( .A(n26071), .B(n30190), .Y(n21404) );
  INVX1 U29805 ( .A(reg_file[3724]), .Y(n30190) );
  NOR2X1 U29806 ( .A(n26071), .B(n30148), .Y(n21403) );
  INVX1 U29807 ( .A(reg_file[3725]), .Y(n30148) );
  NOR2X1 U29808 ( .A(n26072), .B(n30106), .Y(n21402) );
  INVX1 U29809 ( .A(reg_file[3726]), .Y(n30106) );
  NOR2X1 U29810 ( .A(n26072), .B(n30064), .Y(n21401) );
  INVX1 U29811 ( .A(reg_file[3727]), .Y(n30064) );
  NOR2X1 U29812 ( .A(n26072), .B(n30022), .Y(n21400) );
  INVX1 U29813 ( .A(reg_file[3728]), .Y(n30022) );
  NOR2X1 U29814 ( .A(n26072), .B(n29980), .Y(n21399) );
  INVX1 U29815 ( .A(reg_file[3729]), .Y(n29980) );
  NOR2X1 U29816 ( .A(n26072), .B(n29938), .Y(n21398) );
  INVX1 U29817 ( .A(reg_file[3730]), .Y(n29938) );
  NOR2X1 U29818 ( .A(n26072), .B(n29896), .Y(n21397) );
  INVX1 U29819 ( .A(reg_file[3731]), .Y(n29896) );
  NOR2X1 U29820 ( .A(n26072), .B(n29812), .Y(n21396) );
  INVX1 U29821 ( .A(reg_file[3732]), .Y(n29812) );
  NOR2X1 U29822 ( .A(n26072), .B(n29770), .Y(n21395) );
  INVX1 U29823 ( .A(reg_file[3733]), .Y(n29770) );
  NOR2X1 U29824 ( .A(n26072), .B(n29728), .Y(n21394) );
  INVX1 U29825 ( .A(reg_file[3734]), .Y(n29728) );
  NOR2X1 U29826 ( .A(n26072), .B(n29686), .Y(n21393) );
  INVX1 U29827 ( .A(reg_file[3735]), .Y(n29686) );
  NOR2X1 U29828 ( .A(n26072), .B(n29644), .Y(n21392) );
  INVX1 U29829 ( .A(reg_file[3736]), .Y(n29644) );
  NOR2X1 U29830 ( .A(n26072), .B(n29602), .Y(n21391) );
  INVX1 U29831 ( .A(reg_file[3737]), .Y(n29602) );
  NOR2X1 U29832 ( .A(n26072), .B(n29560), .Y(n21390) );
  INVX1 U29833 ( .A(reg_file[3738]), .Y(n29560) );
  NOR2X1 U29834 ( .A(n26072), .B(n29518), .Y(n21389) );
  INVX1 U29835 ( .A(reg_file[3739]), .Y(n29518) );
  NOR2X1 U29836 ( .A(n26072), .B(n29476), .Y(n21388) );
  INVX1 U29837 ( .A(reg_file[3740]), .Y(n29476) );
  NOR2X1 U29838 ( .A(n26072), .B(n29434), .Y(n21387) );
  INVX1 U29839 ( .A(reg_file[3741]), .Y(n29434) );
  NOR2X1 U29840 ( .A(n26072), .B(n29350), .Y(n21386) );
  INVX1 U29841 ( .A(reg_file[3742]), .Y(n29350) );
  NOR2X1 U29842 ( .A(n26073), .B(n29308), .Y(n21385) );
  INVX1 U29843 ( .A(reg_file[3743]), .Y(n29308) );
  NOR2X1 U29844 ( .A(n26073), .B(n29266), .Y(n21384) );
  INVX1 U29845 ( .A(reg_file[3744]), .Y(n29266) );
  NOR2X1 U29846 ( .A(n26073), .B(n29224), .Y(n21383) );
  INVX1 U29847 ( .A(reg_file[3745]), .Y(n29224) );
  NOR2X1 U29848 ( .A(n26073), .B(n29182), .Y(n21382) );
  INVX1 U29849 ( .A(reg_file[3746]), .Y(n29182) );
  NOR2X1 U29850 ( .A(n26073), .B(n29140), .Y(n21381) );
  INVX1 U29851 ( .A(reg_file[3747]), .Y(n29140) );
  NOR2X1 U29852 ( .A(n26073), .B(n29098), .Y(n21380) );
  INVX1 U29853 ( .A(reg_file[3748]), .Y(n29098) );
  NOR2X1 U29854 ( .A(n26073), .B(n29056), .Y(n21379) );
  INVX1 U29855 ( .A(reg_file[3749]), .Y(n29056) );
  NOR2X1 U29856 ( .A(n26073), .B(n29014), .Y(n21378) );
  INVX1 U29857 ( .A(reg_file[3750]), .Y(n29014) );
  NOR2X1 U29858 ( .A(n26073), .B(n28972), .Y(n21377) );
  INVX1 U29859 ( .A(reg_file[3751]), .Y(n28972) );
  NOR2X1 U29860 ( .A(n26073), .B(n28888), .Y(n21376) );
  INVX1 U29861 ( .A(reg_file[3752]), .Y(n28888) );
  NOR2X1 U29862 ( .A(n26073), .B(n28846), .Y(n21375) );
  INVX1 U29863 ( .A(reg_file[3753]), .Y(n28846) );
  NOR2X1 U29864 ( .A(n26073), .B(n28804), .Y(n21374) );
  INVX1 U29865 ( .A(reg_file[3754]), .Y(n28804) );
  NOR2X1 U29866 ( .A(n26073), .B(n28762), .Y(n21373) );
  INVX1 U29867 ( .A(reg_file[3755]), .Y(n28762) );
  NOR2X1 U29868 ( .A(n26073), .B(n28720), .Y(n21372) );
  INVX1 U29869 ( .A(reg_file[3756]), .Y(n28720) );
  NOR2X1 U29870 ( .A(n26073), .B(n28678), .Y(n21371) );
  INVX1 U29871 ( .A(reg_file[3757]), .Y(n28678) );
  NOR2X1 U29872 ( .A(n26073), .B(n28636), .Y(n21370) );
  INVX1 U29873 ( .A(reg_file[3758]), .Y(n28636) );
  NOR2X1 U29874 ( .A(n26073), .B(n28594), .Y(n21369) );
  INVX1 U29875 ( .A(reg_file[3759]), .Y(n28594) );
  NOR2X1 U29876 ( .A(n26074), .B(n28552), .Y(n21368) );
  INVX1 U29877 ( .A(reg_file[3760]), .Y(n28552) );
  NOR2X1 U29878 ( .A(n26074), .B(n28510), .Y(n21367) );
  INVX1 U29879 ( .A(reg_file[3761]), .Y(n28510) );
  NOR2X1 U29880 ( .A(n26074), .B(n28426), .Y(n21366) );
  INVX1 U29881 ( .A(reg_file[3762]), .Y(n28426) );
  NOR2X1 U29882 ( .A(n26074), .B(n28384), .Y(n21365) );
  INVX1 U29883 ( .A(reg_file[3763]), .Y(n28384) );
  NOR2X1 U29884 ( .A(n26074), .B(n28342), .Y(n21364) );
  INVX1 U29885 ( .A(reg_file[3764]), .Y(n28342) );
  NOR2X1 U29886 ( .A(n26074), .B(n28300), .Y(n21363) );
  INVX1 U29887 ( .A(reg_file[3765]), .Y(n28300) );
  NOR2X1 U29888 ( .A(n26074), .B(n28258), .Y(n21362) );
  INVX1 U29889 ( .A(reg_file[3766]), .Y(n28258) );
  NOR2X1 U29890 ( .A(n26074), .B(n28216), .Y(n21361) );
  INVX1 U29891 ( .A(reg_file[3767]), .Y(n28216) );
  NOR2X1 U29892 ( .A(n26074), .B(n28174), .Y(n21360) );
  INVX1 U29893 ( .A(reg_file[3768]), .Y(n28174) );
  NOR2X1 U29894 ( .A(n26074), .B(n28132), .Y(n21359) );
  INVX1 U29895 ( .A(reg_file[3769]), .Y(n28132) );
  NOR2X1 U29896 ( .A(n26074), .B(n28090), .Y(n21358) );
  INVX1 U29897 ( .A(reg_file[3770]), .Y(n28090) );
  NOR2X1 U29898 ( .A(n26074), .B(n28048), .Y(n21357) );
  INVX1 U29899 ( .A(reg_file[3771]), .Y(n28048) );
  NOR2X1 U29900 ( .A(n26074), .B(n27964), .Y(n21356) );
  INVX1 U29901 ( .A(reg_file[3772]), .Y(n27964) );
  NOR2X1 U29902 ( .A(n26074), .B(n27922), .Y(n21355) );
  INVX1 U29903 ( .A(reg_file[3773]), .Y(n27922) );
  NOR2X1 U29904 ( .A(n26074), .B(n27880), .Y(n21354) );
  INVX1 U29905 ( .A(reg_file[3774]), .Y(n27880) );
  NOR2X1 U29906 ( .A(n26074), .B(n27838), .Y(n21353) );
  INVX1 U29907 ( .A(reg_file[3775]), .Y(n27838) );
  NOR2X1 U29908 ( .A(n26074), .B(n27796), .Y(n21352) );
  INVX1 U29909 ( .A(reg_file[3776]), .Y(n27796) );
  NOR2X1 U29910 ( .A(n26075), .B(n27754), .Y(n21351) );
  INVX1 U29911 ( .A(reg_file[3777]), .Y(n27754) );
  NOR2X1 U29912 ( .A(n26075), .B(n27712), .Y(n21350) );
  INVX1 U29913 ( .A(reg_file[3778]), .Y(n27712) );
  NOR2X1 U29914 ( .A(n26075), .B(n27670), .Y(n21349) );
  INVX1 U29915 ( .A(reg_file[3779]), .Y(n27670) );
  NOR2X1 U29916 ( .A(n26075), .B(n27628), .Y(n21348) );
  INVX1 U29917 ( .A(reg_file[3780]), .Y(n27628) );
  NOR2X1 U29918 ( .A(n26075), .B(n27586), .Y(n21347) );
  INVX1 U29919 ( .A(reg_file[3781]), .Y(n27586) );
  NOR2X1 U29920 ( .A(n26075), .B(n27502), .Y(n21346) );
  INVX1 U29921 ( .A(reg_file[3782]), .Y(n27502) );
  NOR2X1 U29922 ( .A(n26075), .B(n27460), .Y(n21345) );
  INVX1 U29923 ( .A(reg_file[3783]), .Y(n27460) );
  NOR2X1 U29924 ( .A(n26075), .B(n27418), .Y(n21344) );
  INVX1 U29925 ( .A(reg_file[3784]), .Y(n27418) );
  NOR2X1 U29926 ( .A(n26075), .B(n27376), .Y(n21343) );
  INVX1 U29927 ( .A(reg_file[3785]), .Y(n27376) );
  NOR2X1 U29928 ( .A(n26075), .B(n27334), .Y(n21342) );
  INVX1 U29929 ( .A(reg_file[3786]), .Y(n27334) );
  NOR2X1 U29930 ( .A(n26075), .B(n27292), .Y(n21341) );
  INVX1 U29931 ( .A(reg_file[3787]), .Y(n27292) );
  NOR2X1 U29932 ( .A(n26075), .B(n27250), .Y(n21340) );
  INVX1 U29933 ( .A(reg_file[3788]), .Y(n27250) );
  NOR2X1 U29934 ( .A(n26075), .B(n27208), .Y(n21339) );
  INVX1 U29935 ( .A(reg_file[3789]), .Y(n27208) );
  NOR2X1 U29936 ( .A(n26075), .B(n27166), .Y(n21338) );
  INVX1 U29937 ( .A(reg_file[3790]), .Y(n27166) );
  NOR2X1 U29938 ( .A(n26075), .B(n27124), .Y(n21337) );
  INVX1 U29939 ( .A(reg_file[3791]), .Y(n27124) );
  NOR2X1 U29940 ( .A(n26075), .B(n27040), .Y(n21336) );
  INVX1 U29941 ( .A(reg_file[3792]), .Y(n27040) );
  NOR2X1 U29942 ( .A(n26075), .B(n26998), .Y(n21335) );
  INVX1 U29943 ( .A(reg_file[3793]), .Y(n26998) );
  NOR2X1 U29944 ( .A(n26076), .B(n26956), .Y(n21334) );
  INVX1 U29945 ( .A(reg_file[3794]), .Y(n26956) );
  NOR2X1 U29946 ( .A(n26076), .B(n26914), .Y(n21333) );
  INVX1 U29947 ( .A(reg_file[3795]), .Y(n26914) );
  NOR2X1 U29948 ( .A(n26076), .B(n26872), .Y(n21332) );
  INVX1 U29949 ( .A(reg_file[3796]), .Y(n26872) );
  NOR2X1 U29950 ( .A(n26076), .B(n26830), .Y(n21331) );
  INVX1 U29951 ( .A(reg_file[3797]), .Y(n26830) );
  NOR2X1 U29952 ( .A(n26076), .B(n26788), .Y(n21330) );
  INVX1 U29953 ( .A(reg_file[3798]), .Y(n26788) );
  NOR2X1 U29954 ( .A(n26076), .B(n26746), .Y(n21329) );
  INVX1 U29955 ( .A(reg_file[3799]), .Y(n26746) );
  NOR2X1 U29956 ( .A(n26076), .B(n26704), .Y(n21328) );
  INVX1 U29957 ( .A(reg_file[3800]), .Y(n26704) );
  NOR2X1 U29958 ( .A(n26076), .B(n26662), .Y(n21327) );
  INVX1 U29959 ( .A(reg_file[3801]), .Y(n26662) );
  NOR2X1 U29960 ( .A(n26076), .B(n26578), .Y(n21326) );
  INVX1 U29961 ( .A(reg_file[3802]), .Y(n26578) );
  NOR2X1 U29962 ( .A(n26076), .B(n26536), .Y(n21325) );
  INVX1 U29963 ( .A(reg_file[3803]), .Y(n26536) );
  NOR2X1 U29964 ( .A(n26076), .B(n26494), .Y(n21324) );
  INVX1 U29965 ( .A(reg_file[3804]), .Y(n26494) );
  NOR2X1 U29966 ( .A(n26076), .B(n26452), .Y(n21323) );
  INVX1 U29967 ( .A(reg_file[3805]), .Y(n26452) );
  NOR2X1 U29968 ( .A(n26076), .B(n26410), .Y(n21322) );
  INVX1 U29969 ( .A(reg_file[3806]), .Y(n26410) );
  NOR2X1 U29970 ( .A(n26076), .B(n26368), .Y(n21321) );
  INVX1 U29971 ( .A(reg_file[3807]), .Y(n26368) );
  NOR2X1 U29972 ( .A(n26076), .B(n26326), .Y(n21320) );
  INVX1 U29973 ( .A(reg_file[3808]), .Y(n26326) );
  NOR2X1 U29974 ( .A(n26076), .B(n26284), .Y(n21319) );
  INVX1 U29975 ( .A(reg_file[3809]), .Y(n26284) );
  NOR2X1 U29976 ( .A(n26076), .B(n26242), .Y(n21318) );
  INVX1 U29977 ( .A(reg_file[3810]), .Y(n26242) );
  NOR2X1 U29978 ( .A(n26077), .B(n26200), .Y(n21317) );
  INVX1 U29979 ( .A(reg_file[3811]), .Y(n26200) );
  NOR2X1 U29980 ( .A(n26077), .B(n31450), .Y(n21316) );
  INVX1 U29981 ( .A(reg_file[3812]), .Y(n31450) );
  NOR2X1 U29982 ( .A(n26077), .B(n31408), .Y(n21315) );
  INVX1 U29983 ( .A(reg_file[3813]), .Y(n31408) );
  NOR2X1 U29984 ( .A(n26077), .B(n31366), .Y(n21314) );
  INVX1 U29985 ( .A(reg_file[3814]), .Y(n31366) );
  NOR2X1 U29986 ( .A(n26077), .B(n31324), .Y(n21313) );
  INVX1 U29987 ( .A(reg_file[3815]), .Y(n31324) );
  NOR2X1 U29988 ( .A(n26077), .B(n31282), .Y(n21312) );
  INVX1 U29989 ( .A(reg_file[3816]), .Y(n31282) );
  NOR2X1 U29990 ( .A(n26077), .B(n31240), .Y(n21311) );
  INVX1 U29991 ( .A(reg_file[3817]), .Y(n31240) );
  NOR2X1 U29992 ( .A(n26077), .B(n31198), .Y(n21310) );
  INVX1 U29993 ( .A(reg_file[3818]), .Y(n31198) );
  NOR2X1 U29994 ( .A(n26077), .B(n31156), .Y(n21309) );
  INVX1 U29995 ( .A(reg_file[3819]), .Y(n31156) );
  NOR2X1 U29996 ( .A(n26077), .B(n31114), .Y(n21308) );
  INVX1 U29997 ( .A(reg_file[3820]), .Y(n31114) );
  NOR2X1 U29998 ( .A(n26077), .B(n31072), .Y(n21307) );
  INVX1 U29999 ( .A(reg_file[3821]), .Y(n31072) );
  NOR2X1 U30000 ( .A(n26077), .B(n30988), .Y(n21306) );
  INVX1 U30001 ( .A(reg_file[3822]), .Y(n30988) );
  NOR2X1 U30002 ( .A(n26077), .B(n30946), .Y(n21305) );
  INVX1 U30003 ( .A(reg_file[3823]), .Y(n30946) );
  NOR2X1 U30004 ( .A(n26077), .B(n30904), .Y(n21304) );
  INVX1 U30005 ( .A(reg_file[3824]), .Y(n30904) );
  NOR2X1 U30006 ( .A(n26077), .B(n30862), .Y(n21303) );
  INVX1 U30007 ( .A(reg_file[3825]), .Y(n30862) );
  NOR2X1 U30008 ( .A(n26077), .B(n30820), .Y(n21302) );
  INVX1 U30009 ( .A(reg_file[3826]), .Y(n30820) );
  NOR2X1 U30010 ( .A(n26077), .B(n30778), .Y(n21301) );
  INVX1 U30011 ( .A(reg_file[3827]), .Y(n30778) );
  NOR2X1 U30012 ( .A(n26078), .B(n30736), .Y(n21300) );
  INVX1 U30013 ( .A(reg_file[3828]), .Y(n30736) );
  NOR2X1 U30014 ( .A(n26078), .B(n30694), .Y(n21299) );
  INVX1 U30015 ( .A(reg_file[3829]), .Y(n30694) );
  NOR2X1 U30016 ( .A(n26078), .B(n30652), .Y(n21298) );
  INVX1 U30017 ( .A(reg_file[3830]), .Y(n30652) );
  NOR2X1 U30018 ( .A(n26078), .B(n30610), .Y(n21297) );
  INVX1 U30019 ( .A(reg_file[3831]), .Y(n30610) );
  NOR2X1 U30020 ( .A(n26078), .B(n30526), .Y(n21296) );
  INVX1 U30021 ( .A(reg_file[3832]), .Y(n30526) );
  NOR2X1 U30022 ( .A(n26078), .B(n30484), .Y(n21295) );
  INVX1 U30023 ( .A(reg_file[3833]), .Y(n30484) );
  NOR2X1 U30024 ( .A(n26078), .B(n30442), .Y(n21294) );
  INVX1 U30025 ( .A(reg_file[3834]), .Y(n30442) );
  NOR2X1 U30026 ( .A(n26078), .B(n30400), .Y(n21293) );
  INVX1 U30027 ( .A(reg_file[3835]), .Y(n30400) );
  NOR2X1 U30028 ( .A(n26078), .B(n30358), .Y(n21292) );
  INVX1 U30029 ( .A(reg_file[3836]), .Y(n30358) );
  NOR2X1 U30030 ( .A(n26078), .B(n30316), .Y(n21291) );
  INVX1 U30031 ( .A(reg_file[3837]), .Y(n30316) );
  NOR2X1 U30032 ( .A(n26078), .B(n30274), .Y(n21290) );
  INVX1 U30033 ( .A(reg_file[3838]), .Y(n30274) );
  NOR2X1 U30034 ( .A(n26078), .B(n30232), .Y(n21289) );
  INVX1 U30035 ( .A(reg_file[3839]), .Y(n30232) );
  NOR2X1 U30036 ( .A(n36753), .B(n35058), .Y(n37016) );
  NAND3X1 U30037 ( .A(n36756), .B(n36754), .C(wraddr[2]), .Y(n35058) );
  INVX1 U30038 ( .A(wraddr[1]), .Y(n36754) );
  MUX2X1 U30039 ( .B(n31510), .A(n25129), .S(n26079), .Y(n21288) );
  INVX1 U30040 ( .A(reg_file[3840]), .Y(n31510) );
  MUX2X1 U30041 ( .B(n29855), .A(n25130), .S(n26079), .Y(n21287) );
  INVX1 U30042 ( .A(reg_file[3841]), .Y(n29855) );
  MUX2X1 U30043 ( .B(n29393), .A(n25131), .S(n26079), .Y(n21286) );
  INVX1 U30044 ( .A(reg_file[3842]), .Y(n29393) );
  MUX2X1 U30045 ( .B(n28931), .A(n25132), .S(n26079), .Y(n21285) );
  INVX1 U30046 ( .A(reg_file[3843]), .Y(n28931) );
  MUX2X1 U30047 ( .B(n28469), .A(n25133), .S(n26079), .Y(n21284) );
  INVX1 U30048 ( .A(reg_file[3844]), .Y(n28469) );
  MUX2X1 U30049 ( .B(n28007), .A(n25134), .S(n26079), .Y(n21283) );
  INVX1 U30050 ( .A(reg_file[3845]), .Y(n28007) );
  MUX2X1 U30051 ( .B(n27545), .A(n25135), .S(n26079), .Y(n21282) );
  INVX1 U30052 ( .A(reg_file[3846]), .Y(n27545) );
  MUX2X1 U30053 ( .B(n27083), .A(n25136), .S(n26079), .Y(n21281) );
  INVX1 U30054 ( .A(reg_file[3847]), .Y(n27083) );
  NOR2X1 U30055 ( .A(n26079), .B(n26621), .Y(n21280) );
  INVX1 U30056 ( .A(reg_file[3848]), .Y(n26621) );
  NOR2X1 U30057 ( .A(n26079), .B(n26146), .Y(n21279) );
  INVX1 U30058 ( .A(reg_file[3849]), .Y(n26146) );
  NOR2X1 U30059 ( .A(n26079), .B(n31031), .Y(n21278) );
  INVX1 U30060 ( .A(reg_file[3850]), .Y(n31031) );
  NOR2X1 U30061 ( .A(n26079), .B(n30569), .Y(n21277) );
  INVX1 U30062 ( .A(reg_file[3851]), .Y(n30569) );
  NOR2X1 U30063 ( .A(n26079), .B(n30191), .Y(n21276) );
  INVX1 U30064 ( .A(reg_file[3852]), .Y(n30191) );
  NOR2X1 U30065 ( .A(n26079), .B(n30149), .Y(n21275) );
  INVX1 U30066 ( .A(reg_file[3853]), .Y(n30149) );
  NOR2X1 U30067 ( .A(n26080), .B(n30107), .Y(n21274) );
  INVX1 U30068 ( .A(reg_file[3854]), .Y(n30107) );
  NOR2X1 U30069 ( .A(n26080), .B(n30065), .Y(n21273) );
  INVX1 U30070 ( .A(reg_file[3855]), .Y(n30065) );
  NOR2X1 U30071 ( .A(n26080), .B(n30023), .Y(n21272) );
  INVX1 U30072 ( .A(reg_file[3856]), .Y(n30023) );
  NOR2X1 U30073 ( .A(n26080), .B(n29981), .Y(n21271) );
  INVX1 U30074 ( .A(reg_file[3857]), .Y(n29981) );
  NOR2X1 U30075 ( .A(n26080), .B(n29939), .Y(n21270) );
  INVX1 U30076 ( .A(reg_file[3858]), .Y(n29939) );
  NOR2X1 U30077 ( .A(n26080), .B(n29897), .Y(n21269) );
  INVX1 U30078 ( .A(reg_file[3859]), .Y(n29897) );
  NOR2X1 U30079 ( .A(n26080), .B(n29813), .Y(n21268) );
  INVX1 U30080 ( .A(reg_file[3860]), .Y(n29813) );
  NOR2X1 U30081 ( .A(n26080), .B(n29771), .Y(n21267) );
  INVX1 U30082 ( .A(reg_file[3861]), .Y(n29771) );
  NOR2X1 U30083 ( .A(n26080), .B(n29729), .Y(n21266) );
  INVX1 U30084 ( .A(reg_file[3862]), .Y(n29729) );
  NOR2X1 U30085 ( .A(n26080), .B(n29687), .Y(n21265) );
  INVX1 U30086 ( .A(reg_file[3863]), .Y(n29687) );
  NOR2X1 U30087 ( .A(n26080), .B(n29645), .Y(n21264) );
  INVX1 U30088 ( .A(reg_file[3864]), .Y(n29645) );
  NOR2X1 U30089 ( .A(n26080), .B(n29603), .Y(n21263) );
  INVX1 U30090 ( .A(reg_file[3865]), .Y(n29603) );
  NOR2X1 U30091 ( .A(n26080), .B(n29561), .Y(n21262) );
  INVX1 U30092 ( .A(reg_file[3866]), .Y(n29561) );
  NOR2X1 U30093 ( .A(n26080), .B(n29519), .Y(n21261) );
  INVX1 U30094 ( .A(reg_file[3867]), .Y(n29519) );
  NOR2X1 U30095 ( .A(n26080), .B(n29477), .Y(n21260) );
  INVX1 U30096 ( .A(reg_file[3868]), .Y(n29477) );
  NOR2X1 U30097 ( .A(n26080), .B(n29435), .Y(n21259) );
  INVX1 U30098 ( .A(reg_file[3869]), .Y(n29435) );
  NOR2X1 U30099 ( .A(n26080), .B(n29351), .Y(n21258) );
  INVX1 U30100 ( .A(reg_file[3870]), .Y(n29351) );
  NOR2X1 U30101 ( .A(n26081), .B(n29309), .Y(n21257) );
  INVX1 U30102 ( .A(reg_file[3871]), .Y(n29309) );
  NOR2X1 U30103 ( .A(n26081), .B(n29267), .Y(n21256) );
  INVX1 U30104 ( .A(reg_file[3872]), .Y(n29267) );
  NOR2X1 U30105 ( .A(n26081), .B(n29225), .Y(n21255) );
  INVX1 U30106 ( .A(reg_file[3873]), .Y(n29225) );
  NOR2X1 U30107 ( .A(n26081), .B(n29183), .Y(n21254) );
  INVX1 U30108 ( .A(reg_file[3874]), .Y(n29183) );
  NOR2X1 U30109 ( .A(n26081), .B(n29141), .Y(n21253) );
  INVX1 U30110 ( .A(reg_file[3875]), .Y(n29141) );
  NOR2X1 U30111 ( .A(n26081), .B(n29099), .Y(n21252) );
  INVX1 U30112 ( .A(reg_file[3876]), .Y(n29099) );
  NOR2X1 U30113 ( .A(n26081), .B(n29057), .Y(n21251) );
  INVX1 U30114 ( .A(reg_file[3877]), .Y(n29057) );
  NOR2X1 U30115 ( .A(n26081), .B(n29015), .Y(n21250) );
  INVX1 U30116 ( .A(reg_file[3878]), .Y(n29015) );
  NOR2X1 U30117 ( .A(n26081), .B(n28973), .Y(n21249) );
  INVX1 U30118 ( .A(reg_file[3879]), .Y(n28973) );
  NOR2X1 U30119 ( .A(n26081), .B(n28889), .Y(n21248) );
  INVX1 U30120 ( .A(reg_file[3880]), .Y(n28889) );
  NOR2X1 U30121 ( .A(n26081), .B(n28847), .Y(n21247) );
  INVX1 U30122 ( .A(reg_file[3881]), .Y(n28847) );
  NOR2X1 U30123 ( .A(n26081), .B(n28805), .Y(n21246) );
  INVX1 U30124 ( .A(reg_file[3882]), .Y(n28805) );
  NOR2X1 U30125 ( .A(n26081), .B(n28763), .Y(n21245) );
  INVX1 U30126 ( .A(reg_file[3883]), .Y(n28763) );
  NOR2X1 U30127 ( .A(n26081), .B(n28721), .Y(n21244) );
  INVX1 U30128 ( .A(reg_file[3884]), .Y(n28721) );
  NOR2X1 U30129 ( .A(n26081), .B(n28679), .Y(n21243) );
  INVX1 U30130 ( .A(reg_file[3885]), .Y(n28679) );
  NOR2X1 U30131 ( .A(n26081), .B(n28637), .Y(n21242) );
  INVX1 U30132 ( .A(reg_file[3886]), .Y(n28637) );
  NOR2X1 U30133 ( .A(n26081), .B(n28595), .Y(n21241) );
  INVX1 U30134 ( .A(reg_file[3887]), .Y(n28595) );
  NOR2X1 U30135 ( .A(n26082), .B(n28553), .Y(n21240) );
  INVX1 U30136 ( .A(reg_file[3888]), .Y(n28553) );
  NOR2X1 U30137 ( .A(n26082), .B(n28511), .Y(n21239) );
  INVX1 U30138 ( .A(reg_file[3889]), .Y(n28511) );
  NOR2X1 U30139 ( .A(n26082), .B(n28427), .Y(n21238) );
  INVX1 U30140 ( .A(reg_file[3890]), .Y(n28427) );
  NOR2X1 U30141 ( .A(n26082), .B(n28385), .Y(n21237) );
  INVX1 U30142 ( .A(reg_file[3891]), .Y(n28385) );
  NOR2X1 U30143 ( .A(n26082), .B(n28343), .Y(n21236) );
  INVX1 U30144 ( .A(reg_file[3892]), .Y(n28343) );
  NOR2X1 U30145 ( .A(n26082), .B(n28301), .Y(n21235) );
  INVX1 U30146 ( .A(reg_file[3893]), .Y(n28301) );
  NOR2X1 U30147 ( .A(n26082), .B(n28259), .Y(n21234) );
  INVX1 U30148 ( .A(reg_file[3894]), .Y(n28259) );
  NOR2X1 U30149 ( .A(n26082), .B(n28217), .Y(n21233) );
  INVX1 U30150 ( .A(reg_file[3895]), .Y(n28217) );
  NOR2X1 U30151 ( .A(n26082), .B(n28175), .Y(n21232) );
  INVX1 U30152 ( .A(reg_file[3896]), .Y(n28175) );
  NOR2X1 U30153 ( .A(n26082), .B(n28133), .Y(n21231) );
  INVX1 U30154 ( .A(reg_file[3897]), .Y(n28133) );
  NOR2X1 U30155 ( .A(n26082), .B(n28091), .Y(n21230) );
  INVX1 U30156 ( .A(reg_file[3898]), .Y(n28091) );
  NOR2X1 U30157 ( .A(n26082), .B(n28049), .Y(n21229) );
  INVX1 U30158 ( .A(reg_file[3899]), .Y(n28049) );
  NOR2X1 U30159 ( .A(n26082), .B(n27965), .Y(n21228) );
  INVX1 U30160 ( .A(reg_file[3900]), .Y(n27965) );
  NOR2X1 U30161 ( .A(n26082), .B(n27923), .Y(n21227) );
  INVX1 U30162 ( .A(reg_file[3901]), .Y(n27923) );
  NOR2X1 U30163 ( .A(n26082), .B(n27881), .Y(n21226) );
  INVX1 U30164 ( .A(reg_file[3902]), .Y(n27881) );
  NOR2X1 U30165 ( .A(n26082), .B(n27839), .Y(n21225) );
  INVX1 U30166 ( .A(reg_file[3903]), .Y(n27839) );
  NOR2X1 U30167 ( .A(n26082), .B(n27797), .Y(n21224) );
  INVX1 U30168 ( .A(reg_file[3904]), .Y(n27797) );
  NOR2X1 U30169 ( .A(n26083), .B(n27755), .Y(n21223) );
  INVX1 U30170 ( .A(reg_file[3905]), .Y(n27755) );
  NOR2X1 U30171 ( .A(n26083), .B(n27713), .Y(n21222) );
  INVX1 U30172 ( .A(reg_file[3906]), .Y(n27713) );
  NOR2X1 U30173 ( .A(n26083), .B(n27671), .Y(n21221) );
  INVX1 U30174 ( .A(reg_file[3907]), .Y(n27671) );
  NOR2X1 U30175 ( .A(n26083), .B(n27629), .Y(n21220) );
  INVX1 U30176 ( .A(reg_file[3908]), .Y(n27629) );
  NOR2X1 U30177 ( .A(n26083), .B(n27587), .Y(n21219) );
  INVX1 U30178 ( .A(reg_file[3909]), .Y(n27587) );
  NOR2X1 U30179 ( .A(n26083), .B(n27503), .Y(n21218) );
  INVX1 U30180 ( .A(reg_file[3910]), .Y(n27503) );
  NOR2X1 U30181 ( .A(n26083), .B(n27461), .Y(n21217) );
  INVX1 U30182 ( .A(reg_file[3911]), .Y(n27461) );
  NOR2X1 U30183 ( .A(n26083), .B(n27419), .Y(n21216) );
  INVX1 U30184 ( .A(reg_file[3912]), .Y(n27419) );
  NOR2X1 U30185 ( .A(n26083), .B(n27377), .Y(n21215) );
  INVX1 U30186 ( .A(reg_file[3913]), .Y(n27377) );
  NOR2X1 U30187 ( .A(n26083), .B(n27335), .Y(n21214) );
  INVX1 U30188 ( .A(reg_file[3914]), .Y(n27335) );
  NOR2X1 U30189 ( .A(n26083), .B(n27293), .Y(n21213) );
  INVX1 U30190 ( .A(reg_file[3915]), .Y(n27293) );
  NOR2X1 U30191 ( .A(n26083), .B(n27251), .Y(n21212) );
  INVX1 U30192 ( .A(reg_file[3916]), .Y(n27251) );
  NOR2X1 U30193 ( .A(n26083), .B(n27209), .Y(n21211) );
  INVX1 U30194 ( .A(reg_file[3917]), .Y(n27209) );
  NOR2X1 U30195 ( .A(n26083), .B(n27167), .Y(n21210) );
  INVX1 U30196 ( .A(reg_file[3918]), .Y(n27167) );
  NOR2X1 U30197 ( .A(n26083), .B(n27125), .Y(n21209) );
  INVX1 U30198 ( .A(reg_file[3919]), .Y(n27125) );
  NOR2X1 U30199 ( .A(n26083), .B(n27041), .Y(n21208) );
  INVX1 U30200 ( .A(reg_file[3920]), .Y(n27041) );
  NOR2X1 U30201 ( .A(n26083), .B(n26999), .Y(n21207) );
  INVX1 U30202 ( .A(reg_file[3921]), .Y(n26999) );
  NOR2X1 U30203 ( .A(n26084), .B(n26957), .Y(n21206) );
  INVX1 U30204 ( .A(reg_file[3922]), .Y(n26957) );
  NOR2X1 U30205 ( .A(n26084), .B(n26915), .Y(n21205) );
  INVX1 U30206 ( .A(reg_file[3923]), .Y(n26915) );
  NOR2X1 U30207 ( .A(n26084), .B(n26873), .Y(n21204) );
  INVX1 U30208 ( .A(reg_file[3924]), .Y(n26873) );
  NOR2X1 U30209 ( .A(n26084), .B(n26831), .Y(n21203) );
  INVX1 U30210 ( .A(reg_file[3925]), .Y(n26831) );
  NOR2X1 U30211 ( .A(n26084), .B(n26789), .Y(n21202) );
  INVX1 U30212 ( .A(reg_file[3926]), .Y(n26789) );
  NOR2X1 U30213 ( .A(n26084), .B(n26747), .Y(n21201) );
  INVX1 U30214 ( .A(reg_file[3927]), .Y(n26747) );
  NOR2X1 U30215 ( .A(n26084), .B(n26705), .Y(n21200) );
  INVX1 U30216 ( .A(reg_file[3928]), .Y(n26705) );
  NOR2X1 U30217 ( .A(n26084), .B(n26663), .Y(n21199) );
  INVX1 U30218 ( .A(reg_file[3929]), .Y(n26663) );
  NOR2X1 U30219 ( .A(n26084), .B(n26579), .Y(n21198) );
  INVX1 U30220 ( .A(reg_file[3930]), .Y(n26579) );
  NOR2X1 U30221 ( .A(n26084), .B(n26537), .Y(n21197) );
  INVX1 U30222 ( .A(reg_file[3931]), .Y(n26537) );
  NOR2X1 U30223 ( .A(n26084), .B(n26495), .Y(n21196) );
  INVX1 U30224 ( .A(reg_file[3932]), .Y(n26495) );
  NOR2X1 U30225 ( .A(n26084), .B(n26453), .Y(n21195) );
  INVX1 U30226 ( .A(reg_file[3933]), .Y(n26453) );
  NOR2X1 U30227 ( .A(n26084), .B(n26411), .Y(n21194) );
  INVX1 U30228 ( .A(reg_file[3934]), .Y(n26411) );
  NOR2X1 U30229 ( .A(n26084), .B(n26369), .Y(n21193) );
  INVX1 U30230 ( .A(reg_file[3935]), .Y(n26369) );
  NOR2X1 U30231 ( .A(n26084), .B(n26327), .Y(n21192) );
  INVX1 U30232 ( .A(reg_file[3936]), .Y(n26327) );
  NOR2X1 U30233 ( .A(n26084), .B(n26285), .Y(n21191) );
  INVX1 U30234 ( .A(reg_file[3937]), .Y(n26285) );
  NOR2X1 U30235 ( .A(n26084), .B(n26243), .Y(n21190) );
  INVX1 U30236 ( .A(reg_file[3938]), .Y(n26243) );
  NOR2X1 U30237 ( .A(n26085), .B(n26201), .Y(n21189) );
  INVX1 U30238 ( .A(reg_file[3939]), .Y(n26201) );
  NOR2X1 U30239 ( .A(n26085), .B(n31451), .Y(n21188) );
  INVX1 U30240 ( .A(reg_file[3940]), .Y(n31451) );
  NOR2X1 U30241 ( .A(n26085), .B(n31409), .Y(n21187) );
  INVX1 U30242 ( .A(reg_file[3941]), .Y(n31409) );
  NOR2X1 U30243 ( .A(n26085), .B(n31367), .Y(n21186) );
  INVX1 U30244 ( .A(reg_file[3942]), .Y(n31367) );
  NOR2X1 U30245 ( .A(n26085), .B(n31325), .Y(n21185) );
  INVX1 U30246 ( .A(reg_file[3943]), .Y(n31325) );
  NOR2X1 U30247 ( .A(n26085), .B(n31283), .Y(n21184) );
  INVX1 U30248 ( .A(reg_file[3944]), .Y(n31283) );
  NOR2X1 U30249 ( .A(n26085), .B(n31241), .Y(n21183) );
  INVX1 U30250 ( .A(reg_file[3945]), .Y(n31241) );
  NOR2X1 U30251 ( .A(n26085), .B(n31199), .Y(n21182) );
  INVX1 U30252 ( .A(reg_file[3946]), .Y(n31199) );
  NOR2X1 U30253 ( .A(n26085), .B(n31157), .Y(n21181) );
  INVX1 U30254 ( .A(reg_file[3947]), .Y(n31157) );
  NOR2X1 U30255 ( .A(n26085), .B(n31115), .Y(n21180) );
  INVX1 U30256 ( .A(reg_file[3948]), .Y(n31115) );
  NOR2X1 U30257 ( .A(n26085), .B(n31073), .Y(n21179) );
  INVX1 U30258 ( .A(reg_file[3949]), .Y(n31073) );
  NOR2X1 U30259 ( .A(n26085), .B(n30989), .Y(n21178) );
  INVX1 U30260 ( .A(reg_file[3950]), .Y(n30989) );
  NOR2X1 U30261 ( .A(n26085), .B(n30947), .Y(n21177) );
  INVX1 U30262 ( .A(reg_file[3951]), .Y(n30947) );
  NOR2X1 U30263 ( .A(n26085), .B(n30905), .Y(n21176) );
  INVX1 U30264 ( .A(reg_file[3952]), .Y(n30905) );
  NOR2X1 U30265 ( .A(n26085), .B(n30863), .Y(n21175) );
  INVX1 U30266 ( .A(reg_file[3953]), .Y(n30863) );
  NOR2X1 U30267 ( .A(n26085), .B(n30821), .Y(n21174) );
  INVX1 U30268 ( .A(reg_file[3954]), .Y(n30821) );
  NOR2X1 U30269 ( .A(n26085), .B(n30779), .Y(n21173) );
  INVX1 U30270 ( .A(reg_file[3955]), .Y(n30779) );
  NOR2X1 U30271 ( .A(n26086), .B(n30737), .Y(n21172) );
  INVX1 U30272 ( .A(reg_file[3956]), .Y(n30737) );
  NOR2X1 U30273 ( .A(n26086), .B(n30695), .Y(n21171) );
  INVX1 U30274 ( .A(reg_file[3957]), .Y(n30695) );
  NOR2X1 U30275 ( .A(n26086), .B(n30653), .Y(n21170) );
  INVX1 U30276 ( .A(reg_file[3958]), .Y(n30653) );
  NOR2X1 U30277 ( .A(n26086), .B(n30611), .Y(n21169) );
  INVX1 U30278 ( .A(reg_file[3959]), .Y(n30611) );
  NOR2X1 U30279 ( .A(n26086), .B(n30527), .Y(n21168) );
  INVX1 U30280 ( .A(reg_file[3960]), .Y(n30527) );
  NOR2X1 U30281 ( .A(n26086), .B(n30485), .Y(n21167) );
  INVX1 U30282 ( .A(reg_file[3961]), .Y(n30485) );
  NOR2X1 U30283 ( .A(n26086), .B(n30443), .Y(n21166) );
  INVX1 U30284 ( .A(reg_file[3962]), .Y(n30443) );
  NOR2X1 U30285 ( .A(n26086), .B(n30401), .Y(n21165) );
  INVX1 U30286 ( .A(reg_file[3963]), .Y(n30401) );
  NOR2X1 U30287 ( .A(n26086), .B(n30359), .Y(n21164) );
  INVX1 U30288 ( .A(reg_file[3964]), .Y(n30359) );
  NOR2X1 U30289 ( .A(n26086), .B(n30317), .Y(n21163) );
  INVX1 U30290 ( .A(reg_file[3965]), .Y(n30317) );
  NOR2X1 U30291 ( .A(n26086), .B(n30275), .Y(n21162) );
  INVX1 U30292 ( .A(reg_file[3966]), .Y(n30275) );
  NOR2X1 U30293 ( .A(n26086), .B(n30233), .Y(n21161) );
  INVX1 U30294 ( .A(reg_file[3967]), .Y(n30233) );
  NOR2X1 U30295 ( .A(n36623), .B(n35317), .Y(n37017) );
  NAND3X1 U30296 ( .A(wraddr[3]), .B(n35320), .C(wraddr[4]), .Y(n36623) );
  INVX1 U30297 ( .A(wraddr[0]), .Y(n35320) );
  MUX2X1 U30298 ( .B(n31511), .A(n25129), .S(n26087), .Y(n21160) );
  NOR2X1 U30299 ( .A(n37019), .B(n37020), .Y(n34913) );
  NAND3X1 U30300 ( .A(n37021), .B(n37022), .C(n37023), .Y(n37020) );
  AND2X1 U30301 ( .A(n37024), .B(n37025), .Y(n37023) );
  AOI22X1 U30302 ( .A(wrdata[55]), .B(n37026), .C(wrdata[47]), .D(n37027), .Y(
        n37025) );
  AOI22X1 U30303 ( .A(wrdata[127]), .B(wrbyteen[15]), .C(wrdata[7]), .D(n37028), .Y(n37024) );
  AOI22X1 U30304 ( .A(wrdata[119]), .B(n37029), .C(wrdata[63]), .D(n37030), 
        .Y(n37022) );
  AOI22X1 U30305 ( .A(wrdata[39]), .B(n37031), .C(wrdata[31]), .D(n37032), .Y(
        n37021) );
  NAND3X1 U30306 ( .A(n37033), .B(n37034), .C(n37035), .Y(n37019) );
  AND2X1 U30307 ( .A(n37036), .B(n37037), .Y(n37035) );
  AOI22X1 U30308 ( .A(wrdata[111]), .B(n37038), .C(wrdata[87]), .D(n37039), 
        .Y(n37037) );
  AOI22X1 U30309 ( .A(wrdata[103]), .B(n37040), .C(wrdata[95]), .D(n37041), 
        .Y(n37036) );
  AOI22X1 U30310 ( .A(wrdata[79]), .B(n37042), .C(wrdata[71]), .D(n37043), .Y(
        n37034) );
  AOI22X1 U30311 ( .A(wrdata[23]), .B(n37044), .C(wrdata[15]), .D(n37045), .Y(
        n37033) );
  INVX1 U30312 ( .A(reg_file[3968]), .Y(n31511) );
  MUX2X1 U30313 ( .B(n29856), .A(n25130), .S(n26087), .Y(n21159) );
  NOR2X1 U30314 ( .A(n37046), .B(n37047), .Y(n34915) );
  NAND3X1 U30315 ( .A(n37048), .B(n37049), .C(n37050), .Y(n37047) );
  AND2X1 U30316 ( .A(n37051), .B(n37052), .Y(n37050) );
  AOI22X1 U30317 ( .A(wrdata[54]), .B(n37026), .C(wrdata[46]), .D(n37027), .Y(
        n37052) );
  AOI22X1 U30318 ( .A(wrdata[126]), .B(wrbyteen[15]), .C(wrdata[6]), .D(n37028), .Y(n37051) );
  AOI22X1 U30319 ( .A(wrdata[118]), .B(n37029), .C(wrdata[62]), .D(n37030), 
        .Y(n37049) );
  AOI22X1 U30320 ( .A(wrdata[38]), .B(n37031), .C(wrdata[30]), .D(n37032), .Y(
        n37048) );
  NAND3X1 U30321 ( .A(n37053), .B(n37054), .C(n37055), .Y(n37046) );
  AND2X1 U30322 ( .A(n37056), .B(n37057), .Y(n37055) );
  AOI22X1 U30323 ( .A(wrdata[110]), .B(n37038), .C(wrdata[86]), .D(n37039), 
        .Y(n37057) );
  AOI22X1 U30324 ( .A(wrdata[102]), .B(n37040), .C(wrdata[94]), .D(n37041), 
        .Y(n37056) );
  AOI22X1 U30325 ( .A(wrdata[78]), .B(n37042), .C(wrdata[70]), .D(n37043), .Y(
        n37054) );
  AOI22X1 U30326 ( .A(wrdata[22]), .B(n37044), .C(wrdata[14]), .D(n37045), .Y(
        n37053) );
  INVX1 U30327 ( .A(reg_file[3969]), .Y(n29856) );
  MUX2X1 U30328 ( .B(n29394), .A(n25131), .S(n26087), .Y(n21158) );
  NOR2X1 U30329 ( .A(n37058), .B(n37059), .Y(n34916) );
  NAND3X1 U30330 ( .A(n37060), .B(n37061), .C(n37062), .Y(n37059) );
  AND2X1 U30331 ( .A(n37063), .B(n37064), .Y(n37062) );
  AOI22X1 U30332 ( .A(wrdata[53]), .B(n37026), .C(wrdata[45]), .D(n37027), .Y(
        n37064) );
  AOI22X1 U30333 ( .A(wrdata[125]), .B(wrbyteen[15]), .C(wrdata[5]), .D(n37028), .Y(n37063) );
  AOI22X1 U30334 ( .A(wrdata[117]), .B(n37029), .C(wrdata[61]), .D(n37030), 
        .Y(n37061) );
  AOI22X1 U30335 ( .A(wrdata[37]), .B(n37031), .C(wrdata[29]), .D(n37032), .Y(
        n37060) );
  NAND3X1 U30336 ( .A(n37065), .B(n37066), .C(n37067), .Y(n37058) );
  AND2X1 U30337 ( .A(n37068), .B(n37069), .Y(n37067) );
  AOI22X1 U30338 ( .A(wrdata[109]), .B(n37038), .C(wrdata[85]), .D(n37039), 
        .Y(n37069) );
  AOI22X1 U30339 ( .A(wrdata[101]), .B(n37040), .C(wrdata[93]), .D(n37041), 
        .Y(n37068) );
  AOI22X1 U30340 ( .A(wrdata[77]), .B(n37042), .C(wrdata[69]), .D(n37043), .Y(
        n37066) );
  AOI22X1 U30341 ( .A(wrdata[21]), .B(n37044), .C(wrdata[13]), .D(n37045), .Y(
        n37065) );
  INVX1 U30342 ( .A(reg_file[3970]), .Y(n29394) );
  MUX2X1 U30343 ( .B(n28932), .A(n25132), .S(n26087), .Y(n21157) );
  NOR2X1 U30344 ( .A(n37070), .B(n37071), .Y(n34917) );
  NAND3X1 U30345 ( .A(n37072), .B(n37073), .C(n37074), .Y(n37071) );
  AND2X1 U30346 ( .A(n37075), .B(n37076), .Y(n37074) );
  AOI22X1 U30347 ( .A(wrdata[52]), .B(n37026), .C(wrdata[44]), .D(n37027), .Y(
        n37076) );
  AOI22X1 U30348 ( .A(wrdata[124]), .B(wrbyteen[15]), .C(wrdata[4]), .D(n37028), .Y(n37075) );
  AOI22X1 U30349 ( .A(wrdata[116]), .B(n37029), .C(wrdata[60]), .D(n37030), 
        .Y(n37073) );
  AOI22X1 U30350 ( .A(wrdata[36]), .B(n37031), .C(wrdata[28]), .D(n37032), .Y(
        n37072) );
  NAND3X1 U30351 ( .A(n37077), .B(n37078), .C(n37079), .Y(n37070) );
  AND2X1 U30352 ( .A(n37080), .B(n37081), .Y(n37079) );
  AOI22X1 U30353 ( .A(wrdata[108]), .B(n37038), .C(wrdata[84]), .D(n37039), 
        .Y(n37081) );
  AOI22X1 U30354 ( .A(wrdata[100]), .B(n37040), .C(wrdata[92]), .D(n37041), 
        .Y(n37080) );
  AOI22X1 U30355 ( .A(wrdata[76]), .B(n37042), .C(wrdata[68]), .D(n37043), .Y(
        n37078) );
  AOI22X1 U30356 ( .A(wrdata[20]), .B(n37044), .C(wrdata[12]), .D(n37045), .Y(
        n37077) );
  INVX1 U30357 ( .A(reg_file[3971]), .Y(n28932) );
  MUX2X1 U30358 ( .B(n28470), .A(n25133), .S(n26087), .Y(n21156) );
  NOR2X1 U30359 ( .A(n37082), .B(n37083), .Y(n34918) );
  NAND3X1 U30360 ( .A(n37084), .B(n37085), .C(n37086), .Y(n37083) );
  AND2X1 U30361 ( .A(n37087), .B(n37088), .Y(n37086) );
  AOI22X1 U30362 ( .A(wrdata[51]), .B(n37026), .C(wrdata[43]), .D(n37027), .Y(
        n37088) );
  AOI22X1 U30363 ( .A(wrdata[123]), .B(wrbyteen[15]), .C(wrdata[3]), .D(n37028), .Y(n37087) );
  AOI22X1 U30364 ( .A(wrdata[115]), .B(n37029), .C(wrdata[59]), .D(n37030), 
        .Y(n37085) );
  AOI22X1 U30365 ( .A(wrdata[35]), .B(n37031), .C(wrdata[27]), .D(n37032), .Y(
        n37084) );
  NAND3X1 U30366 ( .A(n37089), .B(n37090), .C(n37091), .Y(n37082) );
  AND2X1 U30367 ( .A(n37092), .B(n37093), .Y(n37091) );
  AOI22X1 U30368 ( .A(wrdata[107]), .B(n37038), .C(wrdata[83]), .D(n37039), 
        .Y(n37093) );
  AOI22X1 U30369 ( .A(wrdata[99]), .B(n37040), .C(wrdata[91]), .D(n37041), .Y(
        n37092) );
  AOI22X1 U30370 ( .A(wrdata[75]), .B(n37042), .C(wrdata[67]), .D(n37043), .Y(
        n37090) );
  AOI22X1 U30371 ( .A(wrdata[19]), .B(n37044), .C(wrdata[11]), .D(n37045), .Y(
        n37089) );
  INVX1 U30372 ( .A(reg_file[3972]), .Y(n28470) );
  MUX2X1 U30373 ( .B(n28008), .A(n25134), .S(n26087), .Y(n21155) );
  NOR2X1 U30374 ( .A(n37094), .B(n37095), .Y(n34919) );
  NAND3X1 U30375 ( .A(n37096), .B(n37097), .C(n37098), .Y(n37095) );
  AND2X1 U30376 ( .A(n37099), .B(n37100), .Y(n37098) );
  AOI22X1 U30377 ( .A(wrdata[50]), .B(n37026), .C(wrdata[42]), .D(n37027), .Y(
        n37100) );
  AOI22X1 U30378 ( .A(wrdata[122]), .B(wrbyteen[15]), .C(wrdata[2]), .D(n37028), .Y(n37099) );
  AOI22X1 U30379 ( .A(wrdata[114]), .B(n37029), .C(wrdata[58]), .D(n37030), 
        .Y(n37097) );
  AOI22X1 U30380 ( .A(wrdata[34]), .B(n37031), .C(wrdata[26]), .D(n37032), .Y(
        n37096) );
  NAND3X1 U30381 ( .A(n37101), .B(n37102), .C(n37103), .Y(n37094) );
  AND2X1 U30382 ( .A(n37104), .B(n37105), .Y(n37103) );
  AOI22X1 U30383 ( .A(wrdata[106]), .B(n37038), .C(wrdata[82]), .D(n37039), 
        .Y(n37105) );
  AOI22X1 U30384 ( .A(wrdata[98]), .B(n37040), .C(wrdata[90]), .D(n37041), .Y(
        n37104) );
  AOI22X1 U30385 ( .A(wrdata[74]), .B(n37042), .C(wrdata[66]), .D(n37043), .Y(
        n37102) );
  AOI22X1 U30386 ( .A(wrdata[18]), .B(n37044), .C(wrdata[10]), .D(n37045), .Y(
        n37101) );
  INVX1 U30387 ( .A(reg_file[3973]), .Y(n28008) );
  MUX2X1 U30388 ( .B(n27546), .A(n25135), .S(n26087), .Y(n21154) );
  NOR2X1 U30389 ( .A(n37106), .B(n37107), .Y(n34920) );
  NAND3X1 U30390 ( .A(n37108), .B(n37109), .C(n37110), .Y(n37107) );
  AND2X1 U30391 ( .A(n37111), .B(n37112), .Y(n37110) );
  AOI22X1 U30392 ( .A(wrdata[49]), .B(n37026), .C(wrdata[41]), .D(n37027), .Y(
        n37112) );
  AOI22X1 U30393 ( .A(wrdata[121]), .B(wrbyteen[15]), .C(wrdata[1]), .D(n37028), .Y(n37111) );
  AOI22X1 U30394 ( .A(wrdata[113]), .B(n37029), .C(wrdata[57]), .D(n37030), 
        .Y(n37109) );
  AOI22X1 U30395 ( .A(wrdata[33]), .B(n37031), .C(wrdata[25]), .D(n37032), .Y(
        n37108) );
  NAND3X1 U30396 ( .A(n37113), .B(n37114), .C(n37115), .Y(n37106) );
  AND2X1 U30397 ( .A(n37116), .B(n37117), .Y(n37115) );
  AOI22X1 U30398 ( .A(wrdata[105]), .B(n37038), .C(wrdata[81]), .D(n37039), 
        .Y(n37117) );
  AOI22X1 U30399 ( .A(wrdata[97]), .B(n37040), .C(wrdata[89]), .D(n37041), .Y(
        n37116) );
  AOI22X1 U30400 ( .A(wrdata[73]), .B(n37042), .C(wrdata[65]), .D(n37043), .Y(
        n37114) );
  AOI22X1 U30401 ( .A(wrdata[17]), .B(n37044), .C(wrdata[9]), .D(n37045), .Y(
        n37113) );
  INVX1 U30402 ( .A(reg_file[3974]), .Y(n27546) );
  MUX2X1 U30403 ( .B(n27084), .A(n25136), .S(n26087), .Y(n21153) );
  NOR2X1 U30404 ( .A(n37118), .B(n37119), .Y(n34921) );
  NAND3X1 U30405 ( .A(n37120), .B(n37121), .C(n37122), .Y(n37119) );
  AND2X1 U30406 ( .A(n37123), .B(n37124), .Y(n37122) );
  AOI22X1 U30407 ( .A(wrdata[48]), .B(n37026), .C(wrdata[40]), .D(n37027), .Y(
        n37124) );
  NOR2X1 U30408 ( .A(n37125), .B(wrbyteen[6]), .Y(n37027) );
  NOR2X1 U30409 ( .A(n37126), .B(wrbyteen[7]), .Y(n37026) );
  AOI22X1 U30410 ( .A(wrdata[120]), .B(wrbyteen[15]), .C(wrdata[0]), .D(n37028), .Y(n37123) );
  AOI22X1 U30411 ( .A(wrdata[112]), .B(n37029), .C(wrdata[56]), .D(n37030), 
        .Y(n37121) );
  NOR2X1 U30412 ( .A(n37127), .B(wrbyteen[8]), .Y(n37030) );
  AND2X1 U30413 ( .A(wrbyteen[14]), .B(n37128), .Y(n37029) );
  AOI22X1 U30414 ( .A(wrdata[32]), .B(n37031), .C(wrdata[24]), .D(n37032), .Y(
        n37120) );
  NOR2X1 U30415 ( .A(n37129), .B(wrbyteen[4]), .Y(n37032) );
  NOR2X1 U30416 ( .A(n37130), .B(wrbyteen[5]), .Y(n37031) );
  NAND3X1 U30417 ( .A(n37131), .B(n37132), .C(n37133), .Y(n37118) );
  AND2X1 U30418 ( .A(n37134), .B(n37135), .Y(n37133) );
  AOI22X1 U30419 ( .A(wrdata[104]), .B(n37038), .C(wrdata[80]), .D(n37039), 
        .Y(n37135) );
  NOR2X1 U30420 ( .A(n37136), .B(wrbyteen[11]), .Y(n37039) );
  NOR2X1 U30421 ( .A(n37137), .B(wrbyteen[14]), .Y(n37038) );
  AOI22X1 U30422 ( .A(wrdata[96]), .B(n37040), .C(wrdata[88]), .D(n37041), .Y(
        n37134) );
  AND2X1 U30423 ( .A(wrbyteen[11]), .B(n37138), .Y(n37041) );
  NOR2X1 U30424 ( .A(n37138), .B(wrbyteen[13]), .Y(n37040) );
  AOI22X1 U30425 ( .A(wrdata[72]), .B(n37042), .C(wrdata[64]), .D(n37043), .Y(
        n37132) );
  AND2X1 U30426 ( .A(wrbyteen[8]), .B(n37139), .Y(n37043) );
  NOR2X1 U30427 ( .A(n37139), .B(wrbyteen[10]), .Y(n37042) );
  AOI22X1 U30428 ( .A(wrdata[16]), .B(n37044), .C(wrdata[8]), .D(n37045), .Y(
        n37131) );
  NOR2X1 U30429 ( .A(n37028), .B(wrbyteen[2]), .Y(n37045) );
  AND2X1 U30430 ( .A(wrbyteen[2]), .B(n37129), .Y(n37044) );
  INVX1 U30431 ( .A(reg_file[3975]), .Y(n27084) );
  NOR2X1 U30432 ( .A(n26087), .B(n26622), .Y(n21152) );
  INVX1 U30433 ( .A(reg_file[3976]), .Y(n26622) );
  NOR2X1 U30434 ( .A(n26087), .B(n26148), .Y(n21151) );
  INVX1 U30435 ( .A(reg_file[3977]), .Y(n26148) );
  NOR2X1 U30436 ( .A(n26087), .B(n31032), .Y(n21150) );
  INVX1 U30437 ( .A(reg_file[3978]), .Y(n31032) );
  NOR2X1 U30438 ( .A(n26087), .B(n30570), .Y(n21149) );
  INVX1 U30439 ( .A(reg_file[3979]), .Y(n30570) );
  NOR2X1 U30440 ( .A(n26087), .B(n30192), .Y(n21148) );
  INVX1 U30441 ( .A(reg_file[3980]), .Y(n30192) );
  NOR2X1 U30442 ( .A(n26087), .B(n30150), .Y(n21147) );
  INVX1 U30443 ( .A(reg_file[3981]), .Y(n30150) );
  NOR2X1 U30444 ( .A(n26088), .B(n30108), .Y(n21146) );
  INVX1 U30445 ( .A(reg_file[3982]), .Y(n30108) );
  NOR2X1 U30446 ( .A(n26088), .B(n30066), .Y(n21145) );
  INVX1 U30447 ( .A(reg_file[3983]), .Y(n30066) );
  NOR2X1 U30448 ( .A(n26088), .B(n30024), .Y(n21144) );
  INVX1 U30449 ( .A(reg_file[3984]), .Y(n30024) );
  NOR2X1 U30450 ( .A(n26088), .B(n29982), .Y(n21143) );
  INVX1 U30451 ( .A(reg_file[3985]), .Y(n29982) );
  NOR2X1 U30452 ( .A(n26088), .B(n29940), .Y(n21142) );
  INVX1 U30453 ( .A(reg_file[3986]), .Y(n29940) );
  NOR2X1 U30454 ( .A(n26088), .B(n29898), .Y(n21141) );
  INVX1 U30455 ( .A(reg_file[3987]), .Y(n29898) );
  NOR2X1 U30456 ( .A(n26088), .B(n29814), .Y(n21140) );
  INVX1 U30457 ( .A(reg_file[3988]), .Y(n29814) );
  NOR2X1 U30458 ( .A(n26088), .B(n29772), .Y(n21139) );
  INVX1 U30459 ( .A(reg_file[3989]), .Y(n29772) );
  NOR2X1 U30460 ( .A(n26088), .B(n29730), .Y(n21138) );
  INVX1 U30461 ( .A(reg_file[3990]), .Y(n29730) );
  NOR2X1 U30462 ( .A(n26088), .B(n29688), .Y(n21137) );
  INVX1 U30463 ( .A(reg_file[3991]), .Y(n29688) );
  NOR2X1 U30464 ( .A(n26088), .B(n29646), .Y(n21136) );
  INVX1 U30465 ( .A(reg_file[3992]), .Y(n29646) );
  NOR2X1 U30466 ( .A(n26088), .B(n29604), .Y(n21135) );
  INVX1 U30467 ( .A(reg_file[3993]), .Y(n29604) );
  NOR2X1 U30468 ( .A(n26088), .B(n29562), .Y(n21134) );
  INVX1 U30469 ( .A(reg_file[3994]), .Y(n29562) );
  NOR2X1 U30470 ( .A(n26088), .B(n29520), .Y(n21133) );
  INVX1 U30471 ( .A(reg_file[3995]), .Y(n29520) );
  NOR2X1 U30472 ( .A(n26088), .B(n29478), .Y(n21132) );
  INVX1 U30473 ( .A(reg_file[3996]), .Y(n29478) );
  NOR2X1 U30474 ( .A(n26088), .B(n29436), .Y(n21131) );
  INVX1 U30475 ( .A(reg_file[3997]), .Y(n29436) );
  NOR2X1 U30476 ( .A(n26088), .B(n29352), .Y(n21130) );
  INVX1 U30477 ( .A(reg_file[3998]), .Y(n29352) );
  NOR2X1 U30478 ( .A(n26089), .B(n29310), .Y(n21129) );
  INVX1 U30479 ( .A(reg_file[3999]), .Y(n29310) );
  NOR2X1 U30480 ( .A(n26089), .B(n29268), .Y(n21128) );
  INVX1 U30481 ( .A(reg_file[4000]), .Y(n29268) );
  NOR2X1 U30482 ( .A(n26089), .B(n29226), .Y(n21127) );
  INVX1 U30483 ( .A(reg_file[4001]), .Y(n29226) );
  NOR2X1 U30484 ( .A(n26089), .B(n29184), .Y(n21126) );
  INVX1 U30485 ( .A(reg_file[4002]), .Y(n29184) );
  NOR2X1 U30486 ( .A(n26089), .B(n29142), .Y(n21125) );
  INVX1 U30487 ( .A(reg_file[4003]), .Y(n29142) );
  NOR2X1 U30488 ( .A(n26089), .B(n29100), .Y(n21124) );
  INVX1 U30489 ( .A(reg_file[4004]), .Y(n29100) );
  NOR2X1 U30490 ( .A(n26089), .B(n29058), .Y(n21123) );
  INVX1 U30491 ( .A(reg_file[4005]), .Y(n29058) );
  NOR2X1 U30492 ( .A(n26089), .B(n29016), .Y(n21122) );
  INVX1 U30493 ( .A(reg_file[4006]), .Y(n29016) );
  NOR2X1 U30494 ( .A(n26089), .B(n28974), .Y(n21121) );
  INVX1 U30495 ( .A(reg_file[4007]), .Y(n28974) );
  NOR2X1 U30496 ( .A(n26089), .B(n28890), .Y(n21120) );
  INVX1 U30497 ( .A(reg_file[4008]), .Y(n28890) );
  NOR2X1 U30498 ( .A(n26089), .B(n28848), .Y(n21119) );
  INVX1 U30499 ( .A(reg_file[4009]), .Y(n28848) );
  NOR2X1 U30500 ( .A(n26089), .B(n28806), .Y(n21118) );
  INVX1 U30501 ( .A(reg_file[4010]), .Y(n28806) );
  NOR2X1 U30502 ( .A(n26089), .B(n28764), .Y(n21117) );
  INVX1 U30503 ( .A(reg_file[4011]), .Y(n28764) );
  NOR2X1 U30504 ( .A(n26089), .B(n28722), .Y(n21116) );
  INVX1 U30505 ( .A(reg_file[4012]), .Y(n28722) );
  NOR2X1 U30506 ( .A(n26089), .B(n28680), .Y(n21115) );
  INVX1 U30507 ( .A(reg_file[4013]), .Y(n28680) );
  NOR2X1 U30508 ( .A(n26089), .B(n28638), .Y(n21114) );
  INVX1 U30509 ( .A(reg_file[4014]), .Y(n28638) );
  NOR2X1 U30510 ( .A(n26089), .B(n28596), .Y(n21113) );
  INVX1 U30511 ( .A(reg_file[4015]), .Y(n28596) );
  NOR2X1 U30512 ( .A(n26090), .B(n28554), .Y(n21112) );
  INVX1 U30513 ( .A(reg_file[4016]), .Y(n28554) );
  NOR2X1 U30514 ( .A(n26090), .B(n28512), .Y(n21111) );
  INVX1 U30515 ( .A(reg_file[4017]), .Y(n28512) );
  NOR2X1 U30516 ( .A(n26090), .B(n28428), .Y(n21110) );
  INVX1 U30517 ( .A(reg_file[4018]), .Y(n28428) );
  NOR2X1 U30518 ( .A(n26090), .B(n28386), .Y(n21109) );
  INVX1 U30519 ( .A(reg_file[4019]), .Y(n28386) );
  NOR2X1 U30520 ( .A(n26090), .B(n28344), .Y(n21108) );
  INVX1 U30521 ( .A(reg_file[4020]), .Y(n28344) );
  NOR2X1 U30522 ( .A(n26090), .B(n28302), .Y(n21107) );
  INVX1 U30523 ( .A(reg_file[4021]), .Y(n28302) );
  NOR2X1 U30524 ( .A(n26090), .B(n28260), .Y(n21106) );
  INVX1 U30525 ( .A(reg_file[4022]), .Y(n28260) );
  NOR2X1 U30526 ( .A(n26090), .B(n28218), .Y(n21105) );
  INVX1 U30527 ( .A(reg_file[4023]), .Y(n28218) );
  NOR2X1 U30528 ( .A(n26090), .B(n28176), .Y(n21104) );
  INVX1 U30529 ( .A(reg_file[4024]), .Y(n28176) );
  NOR2X1 U30530 ( .A(n26090), .B(n28134), .Y(n21103) );
  INVX1 U30531 ( .A(reg_file[4025]), .Y(n28134) );
  NOR2X1 U30532 ( .A(n26090), .B(n28092), .Y(n21102) );
  INVX1 U30533 ( .A(reg_file[4026]), .Y(n28092) );
  NOR2X1 U30534 ( .A(n26090), .B(n28050), .Y(n21101) );
  INVX1 U30535 ( .A(reg_file[4027]), .Y(n28050) );
  NOR2X1 U30536 ( .A(n26090), .B(n27966), .Y(n21100) );
  INVX1 U30537 ( .A(reg_file[4028]), .Y(n27966) );
  NOR2X1 U30538 ( .A(n26090), .B(n27924), .Y(n21099) );
  INVX1 U30539 ( .A(reg_file[4029]), .Y(n27924) );
  NOR2X1 U30540 ( .A(n26090), .B(n27882), .Y(n21098) );
  INVX1 U30541 ( .A(reg_file[4030]), .Y(n27882) );
  NOR2X1 U30542 ( .A(n26090), .B(n27840), .Y(n21097) );
  INVX1 U30543 ( .A(reg_file[4031]), .Y(n27840) );
  NOR2X1 U30544 ( .A(n26090), .B(n27798), .Y(n21096) );
  INVX1 U30545 ( .A(reg_file[4032]), .Y(n27798) );
  NOR2X1 U30546 ( .A(n26091), .B(n27756), .Y(n21095) );
  INVX1 U30547 ( .A(reg_file[4033]), .Y(n27756) );
  NOR2X1 U30548 ( .A(n26091), .B(n27714), .Y(n21094) );
  INVX1 U30549 ( .A(reg_file[4034]), .Y(n27714) );
  NOR2X1 U30550 ( .A(n26091), .B(n27672), .Y(n21093) );
  INVX1 U30551 ( .A(reg_file[4035]), .Y(n27672) );
  NOR2X1 U30552 ( .A(n26091), .B(n27630), .Y(n21092) );
  INVX1 U30553 ( .A(reg_file[4036]), .Y(n27630) );
  NOR2X1 U30554 ( .A(n26091), .B(n27588), .Y(n21091) );
  INVX1 U30555 ( .A(reg_file[4037]), .Y(n27588) );
  NOR2X1 U30556 ( .A(n26091), .B(n27504), .Y(n21090) );
  INVX1 U30557 ( .A(reg_file[4038]), .Y(n27504) );
  NOR2X1 U30558 ( .A(n26091), .B(n27462), .Y(n21089) );
  INVX1 U30559 ( .A(reg_file[4039]), .Y(n27462) );
  NOR2X1 U30560 ( .A(n26091), .B(n27420), .Y(n21088) );
  INVX1 U30561 ( .A(reg_file[4040]), .Y(n27420) );
  NOR2X1 U30562 ( .A(n26091), .B(n27378), .Y(n21087) );
  INVX1 U30563 ( .A(reg_file[4041]), .Y(n27378) );
  NOR2X1 U30564 ( .A(n26091), .B(n27336), .Y(n21086) );
  INVX1 U30565 ( .A(reg_file[4042]), .Y(n27336) );
  NOR2X1 U30566 ( .A(n26091), .B(n27294), .Y(n21085) );
  INVX1 U30567 ( .A(reg_file[4043]), .Y(n27294) );
  NOR2X1 U30568 ( .A(n26091), .B(n27252), .Y(n21084) );
  INVX1 U30569 ( .A(reg_file[4044]), .Y(n27252) );
  NOR2X1 U30570 ( .A(n26091), .B(n27210), .Y(n21083) );
  INVX1 U30571 ( .A(reg_file[4045]), .Y(n27210) );
  NOR2X1 U30572 ( .A(n26091), .B(n27168), .Y(n21082) );
  INVX1 U30573 ( .A(reg_file[4046]), .Y(n27168) );
  NOR2X1 U30574 ( .A(n26091), .B(n27126), .Y(n21081) );
  INVX1 U30575 ( .A(reg_file[4047]), .Y(n27126) );
  NOR2X1 U30576 ( .A(n26091), .B(n27042), .Y(n21080) );
  INVX1 U30577 ( .A(reg_file[4048]), .Y(n27042) );
  NOR2X1 U30578 ( .A(n26091), .B(n27000), .Y(n21079) );
  INVX1 U30579 ( .A(reg_file[4049]), .Y(n27000) );
  NOR2X1 U30580 ( .A(n26092), .B(n26958), .Y(n21078) );
  INVX1 U30581 ( .A(reg_file[4050]), .Y(n26958) );
  NOR2X1 U30582 ( .A(n26092), .B(n26916), .Y(n21077) );
  INVX1 U30583 ( .A(reg_file[4051]), .Y(n26916) );
  NOR2X1 U30584 ( .A(n26092), .B(n26874), .Y(n21076) );
  INVX1 U30585 ( .A(reg_file[4052]), .Y(n26874) );
  NOR2X1 U30586 ( .A(n26092), .B(n26832), .Y(n21075) );
  INVX1 U30587 ( .A(reg_file[4053]), .Y(n26832) );
  NOR2X1 U30588 ( .A(n26092), .B(n26790), .Y(n21074) );
  INVX1 U30589 ( .A(reg_file[4054]), .Y(n26790) );
  NOR2X1 U30590 ( .A(n26092), .B(n26748), .Y(n21073) );
  INVX1 U30591 ( .A(reg_file[4055]), .Y(n26748) );
  NOR2X1 U30592 ( .A(n26092), .B(n26706), .Y(n21072) );
  INVX1 U30593 ( .A(reg_file[4056]), .Y(n26706) );
  NOR2X1 U30594 ( .A(n26092), .B(n26664), .Y(n21071) );
  INVX1 U30595 ( .A(reg_file[4057]), .Y(n26664) );
  NOR2X1 U30596 ( .A(n26092), .B(n26580), .Y(n21070) );
  INVX1 U30597 ( .A(reg_file[4058]), .Y(n26580) );
  NOR2X1 U30598 ( .A(n26092), .B(n26538), .Y(n21069) );
  INVX1 U30599 ( .A(reg_file[4059]), .Y(n26538) );
  NOR2X1 U30600 ( .A(n26092), .B(n26496), .Y(n21068) );
  INVX1 U30601 ( .A(reg_file[4060]), .Y(n26496) );
  NOR2X1 U30602 ( .A(n26092), .B(n26454), .Y(n21067) );
  INVX1 U30603 ( .A(reg_file[4061]), .Y(n26454) );
  NOR2X1 U30604 ( .A(n26092), .B(n26412), .Y(n21066) );
  INVX1 U30605 ( .A(reg_file[4062]), .Y(n26412) );
  NOR2X1 U30606 ( .A(n26092), .B(n26370), .Y(n21065) );
  INVX1 U30607 ( .A(reg_file[4063]), .Y(n26370) );
  NOR2X1 U30608 ( .A(n26092), .B(n26328), .Y(n21064) );
  INVX1 U30609 ( .A(reg_file[4064]), .Y(n26328) );
  NOR2X1 U30610 ( .A(n26092), .B(n26286), .Y(n21063) );
  INVX1 U30611 ( .A(reg_file[4065]), .Y(n26286) );
  NOR2X1 U30612 ( .A(n26092), .B(n26244), .Y(n21062) );
  INVX1 U30613 ( .A(reg_file[4066]), .Y(n26244) );
  NOR2X1 U30614 ( .A(n26093), .B(n26202), .Y(n21061) );
  INVX1 U30615 ( .A(reg_file[4067]), .Y(n26202) );
  NOR2X1 U30616 ( .A(n26093), .B(n31452), .Y(n21060) );
  INVX1 U30617 ( .A(reg_file[4068]), .Y(n31452) );
  NOR2X1 U30618 ( .A(n26093), .B(n31410), .Y(n21059) );
  INVX1 U30619 ( .A(reg_file[4069]), .Y(n31410) );
  NOR2X1 U30620 ( .A(n26093), .B(n31368), .Y(n21058) );
  INVX1 U30621 ( .A(reg_file[4070]), .Y(n31368) );
  NOR2X1 U30622 ( .A(n26093), .B(n31326), .Y(n21057) );
  INVX1 U30623 ( .A(reg_file[4071]), .Y(n31326) );
  NOR2X1 U30624 ( .A(n26093), .B(n31284), .Y(n21056) );
  INVX1 U30625 ( .A(reg_file[4072]), .Y(n31284) );
  NOR2X1 U30626 ( .A(n26093), .B(n31242), .Y(n21055) );
  INVX1 U30627 ( .A(reg_file[4073]), .Y(n31242) );
  NOR2X1 U30628 ( .A(n26093), .B(n31200), .Y(n21054) );
  INVX1 U30629 ( .A(reg_file[4074]), .Y(n31200) );
  NOR2X1 U30630 ( .A(n26093), .B(n31158), .Y(n21053) );
  INVX1 U30631 ( .A(reg_file[4075]), .Y(n31158) );
  NOR2X1 U30632 ( .A(n26093), .B(n31116), .Y(n21052) );
  INVX1 U30633 ( .A(reg_file[4076]), .Y(n31116) );
  NOR2X1 U30634 ( .A(n26093), .B(n31074), .Y(n21051) );
  INVX1 U30635 ( .A(reg_file[4077]), .Y(n31074) );
  NOR2X1 U30636 ( .A(n26093), .B(n30990), .Y(n21050) );
  INVX1 U30637 ( .A(reg_file[4078]), .Y(n30990) );
  NOR2X1 U30638 ( .A(n26093), .B(n30948), .Y(n21049) );
  INVX1 U30639 ( .A(reg_file[4079]), .Y(n30948) );
  NOR2X1 U30640 ( .A(n26093), .B(n30906), .Y(n21048) );
  INVX1 U30641 ( .A(reg_file[4080]), .Y(n30906) );
  NOR2X1 U30642 ( .A(n26093), .B(n30864), .Y(n21047) );
  INVX1 U30643 ( .A(reg_file[4081]), .Y(n30864) );
  NOR2X1 U30644 ( .A(n26093), .B(n30822), .Y(n21046) );
  INVX1 U30645 ( .A(reg_file[4082]), .Y(n30822) );
  NOR2X1 U30646 ( .A(n26093), .B(n30780), .Y(n21045) );
  INVX1 U30647 ( .A(reg_file[4083]), .Y(n30780) );
  NOR2X1 U30648 ( .A(n26094), .B(n30738), .Y(n21044) );
  INVX1 U30649 ( .A(reg_file[4084]), .Y(n30738) );
  NOR2X1 U30650 ( .A(n26094), .B(n30696), .Y(n21043) );
  INVX1 U30651 ( .A(reg_file[4085]), .Y(n30696) );
  NOR2X1 U30652 ( .A(n26094), .B(n30654), .Y(n21042) );
  INVX1 U30653 ( .A(reg_file[4086]), .Y(n30654) );
  NOR2X1 U30654 ( .A(n26094), .B(n30612), .Y(n21041) );
  INVX1 U30655 ( .A(reg_file[4087]), .Y(n30612) );
  NOR2X1 U30656 ( .A(n26094), .B(n30528), .Y(n21040) );
  INVX1 U30657 ( .A(reg_file[4088]), .Y(n30528) );
  NOR2X1 U30658 ( .A(n26094), .B(n30486), .Y(n21039) );
  INVX1 U30659 ( .A(reg_file[4089]), .Y(n30486) );
  NOR2X1 U30660 ( .A(n26094), .B(n30444), .Y(n21038) );
  INVX1 U30661 ( .A(reg_file[4090]), .Y(n30444) );
  NOR2X1 U30662 ( .A(n26094), .B(n30402), .Y(n21037) );
  INVX1 U30663 ( .A(reg_file[4091]), .Y(n30402) );
  NOR2X1 U30664 ( .A(n26094), .B(n30360), .Y(n21036) );
  INVX1 U30665 ( .A(reg_file[4092]), .Y(n30360) );
  NOR2X1 U30666 ( .A(n26094), .B(n30318), .Y(n21035) );
  INVX1 U30667 ( .A(reg_file[4093]), .Y(n30318) );
  NOR2X1 U30668 ( .A(n26094), .B(n30276), .Y(n21034) );
  INVX1 U30669 ( .A(reg_file[4094]), .Y(n30276) );
  NOR2X1 U30670 ( .A(n26094), .B(n30234), .Y(n21033) );
  INVX1 U30671 ( .A(reg_file[4095]), .Y(n30234) );
  NOR2X1 U30672 ( .A(n36753), .B(n35317), .Y(n37018) );
  NAND3X1 U30673 ( .A(wraddr[1]), .B(n36756), .C(wraddr[2]), .Y(n35317) );
  INVX1 U30674 ( .A(n37140), .Y(n36756) );
  NAND3X1 U30675 ( .A(n37141), .B(n37142), .C(n37143), .Y(n37140) );
  NOR2X1 U30676 ( .A(n37144), .B(n37145), .Y(n37143) );
  NAND2X1 U30677 ( .A(n37146), .B(wren), .Y(n37145) );
  MUX2X1 U30678 ( .B(n37138), .A(wrbyteen[14]), .S(n37137), .Y(n37146) );
  INVX1 U30679 ( .A(wrbyteen[13]), .Y(n37137) );
  OAI21X1 U30680 ( .A(wrbyteen[14]), .B(n37128), .C(wrbyteen[0]), .Y(n37144)
         );
  INVX1 U30681 ( .A(wrbyteen[15]), .Y(n37128) );
  MUX2X1 U30682 ( .B(n37147), .A(n37148), .S(n37127), .Y(n37142) );
  INVX1 U30683 ( .A(wrbyteen[7]), .Y(n37127) );
  OAI21X1 U30684 ( .A(wrbyteen[5]), .B(n37126), .C(n37149), .Y(n37148) );
  AOI21X1 U30685 ( .A(n37150), .B(n37151), .C(wrbyteen[8]), .Y(n37149) );
  NAND3X1 U30686 ( .A(n37130), .B(n37125), .C(n37152), .Y(n37150) );
  MUX2X1 U30687 ( .B(wrbyteen[3]), .A(n37028), .S(wrbyteen[2]), .Y(n37152) );
  INVX1 U30688 ( .A(wrbyteen[1]), .Y(n37028) );
  INVX1 U30689 ( .A(wrbyteen[5]), .Y(n37125) );
  INVX1 U30690 ( .A(wrbyteen[6]), .Y(n37126) );
  NAND3X1 U30691 ( .A(wrbyteen[5]), .B(n37153), .C(wrbyteen[6]), .Y(n37147) );
  INVX1 U30692 ( .A(n37151), .Y(n37153) );
  NAND3X1 U30693 ( .A(wrbyteen[2]), .B(wrbyteen[1]), .C(n37154), .Y(n37151) );
  NOR2X1 U30694 ( .A(n37129), .B(n37130), .Y(n37154) );
  INVX1 U30695 ( .A(wrbyteen[4]), .Y(n37130) );
  INVX1 U30696 ( .A(wrbyteen[3]), .Y(n37129) );
  NOR2X1 U30697 ( .A(n37155), .B(n37156), .Y(n37141) );
  MUX2X1 U30698 ( .B(wrbyteen[8]), .A(n37136), .S(n37139), .Y(n37156) );
  INVX1 U30699 ( .A(wrbyteen[9]), .Y(n37139) );
  INVX1 U30700 ( .A(wrbyteen[10]), .Y(n37136) );
  MUX2X1 U30701 ( .B(n37138), .A(wrbyteen[10]), .S(wrbyteen[11]), .Y(n37155)
         );
  INVX1 U30702 ( .A(wrbyteen[12]), .Y(n37138) );
  NAND3X1 U30703 ( .A(wraddr[3]), .B(wraddr[0]), .C(wraddr[4]), .Y(n36753) );
endmodule

