`timescale 1ns/10ps
/**
 * `timescale time_unit base / precision base
 *
 * -Specifies the time units and precision for delays:
 * -time_unit is the amount of time a delay of 1 represents.
 *	The time unit must be 1 10 or 100
 * -base is the time base for each unit, ranging from seconds
 *	to femtoseconds, and must be: s ms us ns ps or fs
 * -precision and base represent how many decimal points of
 *	precision to use relative to the time units.
 */

/**
 * This is written by Zhiyang Ong -student number 6004919412-
 * for EE577b Homework 4, Question 4
 */

// Testbench for behavioral model for the register file


// Import the modules that will be tested for in this testbench
`include "regfile.v"

// IMPORTANT: To run this, try: ncverilog -f regfile.f +gui
module tb_regfile();
	/**
	 * Depth = number of rows for the register file
	 *
	 * The construct base**exponent is not synthesizable for our
	 * tool and technology library set up. It should be with the latest
	 * version of Verilog, Verilog 2005
	 */
	parameter DEPTH = 8;			// DEPTH = 2^DEPTH_P2 = 2^3
	// Width of the register file
	parameter WIDTH = 8;
	
	
	
	
	
	
	
	// ============================================================
	/**
	 * Declare signal types for testbench to drive and monitor
	 * signals during the simulation of the register file
	 *
	 * The reg data type holds a value until a new value is driven
	 * onto it in an "initial" or "always" block. It can only be
	 * assigned a value in an "always" or "initial" block, and is
	 * used to apply stimulus to the inputs of the DUT.
	 *
	 * The wire type is a passive data type that holds a value driven
	 * onto it by a port, assign statement or reg type. Wires cannot be
	 * assigned values inside "always" and "initial" blocks. They can
	 * be used to hold the values of the DUT's outputs
	 */
	
	// Declare "wire" signals: outputs from the DUT
	// data_out & out_valid output signals
	wire [WIDTH-1:0] d_out;
	
	
	
	
	
	
	
	// ============================================================
	
	// Declare "reg" signals: inputs to the DUT
	// clk, wren
	reg clock,wr_en;
	// data_in
	reg [WIDTH-1:0] d_in;
	// wraddr, rdaddr
	reg [DEPTH-1:0] w_addr,r_addr ;
	
	
	
	
	
	
	
	
	// ============================================================
	// Counter for loop to enumerate all the values of r
	//integer count;
	
	
	
	
	
	
	
	
	
	
	
	
	// ============================================================
	
	/**
	 * Each sequential control block, such as the initial or always
	 * block, will execute concurrently in every module at the start
	 * of the simulation
	 */
	always begin
    	// Clock frequency is arbitrarily chosen; Period=10ns
    	#5 clock = 0;
    	#5 clock = 1;
    end	
	
	
	
	
	
	
	
	
	
	// ============================================================
	
	/**
	 * Instantiate an instance of regfile() so that
	 * inputs can be passed to the Device Under Test (DUT)
	 * Given instance name is "rg"
	 */
	regfile rg (
		// instance_name(signal name),
		// Signal name can be the same as the instance name
		d_out,d_in,w_addr,r_addr,wr_en,clock);
	
	
	
	
	// ============================================================
	
	/**
	 * Initial block start executing sequentially @ t=0
	 * If and when a delay is encountered, the execution of this block
	 * pauses or waits until the delay time has passed, before resuming
	 * execution
	 *
	 * Each intial or always block executes concurrently; that is,
	 * multiple "always" or "initial" blocks will execute simultaneously
	 *
	 * E.g.
	 * always
	 * begin
	 *		#10 clk_50 = ~clk_50; // Invert clock signal every 10 ns
	 *		// Clock signal has a period of 20 ns or 50 MHz
	 * end
	 */
	initial
	begin
		// "$time" indicates the current time in the simulation
		$display($time, " << Starting the simulation >>");
		// @ t=0; reset the sequence detector
		d_in=8'd6;
		w_addr=3'd0;
		r_addr=3'd0;
		wr_en=1;
		
		
		#10
		d_in=8'd7;
		w_addr=3'd0;
		r_addr=3'd0;
		wr_en=0;
		
		// Write...
		#10
		d_in=8'd6;
		w_addr=3'd2;
		r_addr=3'd0;
		wr_en=1;
		
		
		#10
		d_in=8'd5;
		w_addr=3'd3;
		r_addr=3'd1;
		wr_en=1;
		
		
		#10
		d_in=8'd100;
		w_addr=3'd4;
		r_addr=3'd7;
		wr_en=1;
		
		
		#10
		d_in=8'd200;
		w_addr=3'd5;
		r_addr=3'd6;
		wr_en=1;
		
		// Read...
		#10
		d_in=8'd3;
		w_addr=3'd4;
		r_addr=3'd2;
		wr_en=0;
		
		
		#10
		d_in=8'd2;
		w_addr=3'd5;
		r_addr=3'd3;
		wr_en=0;
		
		
		#10
		d_in=8'd1;
		w_addr=3'd6;
		r_addr=3'd4;
		wr_en=0;
		
		
		#10
		d_in=8'd0;
		w_addr=3'd7;
		r_addr=3'd5;
		wr_en=0;
		
		
		#10
		d_in=8'd5;
		w_addr=3'd7;
		r_addr=3'd1;
		wr_en=1;
		
		
		#10
		d_in=8'd0;
		w_addr=3'd2;
		r_addr=3'd7;
		wr_en=0;
		
		
		
		
		
		
		
		
		
		
		
		// end simulation
		#30
		
		$display($time, " << Finishing the simulation >>");
		$finish;
	end

endmodule
