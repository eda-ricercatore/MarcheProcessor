
module shift ( reg_A, reg_B, ctrl_ww, alu_op, result );
  input [0:127] reg_A;
  input [0:127] reg_B;
  input [0:1] ctrl_ww;
  input [0:4] alu_op;
  output [0:127] result;
  wire   n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
         n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038,
         n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046,
         n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054,
         n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062,
         n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070,
         n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
         n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086,
         n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094,
         n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102,
         n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
         n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118,
         n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126,
         n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134,
         n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142,
         n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150,
         n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158,
         n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166,
         n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
         n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182,
         n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190,
         n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
         n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206,
         n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214,
         n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222,
         n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230,
         n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238,
         n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
         n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254,
         n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262,
         n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270,
         n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278,
         n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286,
         n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294,
         n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302,
         n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310,
         n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
         n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326,
         n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334,
         n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342,
         n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350,
         n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358,
         n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366,
         n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374,
         n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382,
         n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
         n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398,
         n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
         n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414,
         n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422,
         n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430,
         n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
         n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446,
         n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454,
         n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
         n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470,
         n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
         n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486,
         n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494,
         n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502,
         n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
         n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
         n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526,
         n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
         n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542,
         n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
         n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558,
         n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566,
         n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574,
         n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
         n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590,
         n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598,
         n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606,
         n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614,
         n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
         n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630,
         n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638,
         n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646,
         n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654,
         n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
         n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670,
         n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
         n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686,
         n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
         n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702,
         n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710,
         n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
         n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
         n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734,
         n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742,
         n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
         n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758,
         n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
         n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774,
         n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782,
         n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
         n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798,
         n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806,
         n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814,
         n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
         n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830,
         n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
         n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846,
         n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854,
         n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862,
         n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
         n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878,
         n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
         n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
         n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902,
         n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
         n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918,
         n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
         n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934,
         n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
         n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950,
         n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
         n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
         n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974,
         n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
         n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990,
         n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998,
         n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006,
         n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
         n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022,
         n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030,
         n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038,
         n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046,
         n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
         n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
         n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070,
         n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078,
         n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086,
         n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094,
         n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102,
         n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110,
         n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118,
         n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
         n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
         n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142,
         n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
         n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
         n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
         n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174,
         n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
         n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190,
         n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
         n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
         n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214,
         n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222,
         n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
         n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238,
         n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246,
         n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
         n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
         n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
         n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278,
         n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286,
         n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294,
         n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
         n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310,
         n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318,
         n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326,
         n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334,
         n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
         n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350,
         n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358,
         n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366,
         n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374,
         n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382,
         n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390,
         n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
         n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406,
         n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
         n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422,
         n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430,
         n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438,
         n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446,
         n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454,
         n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462,
         n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470,
         n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478,
         n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486,
         n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494,
         n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502,
         n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510,
         n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518,
         n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526,
         n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534,
         n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542,
         n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550,
         n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558,
         n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566,
         n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574,
         n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582,
         n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590,
         n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598,
         n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606,
         n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614,
         n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622,
         n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630,
         n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638,
         n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646,
         n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654,
         n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662,
         n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670,
         n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678,
         n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686,
         n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694,
         n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702,
         n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
         n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718,
         n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726,
         n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734,
         n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742,
         n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750,
         n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758,
         n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766,
         n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
         n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782,
         n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790,
         n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798,
         n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
         n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814,
         n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822,
         n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830,
         n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838,
         n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
         n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854,
         n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862,
         n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870,
         n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
         n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886,
         n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894,
         n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902,
         n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910,
         n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
         n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926,
         n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934,
         n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
         n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950,
         n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958,
         n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966,
         n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
         n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982,
         n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990,
         n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998,
         n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006,
         n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014,
         n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022,
         n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030,
         n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038,
         n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046,
         n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054,
         n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062,
         n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070,
         n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078,
         n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
         n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094,
         n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102,
         n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110,
         n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
         n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126,
         n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
         n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142,
         n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150,
         n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158,
         n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166,
         n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174,
         n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182,
         n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190,
         n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198,
         n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206,
         n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214,
         n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222,
         n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
         n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238,
         n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246,
         n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254,
         n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262,
         n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270,
         n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
         n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286,
         n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294,
         n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302,
         n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310,
         n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318,
         n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326,
         n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334,
         n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342,
         n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350,
         n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358,
         n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366,
         n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
         n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382,
         n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390,
         n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398,
         n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406,
         n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414,
         n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422,
         n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430,
         n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438,
         n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
         n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454,
         n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462,
         n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470,
         n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
         n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486,
         n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494,
         n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502,
         n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510,
         n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518,
         n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526,
         n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534,
         n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542,
         n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550,
         n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558,
         n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566,
         n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574,
         n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582,
         n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590,
         n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
         n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606,
         n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614,
         n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622,
         n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630,
         n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638,
         n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646,
         n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654,
         n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662,
         n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670,
         n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678,
         n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686,
         n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694,
         n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702,
         n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710,
         n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718,
         n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726,
         n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734,
         n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742,
         n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750,
         n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758,
         n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
         n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774,
         n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
         n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790,
         n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798,
         n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
         n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814,
         n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822,
         n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830,
         n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838,
         n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846,
         n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
         n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862,
         n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870,
         n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
         n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886,
         n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894,
         n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902,
         n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
         n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918,
         n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
         n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934,
         n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942,
         n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950,
         n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958,
         n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966,
         n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974,
         n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982,
         n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990,
         n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998,
         n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006,
         n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014,
         n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022,
         n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030,
         n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038,
         n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046,
         n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054,
         n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062,
         n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070,
         n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078,
         n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086,
         n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094,
         n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
         n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110,
         n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118,
         n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126,
         n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134,
         n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142,
         n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150,
         n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158,
         n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166,
         n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174,
         n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182,
         n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190,
         n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198,
         n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206,
         n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214,
         n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222,
         n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230,
         n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238,
         n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246,
         n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254,
         n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262,
         n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270,
         n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278,
         n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286,
         n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
         n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
         n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310,
         n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318,
         n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326,
         n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334,
         n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
         n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350,
         n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358,
         n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366,
         n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374,
         n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382,
         n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390,
         n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398,
         n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406,
         n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
         n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422,
         n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430,
         n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
         n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446,
         n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
         n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
         n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470,
         n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478,
         n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486,
         n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494,
         n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
         n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
         n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518,
         n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526,
         n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534,
         n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542,
         n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550,
         n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558,
         n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566,
         n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
         n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582,
         n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590,
         n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598,
         n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606,
         n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614,
         n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622,
         n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630,
         n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638,
         n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
         n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654,
         n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662,
         n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670,
         n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678,
         n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686,
         n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694,
         n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
         n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710,
         n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
         n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726,
         n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734,
         n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742,
         n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750,
         n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758,
         n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766,
         n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
         n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782,
         n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
         n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798,
         n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806,
         n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814,
         n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822,
         n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830,
         n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838,
         n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846,
         n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854,
         n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
         n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870,
         n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878,
         n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886,
         n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894,
         n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902,
         n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910,
         n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918,
         n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
         n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934,
         n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942,
         n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950,
         n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958,
         n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
         n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974,
         n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982,
         n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990,
         n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
         n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006,
         n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014,
         n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022,
         n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030,
         n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038,
         n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046,
         n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054,
         n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
         n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
         n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
         n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086,
         n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094,
         n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102,
         n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
         n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118,
         n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126,
         n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
         n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142,
         n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150,
         n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158,
         n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166,
         n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
         n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182,
         n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190,
         n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198,
         n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
         n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
         n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
         n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
         n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238,
         n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
         n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
         n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262,
         n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270,
         n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
         n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
         n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
         n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302,
         n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310,
         n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318,
         n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326,
         n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334,
         n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342,
         n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
         n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358,
         n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
         n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374,
         n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382,
         n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390,
         n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398,
         n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406,
         n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414,
         n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
         n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430,
         n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
         n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446,
         n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454,
         n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
         n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
         n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478,
         n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
         n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
         n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502,
         n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510,
         n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518,
         n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526,
         n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534,
         n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542,
         n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550,
         n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558,
         n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
         n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574,
         n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582,
         n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590,
         n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598,
         n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606,
         n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614,
         n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622,
         n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630,
         n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
         n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646,
         n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654,
         n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
         n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670,
         n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678,
         n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686,
         n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694,
         n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702,
         n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
         n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
         n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
         n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742,
         n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
         n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758,
         n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766,
         n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774,
         n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
         n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790,
         n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
         n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806,
         n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814,
         n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822,
         n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
         n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
         n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862,
         n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
         n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
         n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886,
         n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894,
         n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
         n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
         n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918,
         n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
         n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934,
         n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
         n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950,
         n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958,
         n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
         n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
         n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982,
         n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
         n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
         n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006,
         n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
         n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022,
         n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030,
         n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
         n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046,
         n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
         n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062,
         n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
         n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
         n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
         n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
         n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102,
         n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
         n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
         n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126,
         n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
         n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
         n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150,
         n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
         n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166,
         n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174,
         n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
         n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
         n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198,
         n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
         n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
         n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222,
         n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
         n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238,
         n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246,
         n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
         n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
         n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270,
         n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278,
         n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
         n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294,
         n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
         n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310,
         n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318,
         n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326,
         n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
         n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342,
         n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350,
         n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
         n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366,
         n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
         n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
         n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390,
         n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
         n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
         n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414,
         n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
         n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
         n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438,
         n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
         n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
         n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462,
         n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470,
         n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478,
         n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
         n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
         n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510,
         n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
         n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526,
         n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534,
         n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
         n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
         n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
         n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566,
         n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
         n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582,
         n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
         n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598,
         n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606,
         n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
         n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
         n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630,
         n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638,
         n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
         n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654,
         n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662,
         n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670,
         n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678,
         n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686,
         n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694,
         n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702,
         n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710,
         n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
         n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726,
         n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
         n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742,
         n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750,
         n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758,
         n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766,
         n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774,
         n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782,
         n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
         n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798,
         n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
         n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814,
         n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822,
         n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
         n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
         n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846,
         n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854,
         n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
         n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870,
         n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878,
         n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886,
         n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894,
         n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902,
         n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910,
         n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918,
         n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926,
         n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
         n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942,
         n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950,
         n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958,
         n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966,
         n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974,
         n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982,
         n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990,
         n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998,
         n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006,
         n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014,
         n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022,
         n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030,
         n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038,
         n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046,
         n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
         n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062,
         n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070,
         n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
         n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086,
         n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
         n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110,
         n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118,
         n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
         n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134,
         n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142,
         n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150,
         n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158,
         n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166,
         n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174,
         n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182,
         n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190,
         n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
         n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206,
         n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214,
         n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
         n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230,
         n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
         n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246,
         n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254,
         n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262,
         n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270,
         n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278,
         n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286,
         n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294,
         n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302,
         n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
         n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318,
         n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326,
         n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
         n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342,
         n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350,
         n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358,
         n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366,
         n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374,
         n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382,
         n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390,
         n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398,
         n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406,
         n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414,
         n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422,
         n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430,
         n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
         n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446,
         n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454,
         n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462,
         n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470,
         n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
         n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
         n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494,
         n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502,
         n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
         n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518,
         n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
         n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
         n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542,
         n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
         n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
         n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566,
         n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574,
         n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582,
         n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590,
         n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
         n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606,
         n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614,
         n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622,
         n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630,
         n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638,
         n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646,
         n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
         n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662,
         n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
         n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678,
         n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686,
         n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694,
         n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702,
         n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710,
         n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718,
         n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726,
         n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734,
         n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
         n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750,
         n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758,
         n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766,
         n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
         n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782,
         n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790,
         n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798,
         n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806,
         n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814,
         n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822,
         n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830,
         n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838,
         n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846,
         n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854,
         n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862,
         n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870,
         n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878,
         n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886,
         n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894,
         n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902,
         n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910,
         n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918,
         n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926,
         n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934,
         n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942,
         n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950,
         n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
         n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966,
         n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
         n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
         n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990,
         n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998,
         n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006,
         n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
         n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
         n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
         n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
         n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046,
         n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054,
         n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062,
         n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070,
         n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078,
         n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
         n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094,
         n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
         n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110,
         n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118,
         n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126,
         n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134,
         n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142,
         n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150,
         n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
         n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166,
         n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
         n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182,
         n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190,
         n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198,
         n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206,
         n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214,
         n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222,
         n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
         n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238,
         n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
         n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254,
         n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262,
         n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270,
         n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278,
         n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286,
         n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294,
         n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
         n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310,
         n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318,
         n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
         n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334,
         n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342,
         n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350,
         n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358,
         n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366,
         n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
         n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382,
         n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
         n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398,
         n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406,
         n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414,
         n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422,
         n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430,
         n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
         n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446,
         n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454,
         n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462,
         n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470,
         n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478,
         n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486,
         n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494,
         n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502,
         n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
         n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
         n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526,
         n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534,
         n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542,
         n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550,
         n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558,
         n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566,
         n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574,
         n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
         n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590,
         n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598,
         n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606,
         n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614,
         n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622,
         n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630,
         n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638,
         n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646,
         n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654,
         n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662,
         n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670,
         n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
         n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
         n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694,
         n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
         n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
         n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718,
         n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
         n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
         n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742,
         n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
         n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
         n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766,
         n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
         n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
         n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
         n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
         n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
         n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
         n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
         n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
         n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
         n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
         n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
         n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
         n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030,
         n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
         n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
         n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054,
         n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
         n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
         n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
         n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
         n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102,
         n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
         n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
         n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
         n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
         n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
         n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
         n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158,
         n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
         n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174,
         n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
         n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
         n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198,
         n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
         n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
         n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222,
         n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230,
         n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
         n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
         n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
         n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
         n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270,
         n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
         n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
         n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294,
         n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
         n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
         n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
         n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342,
         n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
         n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
         n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366,
         n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
         n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
         n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390,
         n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
         n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
         n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
         n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
         n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
         n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446,
         n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462,
         n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
         n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
         n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486,
         n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
         n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
         n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
         n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
         n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
         n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534,
         n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
         n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
         n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
         n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
         n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
         n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
         n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590,
         n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
         n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182,
         n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
         n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
         n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206,
         n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
         n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
         n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230,
         n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238,
         n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
         n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254,
         n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
         n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
         n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278,
         n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
         n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
         n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302,
         n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310,
         n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
         n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326,
         n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
         n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
         n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350,
         n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
         n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366,
         n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374,
         n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382,
         n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
         n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398,
         n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
         n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
         n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422,
         n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
         n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
         n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446,
         n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454,
         n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
         n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470,
         n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
         n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
         n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494,
         n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
         n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
         n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518,
         n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
         n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
         n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542,
         n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
         n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558,
         n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566,
         n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
         n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582,
         n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590,
         n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
         n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
         n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614,
         n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
         n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
         n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638,
         n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646,
         n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654,
         n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662,
         n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670,
         n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
         n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686,
         n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
         n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702,
         n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710,
         n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718,
         n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726,
         n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734,
         n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742,
         n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
         n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758,
         n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
         n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774,
         n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782,
         n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790,
         n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798,
         n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806,
         n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814,
         n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
         n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830,
         n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
         n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846,
         n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854,
         n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862,
         n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
         n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878,
         n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886,
         n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
         n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902,
         n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
         n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918,
         n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926,
         n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
         n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
         n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950,
         n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958,
         n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
         n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974,
         n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
         n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990,
         n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
         n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
         n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014,
         n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022,
         n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030,
         n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
         n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046,
         n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
         n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
         n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
         n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
         n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
         n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
         n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102,
         n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
         n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
         n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
         n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134,
         n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142,
         n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
         n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158,
         n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166,
         n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
         n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
         n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190,
         n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
         n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206,
         n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214,
         n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
         n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230,
         n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238,
         n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246,
         n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
         n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262,
         n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
         n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278,
         n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286,
         n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294,
         n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
         n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310,
         n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318,
         n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
         n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334,
         n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
         n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350,
         n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358,
         n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
         n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374,
         n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382,
         n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390,
         n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
         n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406,
         n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
         n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422,
         n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430,
         n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
         n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
         n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454,
         n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462,
         n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
         n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478,
         n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
         n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
         n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502,
         n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
         n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518,
         n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526,
         n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534,
         n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
         n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550,
         n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
         n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
         n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574,
         n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
         n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590,
         n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598,
         n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606,
         n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
         n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622,
         n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
         n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638,
         n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646,
         n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
         n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662,
         n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670,
         n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678,
         n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
         n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694,
         n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
         n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
         n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718,
         n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726,
         n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734,
         n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742,
         n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
         n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
         n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766,
         n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
         n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
         n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790,
         n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798,
         n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806,
         n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814,
         n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
         n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838,
         n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
         n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
         n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862,
         n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870,
         n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878,
         n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886,
         n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
         n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
         n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910,
         n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
         n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926,
         n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934,
         n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942,
         n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
         n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958,
         n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
         n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
         n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982,
         n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
         n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022,
         n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
         n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038,
         n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
         n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054,
         n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
         n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
         n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
         n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
         n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
         n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102,
         n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110,
         n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
         n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126,
         n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
         n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142,
         n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150,
         n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158,
         n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166,
         n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174,
         n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182,
         n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
         n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198,
         n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
         n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214,
         n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222,
         n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230,
         n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238,
         n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246,
         n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254,
         n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
         n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270,
         n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
         n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286,
         n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294,
         n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302,
         n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
         n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318,
         n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326,
         n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
         n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342,
         n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
         n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358,
         n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366,
         n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374,
         n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
         n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390,
         n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398,
         n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
         n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
         n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
         n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
         n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438,
         n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446,
         n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
         n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486,
         n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
         n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502,
         n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510,
         n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
         n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
         n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534,
         n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542,
         n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
         n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558,
         n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
         n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574,
         n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582,
         n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590,
         n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
         n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606,
         n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614,
         n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
         n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
         n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
         n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646,
         n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654,
         n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662,
         n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
         n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678,
         n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686,
         n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
         n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
         n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
         n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718,
         n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726,
         n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
         n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742,
         n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750,
         n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758,
         n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
         n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
         n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
         n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790,
         n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798,
         n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
         n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
         n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822,
         n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830,
         n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
         n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846,
         n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
         n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
         n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
         n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
         n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886,
         n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894,
         n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902,
         n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
         n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918,
         n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
         n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
         n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942,
         n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
         n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958,
         n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966,
         n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974,
         n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
         n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990,
         n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
         n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006,
         n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014,
         n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
         n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030,
         n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
         n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046,
         n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
         n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062,
         n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
         n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
         n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086,
         n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
         n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102,
         n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110,
         n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118,
         n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
         n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134,
         n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
         n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
         n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158,
         n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166,
         n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174,
         n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182,
         n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190,
         n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
         n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206,
         n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214,
         n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222,
         n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230,
         n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238,
         n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
         n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254,
         n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262,
         n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
         n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278,
         n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286,
         n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294,
         n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302,
         n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310,
         n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318,
         n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326,
         n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334,
         n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
         n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350,
         n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358,
         n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366,
         n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374,
         n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
         n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390,
         n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398,
         n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406,
         n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
         n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422,
         n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430,
         n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438,
         n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446,
         n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454,
         n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462,
         n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470,
         n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478,
         n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486,
         n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494,
         n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502,
         n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510,
         n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
         n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526,
         n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534,
         n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542,
         n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550,
         n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558,
         n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566,
         n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574,
         n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
         n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590,
         n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598,
         n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606,
         n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614,
         n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622,
         n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630,
         n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638,
         n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646,
         n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
         n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662,
         n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670,
         n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678,
         n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686,
         n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694,
         n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702,
         n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710,
         n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
         n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726,
         n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734,
         n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742,
         n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750,
         n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758,
         n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766,
         n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774,
         n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782,
         n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790,
         n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798,
         n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806,
         n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814,
         n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822,
         n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830,
         n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838,
         n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
         n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854,
         n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862,
         n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870,
         n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878,
         n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886,
         n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894,
         n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902,
         n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
         n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918,
         n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926,
         n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934,
         n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942,
         n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950,
         n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958,
         n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966,
         n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974,
         n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982,
         n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990,
         n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998,
         n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
         n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014,
         n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022,
         n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
         n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038,
         n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046,
         n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054,
         n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062,
         n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070,
         n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
         n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086,
         n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094,
         n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102,
         n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110,
         n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118,
         n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126,
         n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134,
         n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142,
         n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
         n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158,
         n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166,
         n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174,
         n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182,
         n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190,
         n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198,
         n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206,
         n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214,
         n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
         n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230,
         n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238,
         n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246,
         n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254,
         n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262,
         n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270,
         n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278,
         n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286,
         n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
         n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
         n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310,
         n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
         n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326,
         n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334,
         n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342,
         n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
         n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358,
         n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
         n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374,
         n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382,
         n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390,
         n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398,
         n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406,
         n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414,
         n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
         n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430,
         n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
         n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
         n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454,
         n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462,
         n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470,
         n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478,
         n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486,
         n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
         n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502,
         n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510,
         n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518,
         n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526,
         n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534,
         n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542,
         n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550,
         n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558,
         n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
         n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574,
         n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582,
         n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590,
         n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598,
         n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606,
         n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614,
         n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622,
         n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630,
         n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
         n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646,
         n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654,
         n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662,
         n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670,
         n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678,
         n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
         n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694,
         n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702,
         n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
         n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718,
         n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726,
         n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734,
         n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742,
         n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750,
         n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
         n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766,
         n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774,
         n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
         n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790,
         n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798,
         n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806,
         n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814,
         n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822,
         n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830,
         n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838,
         n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846,
         n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
         n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862,
         n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
         n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878,
         n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886,
         n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894,
         n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902,
         n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910,
         n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918,
         n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
         n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934,
         n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942,
         n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950,
         n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958,
         n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966,
         n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974,
         n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982,
         n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990,
         n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
         n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006,
         n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
         n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022,
         n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030,
         n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038,
         n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046,
         n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054,
         n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062,
         n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
         n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078,
         n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
         n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094,
         n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102,
         n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110,
         n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118,
         n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126,
         n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134,
         n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
         n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150,
         n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158,
         n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166,
         n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174,
         n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
         n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190,
         n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198,
         n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206,
         n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
         n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222,
         n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230,
         n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238,
         n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246,
         n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254,
         n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262,
         n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270,
         n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
         n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
         n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294,
         n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302,
         n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310,
         n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318,
         n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326,
         n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334,
         n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342,
         n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350,
         n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358,
         n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366,
         n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374,
         n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382,
         n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390,
         n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
         n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406,
         n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414,
         n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422,
         n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430,
         n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438,
         n39439, n39440, n39441;

  INVX2 U20376 ( .A(reg_A[116]), .Y(n25337) );
  INVX1 U20377 ( .A(n26267), .Y(n25023) );
  INVX1 U20378 ( .A(n25932), .Y(n25024) );
  BUFX2 U20379 ( .A(n26034), .Y(n25025) );
  BUFX2 U20380 ( .A(n26210), .Y(n25026) );
  INVX1 U20381 ( .A(n25222), .Y(n25027) );
  INVX1 U20382 ( .A(n25123), .Y(n25028) );
  INVX1 U20383 ( .A(n26999), .Y(n25029) );
  INVX2 U20384 ( .A(n25628), .Y(n25030) );
  INVX2 U20385 ( .A(n26504), .Y(n25031) );
  INVX4 U20386 ( .A(n25342), .Y(n26504) );
  INVX2 U20387 ( .A(n25188), .Y(n25032) );
  INVX2 U20388 ( .A(n25087), .Y(n25382) );
  INVX2 U20389 ( .A(n26990), .Y(n25310) );
  INVX2 U20390 ( .A(n25253), .Y(n25033) );
  INVX2 U20391 ( .A(n25124), .Y(n25034) );
  INVX2 U20392 ( .A(n25234), .Y(n25035) );
  INVX4 U20393 ( .A(n25794), .Y(n25188) );
  INVX4 U20394 ( .A(n26147), .Y(n26267) );
  INVX2 U20395 ( .A(n25637), .Y(n25036) );
  INVX2 U20396 ( .A(n25629), .Y(n25037) );
  INVX2 U20397 ( .A(n25487), .Y(n25038) );
  INVX2 U20398 ( .A(n25243), .Y(n25487) );
  INVX2 U20399 ( .A(n25325), .Y(n25039) );
  INVX4 U20400 ( .A(n25229), .Y(n25325) );
  INVX4 U20401 ( .A(n25475), .Y(n25234) );
  INVX4 U20402 ( .A(n25219), .Y(n25637) );
  INVX4 U20403 ( .A(n25223), .Y(n25629) );
  INVX4 U20404 ( .A(n25252), .Y(n25040) );
  INVX4 U20405 ( .A(n25133), .Y(n25252) );
  INVX4 U20406 ( .A(n25136), .Y(n25041) );
  INVX4 U20407 ( .A(n25254), .Y(n25136) );
  INVX4 U20408 ( .A(n25135), .Y(n25042) );
  INVX4 U20409 ( .A(n25784), .Y(n25135) );
  INVX4 U20410 ( .A(n25125), .Y(n25043) );
  INVX4 U20411 ( .A(n25228), .Y(n25125) );
  INVX4 U20412 ( .A(n25403), .Y(n25044) );
  INVX4 U20413 ( .A(n25473), .Y(n25222) );
  INVX4 U20414 ( .A(n25467), .Y(n25124) );
  INVX4 U20415 ( .A(n25131), .Y(n25253) );
  INVX8 U20416 ( .A(n26703), .Y(n25123) );
  INVX8 U20417 ( .A(n25129), .Y(n25628) );
  INVX2 U20418 ( .A(n30208), .Y(n25045) );
  INVX2 U20419 ( .A(reg_A[74]), .Y(n26438) );
  INVX2 U20420 ( .A(reg_A[87]), .Y(n25965) );
  INVX2 U20421 ( .A(reg_A[41]), .Y(n30463) );
  INVX2 U20422 ( .A(n25339), .Y(n25046) );
  INVX4 U20423 ( .A(n25238), .Y(n25339) );
  INVX2 U20424 ( .A(reg_A[15]), .Y(n29279) );
  INVX2 U20425 ( .A(n25246), .Y(n25047) );
  INVX4 U20426 ( .A(n25336), .Y(n25246) );
  INVX2 U20427 ( .A(reg_A[93]), .Y(n25881) );
  INVX2 U20428 ( .A(n25247), .Y(n25048) );
  INVX4 U20429 ( .A(n25334), .Y(n25247) );
  INVX2 U20430 ( .A(reg_A[40]), .Y(n30744) );
  INVX2 U20431 ( .A(reg_A[55]), .Y(n30043) );
  INVX2 U20432 ( .A(reg_A[14]), .Y(n25208) );
  INVX2 U20433 ( .A(reg_A[47]), .Y(n30068) );
  INVX2 U20434 ( .A(reg_A[104]), .Y(n25298) );
  INVX2 U20435 ( .A(reg_A[8]), .Y(n26701) );
  INVX2 U20436 ( .A(reg_A[28]), .Y(n25244) );
  INVX2 U20437 ( .A(n25257), .Y(n25049) );
  INVX2 U20438 ( .A(reg_A[69]), .Y(n25856) );
  INVX2 U20439 ( .A(reg_A[84]), .Y(n26230) );
  INVX2 U20440 ( .A(reg_A[73]), .Y(n26439) );
  INVX2 U20441 ( .A(reg_A[21]), .Y(n25232) );
  INVX2 U20442 ( .A(reg_A[115]), .Y(n25335) );
  INVX2 U20443 ( .A(reg_A[45]), .Y(n30066) );
  INVX2 U20444 ( .A(n25338), .Y(n25050) );
  INVX2 U20445 ( .A(n25241), .Y(n25051) );
  INVX4 U20446 ( .A(n25331), .Y(n25241) );
  INVX2 U20447 ( .A(n25604), .Y(n25052) );
  INVX4 U20448 ( .A(n25415), .Y(n25604) );
  INVX2 U20449 ( .A(reg_A[6]), .Y(n26677) );
  INVX2 U20450 ( .A(reg_A[100]), .Y(n25436) );
  INVX2 U20451 ( .A(n25517), .Y(n25053) );
  INVX2 U20452 ( .A(reg_A[54]), .Y(n30168) );
  INVX2 U20453 ( .A(reg_A[44]), .Y(n30067) );
  INVX2 U20454 ( .A(n33966), .Y(n33809) );
  INVX2 U20455 ( .A(reg_A[13]), .Y(n25206) );
  INVX2 U20456 ( .A(n26337), .Y(n25838) );
  INVX2 U20457 ( .A(n26338), .Y(n26160) );
  INVX2 U20458 ( .A(reg_A[17]), .Y(n27953) );
  INVX2 U20459 ( .A(n30223), .Y(n30024) );
  INVX2 U20460 ( .A(reg_A[114]), .Y(n25771) );
  INVX2 U20461 ( .A(reg_A[88]), .Y(n26195) );
  INVX2 U20462 ( .A(reg_A[77]), .Y(n26286) );
  INVX2 U20463 ( .A(reg_A[121]), .Y(n25490) );
  INVX2 U20464 ( .A(reg_A[70]), .Y(n26256) );
  INVX2 U20465 ( .A(reg_A[61]), .Y(n29989) );
  INVX2 U20466 ( .A(n30931), .Y(n25203) );
  INVX2 U20467 ( .A(n26599), .Y(n27012) );
  INVX2 U20468 ( .A(n27455), .Y(n26602) );
  INVX2 U20469 ( .A(reg_A[68]), .Y(n26107) );
  INVX2 U20470 ( .A(n34167), .Y(n34000) );
  INVX2 U20471 ( .A(reg_A[105]), .Y(n25296) );
  INVX2 U20472 ( .A(reg_A[109]), .Y(n25474) );
  INVX2 U20473 ( .A(reg_A[79]), .Y(n25864) );
  INVX2 U20474 ( .A(reg_A[53]), .Y(n30299) );
  INVX2 U20475 ( .A(reg_A[51]), .Y(n30009) );
  INVX2 U20476 ( .A(reg_A[49]), .Y(n30174) );
  INVX2 U20477 ( .A(reg_A[1]), .Y(n25177) );
  INVX2 U20478 ( .A(n27575), .Y(n26601) );
  INVX2 U20479 ( .A(reg_A[33]), .Y(n30170) );
  INVX2 U20480 ( .A(reg_A[97]), .Y(n25287) );
  INVX2 U20481 ( .A(reg_A[72]), .Y(n26547) );
  INVX2 U20482 ( .A(reg_A[76]), .Y(n25863) );
  INVX2 U20483 ( .A(reg_A[89]), .Y(n25929) );
  INVX2 U20484 ( .A(reg_A[3]), .Y(n25130) );
  INVX2 U20485 ( .A(reg_A[113]), .Y(n25483) );
  INVX2 U20486 ( .A(reg_A[38]), .Y(n30060) );
  INVX2 U20487 ( .A(n34012), .Y(n32934) );
  INVX2 U20488 ( .A(n25857), .Y(n25054) );
  INVX2 U20489 ( .A(reg_A[20]), .Y(n30587) );
  INVX2 U20490 ( .A(reg_A[52]), .Y(n30378) );
  INVX2 U20491 ( .A(reg_A[111]), .Y(n25452) );
  INVX2 U20492 ( .A(n26663), .Y(n25055) );
  INVX2 U20493 ( .A(n26996), .Y(n26480) );
  INVX2 U20494 ( .A(reg_A[36]), .Y(n30058) );
  INVX2 U20495 ( .A(n32194), .Y(n25608) );
  INVX2 U20496 ( .A(n25122), .Y(n25056) );
  INVX2 U20497 ( .A(reg_A[2]), .Y(n25128) );
  INVX2 U20498 ( .A(n25647), .Y(n25057) );
  INVX2 U20499 ( .A(n25320), .Y(n25647) );
  INVX1 U20500 ( .A(n26038), .Y(n25058) );
  INVX2 U20501 ( .A(n26981), .Y(n26038) );
  INVX2 U20502 ( .A(reg_A[18]), .Y(n25224) );
  INVX2 U20503 ( .A(n26151), .Y(n26186) );
  INVX2 U20504 ( .A(reg_A[32]), .Y(n30395) );
  INVX2 U20505 ( .A(reg_A[19]), .Y(n25220) );
  INVX2 U20506 ( .A(reg_A[99]), .Y(n25396) );
  INVX2 U20507 ( .A(n27523), .Y(n26045) );
  INVX2 U20508 ( .A(reg_A[39]), .Y(n30059) );
  INVX2 U20509 ( .A(reg_A[82]), .Y(n25874) );
  INVX2 U20510 ( .A(reg_A[65]), .Y(n25855) );
  INVX2 U20511 ( .A(n26208), .Y(n26530) );
  INVX2 U20512 ( .A(reg_A[22]), .Y(n25230) );
  INVX2 U20513 ( .A(reg_A[64]), .Y(n25853) );
  INVX2 U20514 ( .A(reg_A[102]), .Y(n25361) );
  INVX2 U20515 ( .A(n36246), .Y(n25355) );
  INVX2 U20516 ( .A(reg_A[50]), .Y(n30008) );
  INVX2 U20517 ( .A(n26432), .Y(n25059) );
  INVX2 U20518 ( .A(reg_A[81]), .Y(n26094) );
  INVX2 U20519 ( .A(n26924), .Y(n25060) );
  INVX2 U20520 ( .A(n30038), .Y(n29987) );
  INVX2 U20521 ( .A(n25097), .Y(n25403) );
  INVX2 U20522 ( .A(n27454), .Y(n26597) );
  INVX2 U20523 ( .A(n36136), .Y(n25399) );
  INVX2 U20524 ( .A(n29558), .Y(n25616) );
  INVX2 U20525 ( .A(reg_A[98]), .Y(n25289) );
  INVX2 U20526 ( .A(reg_A[35]), .Y(n30393) );
  INVX2 U20527 ( .A(n26878), .Y(n25061) );
  INVX2 U20528 ( .A(n25745), .Y(n26878) );
  INVX2 U20529 ( .A(n25264), .Y(n26761) );
  INVX2 U20530 ( .A(reg_A[34]), .Y(n30394) );
  INVX2 U20531 ( .A(n30320), .Y(n30212) );
  INVX2 U20532 ( .A(reg_A[7]), .Y(n25132) );
  INVX2 U20533 ( .A(n29970), .Y(n30846) );
  INVX2 U20534 ( .A(reg_A[16]), .Y(n25250) );
  INVX2 U20535 ( .A(n25491), .Y(n25338) );
  INVX2 U20536 ( .A(n30210), .Y(n30847) );
  INVX2 U20537 ( .A(reg_A[112]), .Y(n25476) );
  INVX2 U20538 ( .A(n29305), .Y(n25258) );
  INVX2 U20539 ( .A(n26758), .Y(n25142) );
  INVX2 U20540 ( .A(reg_A[66]), .Y(n25884) );
  INVX2 U20541 ( .A(reg_A[71]), .Y(n26101) );
  INVX2 U20542 ( .A(n30951), .Y(n25840) );
  INVX2 U20543 ( .A(n35474), .Y(n26032) );
  INVX2 U20544 ( .A(n25748), .Y(n26803) );
  INVX2 U20545 ( .A(reg_A[103]), .Y(n25448) );
  INVX2 U20546 ( .A(n25262), .Y(n25156) );
  INVX2 U20547 ( .A(reg_A[80]), .Y(n25584) );
  INVX2 U20548 ( .A(reg_A[67]), .Y(n25851) );
  INVX2 U20549 ( .A(n31398), .Y(n25607) );
  INVX2 U20550 ( .A(n25568), .Y(n25700) );
  INVX2 U20551 ( .A(n25914), .Y(n26276) );
  INVX2 U20552 ( .A(n26169), .Y(n26149) );
  INVX2 U20553 ( .A(reg_A[48]), .Y(n29655) );
  INVX2 U20554 ( .A(n26801), .Y(n25749) );
  INVX2 U20555 ( .A(n25747), .Y(n26804) );
  INVX2 U20556 ( .A(n26168), .Y(n26148) );
  INVX2 U20557 ( .A(n26927), .Y(n25062) );
  INVX2 U20558 ( .A(n25697), .Y(n25170) );
  INVX2 U20559 ( .A(n25972), .Y(n25984) );
  INVX2 U20560 ( .A(n27438), .Y(n25932) );
  INVX2 U20561 ( .A(n25397), .Y(n25793) );
  INVX2 U20562 ( .A(n26800), .Y(n25750) );
  INVX2 U20563 ( .A(n27253), .Y(n25614) );
  INVX2 U20564 ( .A(n26664), .Y(n25063) );
  INVX4 U20565 ( .A(n26936), .Y(n25613) );
  INVX4 U20566 ( .A(n25492), .Y(n25242) );
  INVX2 U20567 ( .A(n25635), .Y(n25064) );
  INVX4 U20568 ( .A(n25231), .Y(n25635) );
  INVX2 U20569 ( .A(n25235), .Y(n25065) );
  INVX4 U20570 ( .A(n25482), .Y(n25235) );
  INVX4 U20571 ( .A(n27252), .Y(n25615) );
  INVX4 U20572 ( .A(n26719), .Y(n25257) );
  BUFX2 U20573 ( .A(n25122), .Y(n25067) );
  BUFX2 U20574 ( .A(n25122), .Y(n25066) );
  BUFX2 U20575 ( .A(n25122), .Y(n25068) );
  BUFX2 U20576 ( .A(n25122), .Y(n25069) );
  BUFX2 U20577 ( .A(n25122), .Y(n25070) );
  BUFX2 U20578 ( .A(n25122), .Y(n25074) );
  BUFX2 U20579 ( .A(n25122), .Y(n25071) );
  BUFX2 U20580 ( .A(n25122), .Y(n25073) );
  BUFX2 U20581 ( .A(n25122), .Y(n25072) );
  BUFX2 U20582 ( .A(n25122), .Y(n25075) );
  NAND3X1 U20583 ( .A(n25076), .B(n25077), .C(n25078), .Y(result[9]) );
  NOR2X1 U20584 ( .A(n25079), .B(n25080), .Y(n25078) );
  NAND3X1 U20585 ( .A(n25081), .B(n25082), .C(n25083), .Y(n25080) );
  NOR2X1 U20586 ( .A(n25084), .B(n25085), .Y(n25083) );
  OAI21X1 U20587 ( .A(n25086), .B(n25087), .C(n25088), .Y(n25085) );
  AOI21X1 U20588 ( .A(n25089), .B(n25090), .C(n25091), .Y(n25086) );
  OAI21X1 U20589 ( .A(n25092), .B(n25093), .C(n25094), .Y(n25091) );
  OAI21X1 U20590 ( .A(n25095), .B(n25096), .C(n25044), .Y(n25094) );
  OAI21X1 U20591 ( .A(n25098), .B(n25099), .C(n25100), .Y(n25096) );
  AOI22X1 U20592 ( .A(n25101), .B(n25102), .C(n25103), .D(n25104), .Y(n25100)
         );
  OAI21X1 U20593 ( .A(n25105), .B(n25106), .C(n25107), .Y(n25095) );
  AOI22X1 U20594 ( .A(n25108), .B(n25109), .C(n25110), .D(n25111), .Y(n25107)
         );
  INVX1 U20595 ( .A(n25112), .Y(n25089) );
  INVX1 U20596 ( .A(n25113), .Y(n25084) );
  MUX2X1 U20597 ( .B(n25114), .A(n25115), .S(n25116), .Y(n25113) );
  OAI21X1 U20598 ( .A(n25117), .B(n25118), .C(n25119), .Y(n25082) );
  NAND2X1 U20599 ( .A(n25120), .B(n25121), .Y(n25118) );
  AOI22X1 U20600 ( .A(n25075), .B(reg_A[5]), .C(n25123), .D(reg_A[4]), .Y(
        n25121) );
  AOI22X1 U20601 ( .A(n25124), .B(reg_A[1]), .C(n25125), .D(reg_A[9]), .Y(
        n25120) );
  OR2X1 U20602 ( .A(n25126), .B(n25127), .Y(n25117) );
  OAI22X1 U20603 ( .A(n25128), .B(n25129), .C(n25130), .D(n25131), .Y(n25127)
         );
  OAI21X1 U20604 ( .A(n25132), .B(n25133), .C(n25134), .Y(n25126) );
  AOI22X1 U20605 ( .A(n25135), .B(reg_A[8]), .C(n25136), .D(reg_A[6]), .Y(
        n25134) );
  AOI22X1 U20606 ( .A(reg_A[0]), .B(n25137), .C(n25138), .D(reg_A[7]), .Y(
        n25081) );
  NAND3X1 U20607 ( .A(n25139), .B(n25140), .C(n25141), .Y(n25079) );
  AOI21X1 U20608 ( .A(n25142), .B(n25143), .C(n25144), .Y(n25141) );
  OAI22X1 U20609 ( .A(n25145), .B(n25146), .C(n25147), .D(n25148), .Y(n25144)
         );
  AOI22X1 U20610 ( .A(n25149), .B(reg_A[4]), .C(n25150), .D(n25151), .Y(n25140) );
  AOI22X1 U20611 ( .A(n25152), .B(reg_A[12]), .C(n25153), .D(reg_A[11]), .Y(
        n25139) );
  NOR2X1 U20612 ( .A(n25154), .B(n25155), .Y(n25077) );
  OAI21X1 U20613 ( .A(n25156), .B(n25157), .C(n25158), .Y(n25155) );
  AOI22X1 U20614 ( .A(n25159), .B(n25160), .C(n25161), .D(reg_A[3]), .Y(n25158) );
  INVX1 U20615 ( .A(n25162), .Y(n25161) );
  NAND3X1 U20616 ( .A(n25163), .B(n25164), .C(n25165), .Y(n25154) );
  AOI22X1 U20617 ( .A(n25166), .B(n25167), .C(n25168), .D(n25169), .Y(n25165)
         );
  NAND3X1 U20618 ( .A(n25170), .B(n25171), .C(n25172), .Y(n25164) );
  OAI21X1 U20619 ( .A(n25173), .B(n25174), .C(reg_A[8]), .Y(n25163) );
  NOR2X1 U20620 ( .A(n25175), .B(n25176), .Y(n25076) );
  OAI21X1 U20621 ( .A(n25177), .B(n25178), .C(n25179), .Y(n25176) );
  AOI22X1 U20622 ( .A(n25180), .B(reg_A[6]), .C(n25181), .D(reg_A[5]), .Y(
        n25179) );
  OR2X1 U20623 ( .A(n25182), .B(n25183), .Y(n25175) );
  OAI21X1 U20624 ( .A(n25184), .B(n25128), .C(n25185), .Y(n25183) );
  OAI21X1 U20625 ( .A(n25186), .B(n25187), .C(n25188), .Y(n25185) );
  OAI21X1 U20626 ( .A(n25189), .B(n25190), .C(n25191), .Y(n25187) );
  MUX2X1 U20627 ( .B(n25192), .A(n25193), .S(reg_B[14]), .Y(n25191) );
  OAI22X1 U20628 ( .A(n25194), .B(n25195), .C(n25196), .D(n25197), .Y(n25186)
         );
  OAI21X1 U20629 ( .A(n25198), .B(n25199), .C(n25200), .Y(n25182) );
  OAI21X1 U20630 ( .A(n25201), .B(n25202), .C(n25203), .Y(n25200) );
  OAI22X1 U20631 ( .A(n25204), .B(n25146), .C(n25205), .D(n25206), .Y(n25202)
         );
  OAI21X1 U20632 ( .A(n25207), .B(n25208), .C(n25209), .Y(n25201) );
  AOI22X1 U20633 ( .A(n25097), .B(n25210), .C(reg_A[15]), .D(n25211), .Y(
        n25209) );
  NAND3X1 U20634 ( .A(n25212), .B(n25213), .C(n25214), .Y(n25210) );
  AND2X1 U20635 ( .A(n25215), .B(n25216), .Y(n25214) );
  NOR2X1 U20636 ( .A(n25217), .B(n25218), .Y(n25216) );
  OAI21X1 U20637 ( .A(n25036), .B(n25220), .C(n25221), .Y(n25218) );
  AOI22X1 U20638 ( .A(reg_A[17]), .B(n25124), .C(reg_A[20]), .D(n25222), .Y(
        n25221) );
  OAI21X1 U20639 ( .A(n25037), .B(n25224), .C(n25225), .Y(n25217) );
  AOI22X1 U20640 ( .A(reg_A[13]), .B(n25070), .C(reg_A[14]), .D(n25123), .Y(
        n25225) );
  NOR2X1 U20641 ( .A(n25226), .B(n25227), .Y(n25215) );
  OAI22X1 U20642 ( .A(n25146), .B(n25228), .C(n25039), .D(n25230), .Y(n25227)
         );
  OAI21X1 U20643 ( .A(n25064), .B(n25232), .C(n25233), .Y(n25226) );
  AOI22X1 U20644 ( .A(reg_A[23]), .B(n25234), .C(reg_A[24]), .D(n25235), .Y(
        n25233) );
  NOR2X1 U20645 ( .A(n25236), .B(n25237), .Y(n25213) );
  OAI21X1 U20646 ( .A(n25046), .B(n25239), .C(n25240), .Y(n25237) );
  AOI22X1 U20647 ( .A(reg_A[27]), .B(n25241), .C(reg_A[31]), .D(n25242), .Y(
        n25240) );
  OAI21X1 U20648 ( .A(n25038), .B(n25244), .C(n25245), .Y(n25236) );
  AOI22X1 U20649 ( .A(reg_A[26]), .B(n25246), .C(reg_A[25]), .D(n25247), .Y(
        n25245) );
  NOR2X1 U20650 ( .A(n25248), .B(n25249), .Y(n25212) );
  OAI21X1 U20651 ( .A(n25030), .B(n25250), .C(n25251), .Y(n25249) );
  AOI22X1 U20652 ( .A(reg_A[11]), .B(n25252), .C(reg_A[15]), .D(n25253), .Y(
        n25251) );
  OAI21X1 U20653 ( .A(n25041), .B(n25255), .C(n25256), .Y(n25248) );
  AOI22X1 U20654 ( .A(reg_A[30]), .B(n25257), .C(reg_A[10]), .D(n25135), .Y(
        n25256) );
  AOI21X1 U20655 ( .A(n25258), .B(n25259), .C(n25260), .Y(n25199) );
  OAI22X1 U20656 ( .A(n25261), .B(n25262), .C(n25263), .D(n25264), .Y(n25260)
         );
  NAND3X1 U20657 ( .A(n25265), .B(n25266), .C(n25267), .Y(result[99]) );
  NOR2X1 U20658 ( .A(n25268), .B(n25269), .Y(n25267) );
  OR2X1 U20659 ( .A(n25270), .B(n25271), .Y(n25269) );
  OAI21X1 U20660 ( .A(n25272), .B(n25273), .C(n25274), .Y(n25271) );
  AOI22X1 U20661 ( .A(n25275), .B(n25276), .C(n25277), .D(n25278), .Y(n25274)
         );
  OAI21X1 U20662 ( .A(n25279), .B(n25280), .C(n25281), .Y(n25270) );
  AOI22X1 U20663 ( .A(reg_A[100]), .B(n25282), .C(reg_A[99]), .D(n25283), .Y(
        n25281) );
  AOI21X1 U20664 ( .A(reg_A[99]), .B(n25284), .C(n25285), .Y(n25280) );
  OAI22X1 U20665 ( .A(n25286), .B(n25287), .C(n25288), .D(n25289), .Y(n25285)
         );
  NAND3X1 U20666 ( .A(n25290), .B(n25291), .C(n25292), .Y(n25268) );
  AOI21X1 U20667 ( .A(reg_A[106]), .B(n25293), .C(n25294), .Y(n25292) );
  OAI22X1 U20668 ( .A(n25295), .B(n25296), .C(n25297), .D(n25298), .Y(n25294)
         );
  AOI22X1 U20669 ( .A(reg_A[109]), .B(n25299), .C(reg_A[110]), .D(n25300), .Y(
        n25291) );
  AOI22X1 U20670 ( .A(reg_A[108]), .B(n25301), .C(reg_A[107]), .D(n25302), .Y(
        n25290) );
  NOR2X1 U20671 ( .A(n25303), .B(n25304), .Y(n25266) );
  NAND3X1 U20672 ( .A(n25305), .B(n25306), .C(n25307), .Y(n25304) );
  OAI21X1 U20673 ( .A(n25308), .B(n25309), .C(n25310), .Y(n25307) );
  NAND3X1 U20674 ( .A(n25311), .B(n25312), .C(n25313), .Y(n25309) );
  NOR2X1 U20675 ( .A(n25314), .B(n25315), .Y(n25313) );
  OAI22X1 U20676 ( .A(n25316), .B(n25317), .C(n25318), .D(n25319), .Y(n25315)
         );
  OAI22X1 U20677 ( .A(n25057), .B(n25321), .C(n25322), .D(n25323), .Y(n25314)
         );
  AOI22X1 U20678 ( .A(reg_A[127]), .B(n25324), .C(reg_A[113]), .D(n25234), .Y(
        n25312) );
  AOI22X1 U20679 ( .A(reg_A[114]), .B(n25235), .C(reg_A[112]), .D(n25325), .Y(
        n25311) );
  NAND3X1 U20680 ( .A(n25326), .B(n25327), .C(n25328), .Y(n25308) );
  NOR2X1 U20681 ( .A(n25329), .B(n25330), .Y(n25328) );
  OAI22X1 U20682 ( .A(n25331), .B(n25332), .C(n25243), .D(n25333), .Y(n25330)
         );
  OAI22X1 U20683 ( .A(n25334), .B(n25335), .C(n25336), .D(n25337), .Y(n25329)
         );
  AOI22X1 U20684 ( .A(reg_A[121]), .B(n25242), .C(reg_A[122]), .D(n25338), .Y(
        n25327) );
  AOI22X1 U20685 ( .A(reg_A[119]), .B(n25339), .C(reg_A[120]), .D(n25257), .Y(
        n25326) );
  OAI21X1 U20686 ( .A(n25340), .B(n25341), .C(reg_A[96]), .Y(n25306) );
  OAI21X1 U20687 ( .A(n25031), .B(n25343), .C(n25344), .Y(n25341) );
  NAND2X1 U20688 ( .A(n25345), .B(n25346), .Y(n25305) );
  NAND3X1 U20689 ( .A(n25347), .B(n25348), .C(n25349), .Y(n25303) );
  AOI22X1 U20690 ( .A(n25350), .B(n25351), .C(n25352), .D(n25353), .Y(n25349)
         );
  INVX1 U20691 ( .A(n25354), .Y(n25351) );
  OAI21X1 U20692 ( .A(n25355), .B(n25356), .C(n25357), .Y(n25347) );
  NOR2X1 U20693 ( .A(n25358), .B(n25359), .Y(n25265) );
  OAI21X1 U20694 ( .A(n25360), .B(n25361), .C(n25362), .Y(n25359) );
  AOI22X1 U20695 ( .A(reg_A[111]), .B(n25363), .C(reg_A[101]), .D(n25364), .Y(
        n25362) );
  NAND3X1 U20696 ( .A(n25365), .B(n25366), .C(n25367), .Y(n25358) );
  AOI22X1 U20697 ( .A(reg_A[103]), .B(n25368), .C(reg_A[80]), .D(n25369), .Y(
        n25367) );
  OAI21X1 U20698 ( .A(n25370), .B(n25371), .C(n25372), .Y(n25366) );
  OAI22X1 U20699 ( .A(n25272), .B(n25373), .C(n25374), .D(n25375), .Y(n25371)
         );
  INVX1 U20700 ( .A(n25376), .Y(n25272) );
  OAI21X1 U20701 ( .A(n25377), .B(n25289), .C(n25378), .Y(n25370) );
  NAND3X1 U20702 ( .A(reg_B[102]), .B(reg_A[96]), .C(n25379), .Y(n25378) );
  OAI21X1 U20703 ( .A(n25380), .B(n25381), .C(n25382), .Y(n25365) );
  NAND2X1 U20704 ( .A(n25383), .B(n25384), .Y(n25381) );
  AOI22X1 U20705 ( .A(reg_A[101]), .B(n25385), .C(reg_A[99]), .D(n25386), .Y(
        n25384) );
  AOI22X1 U20706 ( .A(reg_A[102]), .B(n25387), .C(n25388), .D(n25389), .Y(
        n25383) );
  NAND3X1 U20707 ( .A(n25390), .B(n25391), .C(n25392), .Y(n25380) );
  AOI22X1 U20708 ( .A(n25393), .B(n25394), .C(reg_A[100]), .D(n25395), .Y(
        n25392) );
  OAI21X1 U20709 ( .A(n25396), .B(n25397), .C(n25398), .Y(n25394) );
  AOI22X1 U20710 ( .A(reg_A[102]), .B(n25355), .C(reg_A[101]), .D(n25399), .Y(
        n25398) );
  INVX1 U20711 ( .A(n25400), .Y(n25391) );
  AOI21X1 U20712 ( .A(n25401), .B(n25402), .C(n25403), .Y(n25400) );
  AOI22X1 U20713 ( .A(n25404), .B(n25405), .C(n25406), .D(n25407), .Y(n25402)
         );
  AOI22X1 U20714 ( .A(n25408), .B(n25409), .C(n25410), .D(reg_B[123]), .Y(
        n25401) );
  AOI22X1 U20715 ( .A(n25411), .B(reg_B[108]), .C(n25412), .D(reg_A[103]), .Y(
        n25390) );
  NOR2X1 U20716 ( .A(n25373), .B(n25413), .Y(n25412) );
  NOR2X1 U20717 ( .A(n25414), .B(n25415), .Y(n25411) );
  NAND3X1 U20718 ( .A(n25416), .B(n25417), .C(n25418), .Y(result[98]) );
  NOR2X1 U20719 ( .A(n25419), .B(n25420), .Y(n25418) );
  NAND3X1 U20720 ( .A(n25421), .B(n25422), .C(n25423), .Y(n25420) );
  AOI22X1 U20721 ( .A(n25357), .B(reg_B[126]), .C(n25277), .D(n25276), .Y(
        n25423) );
  OAI21X1 U20722 ( .A(n25424), .B(n25425), .C(n25426), .Y(n25276) );
  NAND3X1 U20723 ( .A(n25427), .B(n25428), .C(reg_A[98]), .Y(n25426) );
  OAI21X1 U20724 ( .A(n25429), .B(n25430), .C(n25203), .Y(n25422) );
  NAND3X1 U20725 ( .A(n25431), .B(n25432), .C(n25433), .Y(n25430) );
  AOI21X1 U20726 ( .A(reg_A[98]), .B(n25434), .C(n25435), .Y(n25433) );
  OAI22X1 U20727 ( .A(n25436), .B(n25437), .C(n25361), .D(n25438), .Y(n25435)
         );
  AOI22X1 U20728 ( .A(n25439), .B(reg_A[108]), .C(n25440), .D(reg_A[104]), .Y(
        n25432) );
  AOI22X1 U20729 ( .A(reg_A[99]), .B(n25441), .C(n25442), .D(reg_A[101]), .Y(
        n25431) );
  NAND3X1 U20730 ( .A(n25443), .B(n25444), .C(n25445), .Y(n25429) );
  NOR2X1 U20731 ( .A(n25446), .B(n25447), .Y(n25445) );
  OAI22X1 U20732 ( .A(n25448), .B(n25449), .C(n25450), .D(n25451), .Y(n25447)
         );
  OAI21X1 U20733 ( .A(n25452), .B(n25453), .C(n25454), .Y(n25446) );
  OAI21X1 U20734 ( .A(n25455), .B(n25456), .C(n25044), .Y(n25454) );
  NAND3X1 U20735 ( .A(n25457), .B(n25458), .C(n25459), .Y(n25456) );
  NOR2X1 U20736 ( .A(n25460), .B(n25461), .Y(n25459) );
  OAI21X1 U20737 ( .A(n25043), .B(n25289), .C(n25462), .Y(n25461) );
  AOI22X1 U20738 ( .A(reg_A[99]), .B(n25135), .C(reg_A[100]), .D(n25252), .Y(
        n25462) );
  NAND2X1 U20739 ( .A(n25463), .B(n25464), .Y(n25460) );
  AOI22X1 U20740 ( .A(reg_A[101]), .B(n25136), .C(reg_A[104]), .D(n25253), .Y(
        n25464) );
  AOI22X1 U20741 ( .A(reg_A[102]), .B(n25070), .C(reg_A[103]), .D(n25123), .Y(
        n25463) );
  NOR2X1 U20742 ( .A(n25465), .B(n25466), .Y(n25458) );
  OAI22X1 U20743 ( .A(n25034), .B(n25468), .C(n25129), .D(n25296), .Y(n25466)
         );
  OAI22X1 U20744 ( .A(n25036), .B(n25469), .C(n25037), .D(n25470), .Y(n25465)
         );
  NOR2X1 U20745 ( .A(n25471), .B(n25472), .Y(n25457) );
  OAI22X1 U20746 ( .A(n25064), .B(n25450), .C(n25473), .D(n25474), .Y(n25472)
         );
  OAI22X1 U20747 ( .A(n25039), .B(n25452), .C(n25035), .D(n25476), .Y(n25471)
         );
  NAND3X1 U20748 ( .A(n25477), .B(n25478), .C(n25479), .Y(n25455) );
  NOR2X1 U20749 ( .A(n25480), .B(n25481), .Y(n25479) );
  OAI21X1 U20750 ( .A(n25065), .B(n25483), .C(n25484), .Y(n25481) );
  AOI22X1 U20751 ( .A(reg_A[115]), .B(n25246), .C(reg_A[114]), .D(n25247), .Y(
        n25484) );
  NAND2X1 U20752 ( .A(n25485), .B(n25486), .Y(n25480) );
  AOI22X1 U20753 ( .A(reg_A[117]), .B(n25487), .C(reg_A[116]), .D(n25241), .Y(
        n25486) );
  AOI22X1 U20754 ( .A(reg_A[118]), .B(n25339), .C(reg_A[119]), .D(n25257), .Y(
        n25485) );
  NOR2X1 U20755 ( .A(n25488), .B(n25489), .Y(n25478) );
  OAI22X1 U20756 ( .A(n25490), .B(n25491), .C(n25492), .D(n25493), .Y(n25489)
         );
  OAI22X1 U20757 ( .A(n25494), .B(n25320), .C(n25322), .D(n25321), .Y(n25488)
         );
  NOR2X1 U20758 ( .A(n25495), .B(n25496), .Y(n25477) );
  OAI22X1 U20759 ( .A(n25323), .B(n25316), .C(n25318), .D(n25317), .Y(n25496)
         );
  OAI22X1 U20760 ( .A(n25497), .B(n25498), .C(n25319), .D(n25499), .Y(n25495)
         );
  AOI22X1 U20761 ( .A(n25500), .B(reg_A[107]), .C(n25501), .D(reg_A[106]), .Y(
        n25444) );
  AOI22X1 U20762 ( .A(n25502), .B(reg_A[105]), .C(n25503), .D(reg_A[109]), .Y(
        n25443) );
  NAND2X1 U20763 ( .A(n25504), .B(n25505), .Y(n25419) );
  AOI22X1 U20764 ( .A(n25506), .B(reg_A[100]), .C(n25507), .D(reg_A[101]), .Y(
        n25505) );
  AOI22X1 U20765 ( .A(n25508), .B(reg_A[102]), .C(n25509), .D(reg_A[103]), .Y(
        n25504) );
  NOR2X1 U20766 ( .A(n25510), .B(n25511), .Y(n25417) );
  OAI21X1 U20767 ( .A(n25512), .B(n25513), .C(n25514), .Y(n25511) );
  NAND2X1 U20768 ( .A(reg_A[98]), .B(n25515), .Y(n25514) );
  OAI21X1 U20769 ( .A(n25516), .B(n25517), .C(n25518), .Y(n25515) );
  INVX1 U20770 ( .A(n25353), .Y(n25512) );
  OAI21X1 U20771 ( .A(n25424), .B(n25519), .C(n25520), .Y(n25353) );
  NAND3X1 U20772 ( .A(reg_A[98]), .B(n25521), .C(n25522), .Y(n25520) );
  OAI21X1 U20773 ( .A(n25523), .B(n25524), .C(n25348), .Y(n25510) );
  OR2X1 U20774 ( .A(n25525), .B(n25343), .Y(n25524) );
  NOR2X1 U20775 ( .A(n25526), .B(n25527), .Y(n25416) );
  OAI21X1 U20776 ( .A(n25528), .B(n25424), .C(n25529), .Y(n25527) );
  OAI21X1 U20777 ( .A(n25530), .B(n25531), .C(n25382), .Y(n25529) );
  NAND2X1 U20778 ( .A(n25532), .B(n25533), .Y(n25531) );
  AOI22X1 U20779 ( .A(reg_A[100]), .B(n25385), .C(reg_A[98]), .D(n25386), .Y(
        n25533) );
  AOI22X1 U20780 ( .A(reg_A[101]), .B(n25387), .C(n25534), .D(n25535), .Y(
        n25532) );
  NAND3X1 U20781 ( .A(n25536), .B(n25537), .C(n25538), .Y(n25530) );
  AOI22X1 U20782 ( .A(n25393), .B(n25539), .C(reg_A[99]), .D(n25395), .Y(
        n25538) );
  OAI21X1 U20783 ( .A(n25289), .B(n25397), .C(n25540), .Y(n25539) );
  AOI22X1 U20784 ( .A(reg_A[101]), .B(n25355), .C(reg_A[100]), .D(n25399), .Y(
        n25540) );
  OAI21X1 U20785 ( .A(n25541), .B(n25542), .C(n25044), .Y(n25537) );
  OAI22X1 U20786 ( .A(n25543), .B(n25544), .C(n25545), .D(n25546), .Y(n25542)
         );
  INVX1 U20787 ( .A(n25547), .Y(n25543) );
  OAI22X1 U20788 ( .A(n25548), .B(n25549), .C(n25550), .D(n25551), .Y(n25541)
         );
  INVX1 U20789 ( .A(n25552), .Y(n25548) );
  AOI21X1 U20790 ( .A(n25553), .B(n25554), .C(n25555), .Y(n25536) );
  AOI21X1 U20791 ( .A(n25556), .B(n25557), .C(n25558), .Y(n25555) );
  AOI22X1 U20792 ( .A(reg_A[103]), .B(n25559), .C(reg_A[105]), .D(n25560), .Y(
        n25557) );
  AOI22X1 U20793 ( .A(reg_A[102]), .B(n25561), .C(reg_A[104]), .D(n25562), .Y(
        n25556) );
  OAI21X1 U20794 ( .A(n25354), .B(n25273), .C(n25563), .Y(n25526) );
  OAI21X1 U20795 ( .A(n25564), .B(n25565), .C(reg_A[97]), .Y(n25563) );
  OAI21X1 U20796 ( .A(n25377), .B(n25517), .C(n25566), .Y(n25565) );
  INVX1 U20797 ( .A(n25567), .Y(n25377) );
  OAI21X1 U20798 ( .A(n25568), .B(n25569), .C(n25570), .Y(n25567) );
  AOI21X1 U20799 ( .A(n25571), .B(n25572), .C(n25573), .Y(n25570) );
  AOI22X1 U20800 ( .A(n25574), .B(reg_A[98]), .C(reg_A[96]), .D(n25575), .Y(
        n25354) );
  NAND3X1 U20801 ( .A(n25576), .B(n25577), .C(n25578), .Y(result[97]) );
  NOR2X1 U20802 ( .A(n25579), .B(n25580), .Y(n25578) );
  NAND2X1 U20803 ( .A(n25581), .B(n25421), .Y(n25580) );
  INVX1 U20804 ( .A(n25582), .Y(n25421) );
  OAI21X1 U20805 ( .A(n25583), .B(n25584), .C(n25585), .Y(n25582) );
  NAND3X1 U20806 ( .A(n25372), .B(n25586), .C(reg_A[96]), .Y(n25585) );
  OAI21X1 U20807 ( .A(n25427), .B(n25403), .C(n25587), .Y(n25586) );
  AOI22X1 U20808 ( .A(n25588), .B(reg_B[110]), .C(n25589), .D(n25590), .Y(
        n25587) );
  NOR2X1 U20809 ( .A(n25415), .B(n25591), .Y(n25588) );
  AOI22X1 U20810 ( .A(n25357), .B(n25397), .C(n25203), .D(n25592), .Y(n25581)
         );
  NAND3X1 U20811 ( .A(n25593), .B(n25594), .C(n25595), .Y(n25592) );
  NOR2X1 U20812 ( .A(n25596), .B(n25597), .Y(n25595) );
  OAI22X1 U20813 ( .A(n25598), .B(n25396), .C(n25599), .D(n25436), .Y(n25597)
         );
  OAI21X1 U20814 ( .A(n25600), .B(n25361), .C(n25601), .Y(n25596) );
  OAI21X1 U20815 ( .A(n25602), .B(n25603), .C(n25604), .Y(n25601) );
  NAND2X1 U20816 ( .A(n25605), .B(n25606), .Y(n25603) );
  AOI22X1 U20817 ( .A(reg_A[107]), .B(n25607), .C(reg_A[111]), .D(n25608), .Y(
        n25606) );
  AOI22X1 U20818 ( .A(reg_A[109]), .B(n25609), .C(reg_A[110]), .D(n25610), .Y(
        n25605) );
  NAND2X1 U20819 ( .A(n25611), .B(n25612), .Y(n25602) );
  AOI22X1 U20820 ( .A(reg_A[104]), .B(n25613), .C(reg_A[106]), .D(n25614), .Y(
        n25612) );
  AOI22X1 U20821 ( .A(reg_A[105]), .B(n25615), .C(reg_A[108]), .D(n25616), .Y(
        n25611) );
  AOI21X1 U20822 ( .A(reg_A[98]), .B(n25617), .C(n25618), .Y(n25594) );
  OAI21X1 U20823 ( .A(n25619), .B(n25287), .C(n25620), .Y(n25618) );
  OAI21X1 U20824 ( .A(n25621), .B(n25622), .C(n25044), .Y(n25620) );
  NAND2X1 U20825 ( .A(n25623), .B(n25624), .Y(n25622) );
  NOR2X1 U20826 ( .A(n25625), .B(n25626), .Y(n25624) );
  OAI21X1 U20827 ( .A(n25034), .B(n25296), .C(n25627), .Y(n25626) );
  AOI22X1 U20828 ( .A(reg_A[104]), .B(n25628), .C(reg_A[106]), .D(n25629), .Y(
        n25627) );
  OAI21X1 U20829 ( .A(n25319), .B(n25498), .C(n25630), .Y(n25625) );
  AOI22X1 U20830 ( .A(n25631), .B(reg_A[127]), .C(n25324), .D(reg_A[125]), .Y(
        n25630) );
  NOR2X1 U20831 ( .A(n25632), .B(n25633), .Y(n25623) );
  OAI21X1 U20832 ( .A(n25039), .B(n25450), .C(n25634), .Y(n25633) );
  AOI22X1 U20833 ( .A(reg_A[112]), .B(n25235), .C(reg_A[109]), .D(n25635), .Y(
        n25634) );
  OAI21X1 U20834 ( .A(n25035), .B(n25452), .C(n25636), .Y(n25632) );
  AOI22X1 U20835 ( .A(reg_A[108]), .B(n25222), .C(reg_A[107]), .D(n25637), .Y(
        n25636) );
  NAND2X1 U20836 ( .A(n25638), .B(n25639), .Y(n25621) );
  NOR2X1 U20837 ( .A(n25640), .B(n25641), .Y(n25639) );
  OAI21X1 U20838 ( .A(n25050), .B(n25493), .C(n25642), .Y(n25641) );
  AOI22X1 U20839 ( .A(reg_A[115]), .B(n25241), .C(reg_A[119]), .D(n25242), .Y(
        n25642) );
  OAI21X1 U20840 ( .A(n25038), .B(n25337), .C(n25643), .Y(n25640) );
  AOI22X1 U20841 ( .A(reg_A[114]), .B(n25246), .C(reg_A[113]), .D(n25247), .Y(
        n25643) );
  NOR2X1 U20842 ( .A(n25644), .B(n25645), .Y(n25638) );
  OAI21X1 U20843 ( .A(n25321), .B(n25316), .C(n25646), .Y(n25645) );
  AOI22X1 U20844 ( .A(n25647), .B(reg_A[121]), .C(n25648), .D(reg_A[124]), .Y(
        n25646) );
  OAI21X1 U20845 ( .A(n25494), .B(n25322), .C(n25649), .Y(n25644) );
  AOI22X1 U20846 ( .A(reg_A[117]), .B(n25339), .C(reg_A[118]), .D(n25257), .Y(
        n25649) );
  AOI22X1 U20847 ( .A(reg_A[101]), .B(n25650), .C(reg_A[103]), .D(n25651), .Y(
        n25593) );
  OAI21X1 U20848 ( .A(n25361), .B(n25652), .C(n25653), .Y(n25579) );
  AOI22X1 U20849 ( .A(n25507), .B(reg_A[100]), .C(n25508), .D(reg_A[101]), .Y(
        n25653) );
  AOI21X1 U20850 ( .A(reg_A[96]), .B(n25654), .C(n25655), .Y(n25577) );
  OAI21X1 U20851 ( .A(n25656), .B(n25657), .C(n25658), .Y(n25655) );
  OAI21X1 U20852 ( .A(n25659), .B(n25660), .C(n25382), .Y(n25658) );
  NAND2X1 U20853 ( .A(n25661), .B(n25662), .Y(n25660) );
  AOI21X1 U20854 ( .A(reg_A[97]), .B(n25386), .C(n25663), .Y(n25662) );
  OAI21X1 U20855 ( .A(n25664), .B(n25396), .C(n25665), .Y(n25663) );
  OAI21X1 U20856 ( .A(n25666), .B(n25667), .C(n25388), .Y(n25665) );
  OAI22X1 U20857 ( .A(n25668), .B(n25448), .C(n25669), .D(n25670), .Y(n25667)
         );
  OAI22X1 U20858 ( .A(n25671), .B(n25298), .C(n25672), .D(n25361), .Y(n25666)
         );
  AOI22X1 U20859 ( .A(reg_A[100]), .B(n25387), .C(n25534), .D(n25673), .Y(
        n25661) );
  INVX1 U20860 ( .A(n25674), .Y(n25534) );
  INVX1 U20861 ( .A(n25675), .Y(n25387) );
  NAND3X1 U20862 ( .A(n25676), .B(n25677), .C(n25678), .Y(n25659) );
  AOI22X1 U20863 ( .A(n25393), .B(n25679), .C(reg_A[98]), .D(n25395), .Y(
        n25678) );
  OAI21X1 U20864 ( .A(n25568), .B(n25569), .C(n25680), .Y(n25395) );
  OAI21X1 U20865 ( .A(n25287), .B(n25397), .C(n25681), .Y(n25679) );
  AOI22X1 U20866 ( .A(reg_A[100]), .B(n25355), .C(n25399), .D(reg_A[99]), .Y(
        n25681) );
  INVX1 U20867 ( .A(n25682), .Y(n25677) );
  AOI21X1 U20868 ( .A(n25683), .B(n25684), .C(n25403), .Y(n25682) );
  AOI22X1 U20869 ( .A(n25685), .B(n25405), .C(n25686), .D(n25407), .Y(n25684)
         );
  AOI22X1 U20870 ( .A(n25687), .B(n25409), .C(n25688), .D(reg_B[123]), .Y(
        n25683) );
  AOI22X1 U20871 ( .A(n25553), .B(n25689), .C(n25690), .D(n25691), .Y(n25676)
         );
  NAND2X1 U20872 ( .A(n25692), .B(n25372), .Y(n25657) );
  NAND3X1 U20873 ( .A(n25693), .B(n25694), .C(n25695), .Y(n25654) );
  AOI21X1 U20874 ( .A(n25379), .B(n25372), .C(n25696), .Y(n25695) );
  INVX1 U20875 ( .A(n25564), .Y(n25694) );
  OAI21X1 U20876 ( .A(n25680), .B(n25697), .C(n25698), .Y(n25564) );
  NAND3X1 U20877 ( .A(n25427), .B(n25699), .C(n25700), .Y(n25698) );
  AOI21X1 U20878 ( .A(n25506), .B(reg_A[99]), .C(n25701), .Y(n25576) );
  OAI21X1 U20879 ( .A(n25448), .B(n25702), .C(n25703), .Y(n25701) );
  OAI21X1 U20880 ( .A(n25704), .B(n25705), .C(reg_A[97]), .Y(n25703) );
  OAI21X1 U20881 ( .A(n25516), .B(n25517), .C(n25706), .Y(n25705) );
  INVX1 U20882 ( .A(n25707), .Y(n25516) );
  OAI21X1 U20883 ( .A(n25569), .B(n25397), .C(n25708), .Y(n25707) );
  AOI21X1 U20884 ( .A(n25709), .B(n25571), .C(n25710), .Y(n25708) );
  INVX1 U20885 ( .A(n25711), .Y(n25710) );
  NAND3X1 U20886 ( .A(n25712), .B(n25713), .C(n25714), .Y(result[96]) );
  NOR2X1 U20887 ( .A(n25715), .B(n25716), .Y(n25714) );
  OAI22X1 U20888 ( .A(n25289), .B(n25717), .C(n25396), .D(n25718), .Y(n25716)
         );
  OAI21X1 U20889 ( .A(n25287), .B(n25719), .C(n25720), .Y(n25715) );
  AOI22X1 U20890 ( .A(n25721), .B(reg_A[80]), .C(n25722), .D(reg_A[100]), .Y(
        n25720) );
  AOI21X1 U20891 ( .A(n25310), .B(n25723), .C(n25724), .Y(n25713) );
  OAI21X1 U20892 ( .A(n25725), .B(n25726), .C(n25727), .Y(n25724) );
  OAI21X1 U20893 ( .A(n25728), .B(n25729), .C(n25730), .Y(n25727) );
  NAND3X1 U20894 ( .A(n25731), .B(n25732), .C(n25733), .Y(n25729) );
  NOR2X1 U20895 ( .A(n25734), .B(n25735), .Y(n25733) );
  OAI22X1 U20896 ( .A(n25736), .B(n25424), .C(n25737), .D(n25474), .Y(n25735)
         );
  OAI22X1 U20897 ( .A(n25738), .B(n25469), .C(n25739), .D(n25452), .Y(n25734)
         );
  AOI22X1 U20898 ( .A(reg_A[104]), .B(n25615), .C(reg_A[107]), .D(n25616), .Y(
        n25732) );
  AOI22X1 U20899 ( .A(reg_A[106]), .B(n25607), .C(reg_A[110]), .D(n25608), .Y(
        n25731) );
  NAND3X1 U20900 ( .A(n25740), .B(n25741), .C(n25742), .Y(n25728) );
  NOR2X1 U20901 ( .A(n25743), .B(n25744), .Y(n25742) );
  OAI22X1 U20902 ( .A(n25061), .B(n25361), .C(n25746), .D(n25289), .Y(n25744)
         );
  OAI22X1 U20903 ( .A(n25747), .B(n25396), .C(n25748), .D(n25287), .Y(n25743)
         );
  AOI22X1 U20904 ( .A(reg_A[103]), .B(n25613), .C(reg_A[100]), .D(n25749), .Y(
        n25741) );
  AOI22X1 U20905 ( .A(reg_A[101]), .B(n25750), .C(reg_A[105]), .D(n25614), .Y(
        n25740) );
  AOI21X1 U20906 ( .A(reg_A[101]), .B(n25751), .C(n25752), .Y(n25725) );
  OAI22X1 U20907 ( .A(n25753), .B(n25448), .C(n25754), .D(n25361), .Y(n25752)
         );
  NAND2X1 U20908 ( .A(n25755), .B(n25756), .Y(n25723) );
  NOR2X1 U20909 ( .A(n25757), .B(n25758), .Y(n25756) );
  NAND3X1 U20910 ( .A(n25759), .B(n25760), .C(n25761), .Y(n25758) );
  NOR2X1 U20911 ( .A(n25762), .B(n25763), .Y(n25761) );
  OAI22X1 U20912 ( .A(n25494), .B(n25316), .C(n25321), .D(n25318), .Y(n25763)
         );
  OAI22X1 U20913 ( .A(n25493), .B(n25320), .C(n25490), .D(n25322), .Y(n25762)
         );
  AOI22X1 U20914 ( .A(n25631), .B(reg_A[126]), .C(n25764), .D(reg_A[127]), .Y(
        n25760) );
  AOI22X1 U20915 ( .A(n25324), .B(reg_A[124]), .C(n25765), .D(reg_A[125]), .Y(
        n25759) );
  NAND3X1 U20916 ( .A(n25766), .B(n25767), .C(n25768), .Y(n25757) );
  NOR2X1 U20917 ( .A(n25769), .B(n25770), .Y(n25768) );
  OAI22X1 U20918 ( .A(n25051), .B(n25771), .C(n25243), .D(n25335), .Y(n25770)
         );
  OAI22X1 U20919 ( .A(n25048), .B(n25476), .C(n25336), .D(n25483), .Y(n25769)
         );
  AOI22X1 U20920 ( .A(reg_A[118]), .B(n25242), .C(reg_A[119]), .D(n25338), .Y(
        n25767) );
  AOI22X1 U20921 ( .A(reg_A[116]), .B(n25339), .C(reg_A[117]), .D(n25257), .Y(
        n25766) );
  NOR2X1 U20922 ( .A(n25772), .B(n25773), .Y(n25755) );
  NAND3X1 U20923 ( .A(n25774), .B(n25775), .C(n25776), .Y(n25773) );
  NOR2X1 U20924 ( .A(n25777), .B(n25778), .Y(n25776) );
  OAI22X1 U20925 ( .A(n25043), .B(n25424), .C(n25039), .D(n25474), .Y(n25778)
         );
  OAI22X1 U20926 ( .A(n25064), .B(n25469), .C(n25065), .D(n25452), .Y(n25777)
         );
  AOI22X1 U20927 ( .A(reg_A[104]), .B(n25124), .C(reg_A[107]), .D(n25222), .Y(
        n25775) );
  AOI22X1 U20928 ( .A(reg_A[106]), .B(n25637), .C(reg_A[110]), .D(n25234), .Y(
        n25774) );
  NAND3X1 U20929 ( .A(n25779), .B(n25780), .C(n25781), .Y(n25772) );
  NOR2X1 U20930 ( .A(n25782), .B(n25783), .Y(n25781) );
  OAI22X1 U20931 ( .A(n25033), .B(n25361), .C(n25040), .D(n25289), .Y(n25783)
         );
  OAI22X1 U20932 ( .A(n25041), .B(n25396), .C(n25042), .D(n25287), .Y(n25782)
         );
  AOI22X1 U20933 ( .A(reg_A[103]), .B(n25628), .C(reg_A[100]), .D(n25066), .Y(
        n25780) );
  AOI22X1 U20934 ( .A(reg_A[101]), .B(n25123), .C(reg_A[105]), .D(n25629), .Y(
        n25779) );
  AND2X1 U20935 ( .A(n25785), .B(n25786), .Y(n25712) );
  OAI21X1 U20936 ( .A(n25787), .B(n25788), .C(reg_A[96]), .Y(n25786) );
  NAND2X1 U20937 ( .A(n25789), .B(n25790), .Y(n25788) );
  INVX1 U20938 ( .A(n25704), .Y(n25790) );
  OAI21X1 U20939 ( .A(n25791), .B(n25697), .C(n25792), .Y(n25704) );
  NAND3X1 U20940 ( .A(n25427), .B(n25699), .C(n25793), .Y(n25792) );
  INVX1 U20941 ( .A(n25386), .Y(n25791) );
  OAI21X1 U20942 ( .A(n25032), .B(n25591), .C(n25795), .Y(n25787) );
  OAI21X1 U20943 ( .A(n25796), .B(n25797), .C(n25382), .Y(n25785) );
  OR2X1 U20944 ( .A(n25798), .B(n25799), .Y(n25797) );
  OAI22X1 U20945 ( .A(n25800), .B(n25674), .C(n25680), .D(n25287), .Y(n25799)
         );
  NOR2X1 U20946 ( .A(n25801), .B(n25573), .Y(n25680) );
  NOR2X1 U20947 ( .A(n25802), .B(n25590), .Y(n25573) );
  INVX1 U20948 ( .A(n25803), .Y(n25800) );
  OAI21X1 U20949 ( .A(n25675), .B(n25396), .C(n25804), .Y(n25798) );
  OAI21X1 U20950 ( .A(n25805), .B(n25806), .C(n25044), .Y(n25804) );
  OAI22X1 U20951 ( .A(n25807), .B(n25544), .C(n25808), .D(n25546), .Y(n25806)
         );
  INVX1 U20952 ( .A(n25809), .Y(n25807) );
  OAI21X1 U20953 ( .A(n25810), .B(n25549), .C(n25811), .Y(n25805) );
  AOI22X1 U20954 ( .A(n25427), .B(n25812), .C(reg_B[123]), .D(n25813), .Y(
        n25811) );
  NAND2X1 U20955 ( .A(n25814), .B(n25815), .Y(n25812) );
  AOI22X1 U20956 ( .A(n25355), .B(reg_A[99]), .C(n25399), .D(reg_A[98]), .Y(
        n25815) );
  AOI22X1 U20957 ( .A(n25793), .B(reg_A[96]), .C(n25700), .D(reg_A[97]), .Y(
        n25814) );
  AOI21X1 U20958 ( .A(n25575), .B(n25379), .C(n25816), .Y(n25675) );
  NAND3X1 U20959 ( .A(n25817), .B(n25818), .C(n25819), .Y(n25796) );
  AOI22X1 U20960 ( .A(reg_A[98]), .B(n25385), .C(reg_A[96]), .D(n25386), .Y(
        n25819) );
  OAI21X1 U20961 ( .A(n25820), .B(n25656), .C(n25711), .Y(n25386) );
  INVX1 U20962 ( .A(n25664), .Y(n25385) );
  NOR2X1 U20963 ( .A(n25821), .B(n25822), .Y(n25664) );
  OAI21X1 U20964 ( .A(n25823), .B(n25824), .C(n25388), .Y(n25818) );
  OAI22X1 U20965 ( .A(n25668), .B(n25361), .C(n25669), .D(n25436), .Y(n25824)
         );
  OAI22X1 U20966 ( .A(n25671), .B(n25448), .C(n25672), .D(n25670), .Y(n25823)
         );
  AOI22X1 U20967 ( .A(n25553), .B(n25825), .C(n25690), .D(n25826), .Y(n25817)
         );
  NOR2X1 U20968 ( .A(n25827), .B(n25415), .Y(n25553) );
  NAND3X1 U20969 ( .A(n25828), .B(n25829), .C(n25830), .Y(result[95]) );
  NOR2X1 U20970 ( .A(n25831), .B(n25832), .Y(n25830) );
  OR2X1 U20971 ( .A(n25833), .B(n25834), .Y(n25832) );
  OAI21X1 U20972 ( .A(n25835), .B(n25836), .C(n25837), .Y(n25834) );
  AOI22X1 U20973 ( .A(n25838), .B(n25839), .C(n25840), .D(n25841), .Y(n25837)
         );
  NAND2X1 U20974 ( .A(n25842), .B(n25843), .Y(n25841) );
  NOR2X1 U20975 ( .A(n25844), .B(n25845), .Y(n25843) );
  NAND3X1 U20976 ( .A(n25846), .B(n25847), .C(n25848), .Y(n25845) );
  NOR2X1 U20977 ( .A(n25849), .B(n25850), .Y(n25848) );
  OAI22X1 U20978 ( .A(n25499), .B(n25851), .C(n25852), .D(n25853), .Y(n25850)
         );
  OAI22X1 U20979 ( .A(n25854), .B(n25855), .C(n25316), .D(n25856), .Y(n25849)
         );
  AOI22X1 U20980 ( .A(reg_A[74]), .B(n25257), .C(reg_A[70]), .D(n25857), .Y(
        n25847) );
  AOI22X1 U20981 ( .A(reg_A[71]), .B(n25647), .C(reg_A[68]), .D(n25648), .Y(
        n25846) );
  NAND3X1 U20982 ( .A(n25858), .B(n25859), .C(n25860), .Y(n25844) );
  NOR2X1 U20983 ( .A(n25861), .B(n25862), .Y(n25860) );
  OAI22X1 U20984 ( .A(n25038), .B(n25863), .C(n25334), .D(n25864), .Y(n25862)
         );
  OAI21X1 U20985 ( .A(n25047), .B(n25865), .C(n25836), .Y(n25861) );
  AOI22X1 U20986 ( .A(reg_A[77]), .B(n25241), .C(reg_A[73]), .D(n25242), .Y(
        n25859) );
  AOI22X1 U20987 ( .A(reg_A[72]), .B(n25338), .C(reg_A[75]), .D(n25339), .Y(
        n25858) );
  NOR2X1 U20988 ( .A(n25866), .B(n25867), .Y(n25842) );
  NAND3X1 U20989 ( .A(n25868), .B(n25869), .C(n25870), .Y(n25867) );
  NOR2X1 U20990 ( .A(n25871), .B(n25872), .Y(n25870) );
  OAI22X1 U20991 ( .A(n25043), .B(n25873), .C(n25039), .D(n25874), .Y(n25872)
         );
  OAI22X1 U20992 ( .A(n25064), .B(n25875), .C(n25482), .D(n25584), .Y(n25871)
         );
  AOI22X1 U20993 ( .A(reg_A[86]), .B(n25629), .C(reg_A[84]), .D(n25222), .Y(
        n25869) );
  AOI22X1 U20994 ( .A(reg_A[85]), .B(n25637), .C(reg_A[81]), .D(n25234), .Y(
        n25868) );
  NAND3X1 U20995 ( .A(n25876), .B(n25877), .C(n25878), .Y(n25866) );
  NOR2X1 U20996 ( .A(n25879), .B(n25880), .Y(n25878) );
  OAI22X1 U20997 ( .A(n25040), .B(n25881), .C(n25254), .D(n25882), .Y(n25880)
         );
  OAI22X1 U20998 ( .A(n25042), .B(n25883), .C(n25498), .D(n25884), .Y(n25879)
         );
  AOI22X1 U20999 ( .A(reg_A[89]), .B(n25253), .C(reg_A[88]), .D(n25628), .Y(
        n25877) );
  AOI22X1 U21000 ( .A(reg_A[91]), .B(n25070), .C(reg_A[90]), .D(n25123), .Y(
        n25876) );
  OAI21X1 U21001 ( .A(n25885), .B(n25886), .C(n25887), .Y(n25839) );
  AOI22X1 U21002 ( .A(n25888), .B(n25889), .C(n25890), .D(n25891), .Y(n25887)
         );
  OAI21X1 U21003 ( .A(reg_B[92]), .B(n25794), .C(n25031), .Y(n25889) );
  MUX2X1 U21004 ( .B(n25873), .A(n25883), .S(reg_B[95]), .Y(n25888) );
  AOI21X1 U21005 ( .A(reg_A[87]), .B(n25892), .C(n25893), .Y(n25885) );
  OAI22X1 U21006 ( .A(n25894), .B(n25873), .C(n25895), .D(n25896), .Y(n25893)
         );
  OAI21X1 U21007 ( .A(n25897), .B(n25898), .C(n25899), .Y(n25833) );
  AOI22X1 U21008 ( .A(n25900), .B(n25901), .C(n25902), .D(n25903), .Y(n25899)
         );
  AOI21X1 U21009 ( .A(n25904), .B(n25188), .C(n25905), .Y(n25897) );
  OAI22X1 U21010 ( .A(n25906), .B(n25886), .C(n25907), .D(n25342), .Y(n25905)
         );
  NAND2X1 U21011 ( .A(n25908), .B(n25909), .Y(n25831) );
  AOI21X1 U21012 ( .A(n25910), .B(n25911), .C(n25912), .Y(n25909) );
  OAI21X1 U21013 ( .A(n25913), .B(n25914), .C(n25915), .Y(n25912) );
  OAI21X1 U21014 ( .A(n25916), .B(n25917), .C(n25918), .Y(n25915) );
  NAND3X1 U21015 ( .A(n25919), .B(n25920), .C(n25921), .Y(n25917) );
  NOR2X1 U21016 ( .A(n25922), .B(n25923), .Y(n25921) );
  OAI22X1 U21017 ( .A(n25736), .B(n25873), .C(n25737), .D(n25874), .Y(n25923)
         );
  OAI22X1 U21018 ( .A(n25738), .B(n25875), .C(n25739), .D(n25584), .Y(n25922)
         );
  AOI22X1 U21019 ( .A(reg_A[87]), .B(n25615), .C(reg_A[84]), .D(n25616), .Y(
        n25920) );
  AOI22X1 U21020 ( .A(reg_A[85]), .B(n25607), .C(reg_A[81]), .D(n25608), .Y(
        n25919) );
  NAND3X1 U21021 ( .A(n25924), .B(n25925), .C(n25926), .Y(n25916) );
  NOR2X1 U21022 ( .A(n25927), .B(n25928), .Y(n25926) );
  OAI22X1 U21023 ( .A(n25061), .B(n25929), .C(n25746), .D(n25881), .Y(n25928)
         );
  OAI22X1 U21024 ( .A(n25747), .B(n25882), .C(n25748), .D(n25883), .Y(n25927)
         );
  AOI22X1 U21025 ( .A(reg_A[88]), .B(n25613), .C(reg_A[91]), .D(n25749), .Y(
        n25925) );
  AOI22X1 U21026 ( .A(reg_A[90]), .B(n25750), .C(reg_A[86]), .D(n25614), .Y(
        n25924) );
  AOI22X1 U21027 ( .A(n25699), .B(n25930), .C(n25931), .D(n25932), .Y(n25913)
         );
  INVX1 U21028 ( .A(n25933), .Y(n25931) );
  INVX1 U21029 ( .A(n25934), .Y(n25911) );
  AOI21X1 U21030 ( .A(n25935), .B(n25936), .C(n25937), .Y(n25908) );
  OAI22X1 U21031 ( .A(n25938), .B(n25939), .C(n25940), .D(n25941), .Y(n25937)
         );
  NOR2X1 U21032 ( .A(n25942), .B(n25943), .Y(n25829) );
  OAI21X1 U21033 ( .A(n25944), .B(n25945), .C(n25946), .Y(n25943) );
  AOI22X1 U21034 ( .A(n25947), .B(reg_A[90]), .C(n25948), .D(reg_A[91]), .Y(
        n25946) );
  OAI21X1 U21035 ( .A(n25949), .B(n25950), .C(n25951), .Y(n25942) );
  AOI21X1 U21036 ( .A(reg_A[95]), .B(n25952), .C(n25953), .Y(n25951) );
  AOI21X1 U21037 ( .A(n25954), .B(n25955), .C(n25697), .Y(n25953) );
  AOI21X1 U21038 ( .A(n25589), .B(n25956), .C(n25957), .Y(n25955) );
  OAI21X1 U21039 ( .A(n25958), .B(n25959), .C(n25960), .Y(n25957) );
  OAI21X1 U21040 ( .A(n25961), .B(n25962), .C(n25963), .Y(n25960) );
  OAI22X1 U21041 ( .A(n25964), .B(n25965), .C(n25966), .D(n25873), .Y(n25962)
         );
  OAI21X1 U21042 ( .A(n25967), .B(n25864), .C(n25968), .Y(n25961) );
  AOI22X1 U21043 ( .A(reg_A[71]), .B(n25969), .C(reg_B[93]), .D(n25970), .Y(
        n25968) );
  MUX2X1 U21044 ( .B(n25902), .A(n25971), .S(reg_B[93]), .Y(n25959) );
  NOR2X1 U21045 ( .A(n25972), .B(n25973), .Y(n25971) );
  INVX1 U21046 ( .A(n25974), .Y(n25958) );
  OAI22X1 U21047 ( .A(n25975), .B(n25976), .C(n25914), .D(n25977), .Y(n25956)
         );
  MUX2X1 U21048 ( .B(reg_A[93]), .A(reg_A[89]), .S(reg_B[93]), .Y(n25977) );
  INVX1 U21049 ( .A(n25978), .Y(n25975) );
  AOI22X1 U21050 ( .A(n25604), .B(n25979), .C(n25980), .D(n25981), .Y(n25954)
         );
  OAI21X1 U21051 ( .A(n25982), .B(n25914), .C(n25983), .Y(n25979) );
  AOI22X1 U21052 ( .A(n25984), .B(n25985), .C(reg_B[95]), .D(n25986), .Y(
        n25983) );
  INVX1 U21053 ( .A(n25987), .Y(n25985) );
  AOI22X1 U21054 ( .A(n25988), .B(reg_A[87]), .C(reg_A[83]), .D(n25989), .Y(
        n25987) );
  INVX1 U21055 ( .A(n25990), .Y(n25982) );
  INVX1 U21056 ( .A(n25991), .Y(n25949) );
  NOR2X1 U21057 ( .A(n25992), .B(n25993), .Y(n25828) );
  OAI21X1 U21058 ( .A(n25994), .B(n25995), .C(n25996), .Y(n25993) );
  OAI21X1 U21059 ( .A(n25997), .B(n25998), .C(n25999), .Y(n25996) );
  NAND2X1 U21060 ( .A(n26000), .B(n26001), .Y(n25998) );
  AOI22X1 U21061 ( .A(reg_A[88]), .B(n26002), .C(reg_A[91]), .D(n26003), .Y(
        n26001) );
  AOI22X1 U21062 ( .A(reg_A[90]), .B(n25751), .C(reg_A[95]), .D(n26004), .Y(
        n26000) );
  NAND2X1 U21063 ( .A(n26005), .B(n26006), .Y(n25997) );
  AOI22X1 U21064 ( .A(reg_A[94]), .B(n26007), .C(reg_A[92]), .D(n26008), .Y(
        n26006) );
  AOI22X1 U21065 ( .A(reg_A[93]), .B(n26009), .C(reg_A[89]), .D(n26010), .Y(
        n26005) );
  OAI21X1 U21066 ( .A(n26011), .B(n26012), .C(n26013), .Y(n25992) );
  AOI22X1 U21067 ( .A(n26014), .B(n26015), .C(reg_A[94]), .D(n26016), .Y(
        n26013) );
  OR2X1 U21068 ( .A(n26017), .B(n26018), .Y(result[94]) );
  NAND3X1 U21069 ( .A(n26019), .B(n26020), .C(n26021), .Y(n26018) );
  NOR2X1 U21070 ( .A(n26022), .B(n26023), .Y(n26021) );
  OAI21X1 U21071 ( .A(n26012), .B(n26024), .C(n26025), .Y(n26023) );
  AOI22X1 U21072 ( .A(reg_A[90]), .B(n26026), .C(n26027), .D(n26028), .Y(
        n26025) );
  INVX1 U21073 ( .A(n26011), .Y(n26027) );
  OAI21X1 U21074 ( .A(n26029), .B(n26030), .C(n26031), .Y(n26011) );
  AOI22X1 U21075 ( .A(n26032), .B(n26033), .C(n25025), .D(n26035), .Y(n26031)
         );
  OAI21X1 U21076 ( .A(reg_A[94]), .B(n25063), .C(n26037), .Y(n26033) );
  AOI22X1 U21077 ( .A(n26038), .B(n26039), .C(reg_B[0]), .D(n26040), .Y(n26037) );
  OAI21X1 U21078 ( .A(n26041), .B(n25929), .C(n26042), .Y(n26022) );
  AOI22X1 U21079 ( .A(reg_A[88]), .B(n26043), .C(reg_A[94]), .D(n26044), .Y(
        n26042) );
  AOI21X1 U21080 ( .A(n26045), .B(n26046), .C(n26047), .Y(n26020) );
  INVX1 U21081 ( .A(n26048), .Y(n26047) );
  AOI22X1 U21082 ( .A(n25986), .B(n26049), .C(n25981), .D(n26050), .Y(n26048)
         );
  NAND2X1 U21083 ( .A(n26051), .B(n26052), .Y(n25981) );
  MUX2X1 U21084 ( .B(n26053), .A(n26054), .S(reg_B[94]), .Y(n26052) );
  OAI21X1 U21085 ( .A(n25964), .B(n26039), .C(n26055), .Y(n26053) );
  AOI22X1 U21086 ( .A(reg_A[78]), .B(n26056), .C(reg_A[94]), .D(n26057), .Y(
        n26055) );
  AOI22X1 U21087 ( .A(n26058), .B(reg_A[70]), .C(n26059), .D(n26060), .Y(
        n26051) );
  AND2X1 U21088 ( .A(n26061), .B(n25838), .Y(n26058) );
  OAI21X1 U21089 ( .A(n26062), .B(n26063), .C(n26064), .Y(n25986) );
  MUX2X1 U21090 ( .B(n26065), .A(n26066), .S(reg_B[94]), .Y(n26064) );
  OAI22X1 U21091 ( .A(n26067), .B(n25883), .C(n26068), .D(n26069), .Y(n26065)
         );
  AOI22X1 U21092 ( .A(n25838), .B(reg_A[86]), .C(n26059), .D(reg_A[82]), .Y(
        n26062) );
  NAND3X1 U21093 ( .A(n26070), .B(n26071), .C(n26072), .Y(n26046) );
  NOR2X1 U21094 ( .A(n26073), .B(n26074), .Y(n26072) );
  OAI22X1 U21095 ( .A(n25598), .B(n25882), .C(n25599), .D(n25973), .Y(n26074)
         );
  OAI21X1 U21096 ( .A(n25600), .B(n25929), .C(n26075), .Y(n26073) );
  OAI21X1 U21097 ( .A(n26076), .B(n26077), .C(n25604), .Y(n26075) );
  NAND2X1 U21098 ( .A(n26078), .B(n26079), .Y(n26077) );
  AOI22X1 U21099 ( .A(reg_A[84]), .B(n25607), .C(reg_A[80]), .D(n25608), .Y(
        n26079) );
  AOI22X1 U21100 ( .A(reg_A[82]), .B(n25609), .C(reg_A[81]), .D(n25610), .Y(
        n26078) );
  NAND2X1 U21101 ( .A(n26080), .B(n26081), .Y(n26076) );
  AOI22X1 U21102 ( .A(reg_A[87]), .B(n25613), .C(reg_A[85]), .D(n25614), .Y(
        n26081) );
  AOI22X1 U21103 ( .A(reg_A[86]), .B(n25615), .C(reg_A[83]), .D(n25616), .Y(
        n26080) );
  AOI21X1 U21104 ( .A(reg_A[93]), .B(n25617), .C(n26082), .Y(n26071) );
  OAI21X1 U21105 ( .A(n25619), .B(n25883), .C(n26083), .Y(n26082) );
  OAI21X1 U21106 ( .A(n26084), .B(n26085), .C(n25044), .Y(n26083) );
  NAND2X1 U21107 ( .A(n26086), .B(n26087), .Y(n26085) );
  NOR2X1 U21108 ( .A(n26088), .B(n26089), .Y(n26087) );
  OAI21X1 U21109 ( .A(n25034), .B(n26039), .C(n26090), .Y(n26089) );
  AOI22X1 U21110 ( .A(reg_A[87]), .B(n25628), .C(reg_A[85]), .D(n25629), .Y(
        n26090) );
  OAI21X1 U21111 ( .A(n25498), .B(n25855), .C(n26091), .Y(n26088) );
  AOI22X1 U21112 ( .A(reg_A[64]), .B(n25631), .C(reg_A[66]), .D(n25324), .Y(
        n26091) );
  NOR2X1 U21113 ( .A(n26092), .B(n26093), .Y(n26086) );
  OAI21X1 U21114 ( .A(n25039), .B(n26094), .C(n26095), .Y(n26093) );
  AOI22X1 U21115 ( .A(reg_A[79]), .B(n25235), .C(reg_A[82]), .D(n25635), .Y(
        n26095) );
  OAI21X1 U21116 ( .A(n25035), .B(n25584), .C(n26096), .Y(n26092) );
  AOI22X1 U21117 ( .A(reg_A[83]), .B(n25222), .C(reg_A[84]), .D(n25637), .Y(
        n26096) );
  NAND2X1 U21118 ( .A(n26097), .B(n26098), .Y(n26084) );
  NOR2X1 U21119 ( .A(n26099), .B(n26100), .Y(n26098) );
  OAI21X1 U21120 ( .A(n25050), .B(n26101), .C(n26102), .Y(n26100) );
  AOI22X1 U21121 ( .A(reg_A[76]), .B(n25241), .C(reg_A[72]), .D(n25242), .Y(
        n26102) );
  OAI21X1 U21122 ( .A(n25038), .B(n26103), .C(n26104), .Y(n26099) );
  AOI22X1 U21123 ( .A(reg_A[77]), .B(n25246), .C(reg_A[78]), .D(n25247), .Y(
        n26104) );
  NOR2X1 U21124 ( .A(n26105), .B(n26106), .Y(n26097) );
  OAI21X1 U21125 ( .A(n25059), .B(n26107), .C(n26108), .Y(n26106) );
  AOI22X1 U21126 ( .A(reg_A[70]), .B(n25647), .C(reg_A[67]), .D(n25648), .Y(
        n26108) );
  OAI21X1 U21127 ( .A(n25054), .B(n25856), .C(n26109), .Y(n26105) );
  AOI22X1 U21128 ( .A(reg_A[74]), .B(n25339), .C(reg_A[73]), .D(n25257), .Y(
        n26109) );
  AOI22X1 U21129 ( .A(reg_A[90]), .B(n25650), .C(reg_A[88]), .D(n25651), .Y(
        n26070) );
  INVX1 U21130 ( .A(n26110), .Y(n26019) );
  OAI21X1 U21131 ( .A(n26111), .B(n26112), .C(n26113), .Y(n26110) );
  AOI22X1 U21132 ( .A(n26114), .B(n25903), .C(n26115), .D(n26116), .Y(n26113)
         );
  NAND3X1 U21133 ( .A(n26117), .B(n26118), .C(n26119), .Y(n26017) );
  NOR2X1 U21134 ( .A(n26120), .B(n26121), .Y(n26119) );
  OAI21X1 U21135 ( .A(n26122), .B(n25881), .C(n26123), .Y(n26121) );
  AOI22X1 U21136 ( .A(n26124), .B(n26014), .C(n26015), .D(n26125), .Y(n26123)
         );
  AOI21X1 U21137 ( .A(n26126), .B(n26059), .C(n26127), .Y(n26015) );
  INVX1 U21138 ( .A(n26128), .Y(n26127) );
  AOI22X1 U21139 ( .A(n25838), .B(n26129), .C(reg_B[94]), .D(n26130), .Y(
        n26128) );
  OAI21X1 U21140 ( .A(reg_A[86]), .B(n26131), .C(n26132), .Y(n26129) );
  AOI22X1 U21141 ( .A(reg_B[91]), .B(n26133), .C(n26134), .D(n25883), .Y(
        n26132) );
  INVX1 U21142 ( .A(n26135), .Y(n26124) );
  OAI21X1 U21143 ( .A(n25873), .B(n26136), .C(n26137), .Y(n26120) );
  AOI22X1 U21144 ( .A(reg_B[93]), .B(n26138), .C(n26139), .D(n26140), .Y(
        n26137) );
  INVX1 U21145 ( .A(n26141), .Y(n26140) );
  NOR2X1 U21146 ( .A(n26142), .B(n26143), .Y(n26118) );
  OAI22X1 U21147 ( .A(n26144), .B(n26145), .C(n26146), .D(n26147), .Y(n26143)
         );
  AOI22X1 U21148 ( .A(n26148), .B(n25990), .C(n26149), .D(n26150), .Y(n26146)
         );
  OAI21X1 U21149 ( .A(n26151), .B(n26152), .C(n26153), .Y(n26142) );
  NAND3X1 U21150 ( .A(n25988), .B(n25188), .C(n26154), .Y(n26153) );
  INVX1 U21151 ( .A(n26155), .Y(n26154) );
  MUX2X1 U21152 ( .B(n25978), .A(n26156), .S(reg_B[95]), .Y(n26152) );
  NAND2X1 U21153 ( .A(n26157), .B(n26158), .Y(n25978) );
  AOI22X1 U21154 ( .A(n26159), .B(reg_A[88]), .C(n26160), .D(reg_A[92]), .Y(
        n26158) );
  AOI22X1 U21155 ( .A(n25838), .B(reg_A[94]), .C(n26059), .D(reg_A[90]), .Y(
        n26157) );
  AOI21X1 U21156 ( .A(reg_A[91]), .B(n26161), .C(n26162), .Y(n26117) );
  OAI21X1 U21157 ( .A(n26163), .B(n25882), .C(n26164), .Y(n26162) );
  OAI21X1 U21158 ( .A(n26165), .B(n26166), .C(n26167), .Y(n26164) );
  OAI22X1 U21159 ( .A(n25881), .B(n26168), .C(n25973), .D(n26169), .Y(n26166)
         );
  OAI21X1 U21160 ( .A(n25914), .B(n25882), .C(n26170), .Y(n26165) );
  NAND3X1 U21161 ( .A(n26171), .B(n26172), .C(n26173), .Y(result[93]) );
  NOR2X1 U21162 ( .A(n26174), .B(n26175), .Y(n26173) );
  NAND3X1 U21163 ( .A(n26176), .B(n26177), .C(n26178), .Y(n26175) );
  AOI21X1 U21164 ( .A(n26179), .B(reg_A[93]), .C(n26180), .Y(n26178) );
  OAI22X1 U21165 ( .A(n26112), .B(n26111), .C(n26181), .D(n26182), .Y(n26180)
         );
  MUX2X1 U21166 ( .B(n26183), .A(n26184), .S(reg_B[95]), .Y(n26177) );
  AND2X1 U21167 ( .A(n26185), .B(n25170), .Y(n26184) );
  AND2X1 U21168 ( .A(n26156), .B(n26186), .Y(n26183) );
  OAI21X1 U21169 ( .A(n25929), .B(n25898), .C(n26187), .Y(n26156) );
  AOI22X1 U21170 ( .A(n26160), .B(reg_A[91]), .C(n25838), .D(reg_A[93]), .Y(
        n26187) );
  MUX2X1 U21171 ( .B(n25991), .A(n26188), .S(reg_B[94]), .Y(n26176) );
  AND2X1 U21172 ( .A(n25188), .B(n26189), .Y(n26188) );
  OAI22X1 U21173 ( .A(n26190), .B(n26191), .C(n25342), .D(n26192), .Y(n25991)
         );
  MUX2X1 U21174 ( .B(n26193), .A(n26194), .S(reg_B[93]), .Y(n26192) );
  MUX2X1 U21175 ( .B(n25929), .A(n26195), .S(reg_B[95]), .Y(n26194) );
  OAI21X1 U21176 ( .A(n26196), .B(n26197), .C(n25188), .Y(n26191) );
  OAI22X1 U21177 ( .A(n26198), .B(n26199), .C(n26193), .D(n26067), .Y(n26190)
         );
  MUX2X1 U21178 ( .B(n25881), .A(n25882), .S(reg_B[95]), .Y(n26193) );
  NAND3X1 U21179 ( .A(n26200), .B(n26201), .C(n26202), .Y(n26174) );
  AOI21X1 U21180 ( .A(n26203), .B(n26028), .C(n26204), .Y(n26202) );
  OAI22X1 U21181 ( .A(n26205), .B(n26068), .C(n26206), .D(n25973), .Y(n26204)
         );
  INVX1 U21182 ( .A(n26024), .Y(n26203) );
  OAI21X1 U21183 ( .A(n26207), .B(n26208), .C(n26209), .Y(n26024) );
  AOI22X1 U21184 ( .A(n25026), .B(n25934), .C(n25938), .D(n26030), .Y(n26209)
         );
  INVX1 U21185 ( .A(n26211), .Y(n25938) );
  MUX2X1 U21186 ( .B(n26212), .A(n26213), .S(reg_B[2]), .Y(n26211) );
  OAI21X1 U21187 ( .A(reg_A[93]), .B(n25063), .C(n26214), .Y(n26212) );
  AOI22X1 U21188 ( .A(n26038), .B(n26215), .C(reg_B[0]), .D(n26216), .Y(n26214) );
  OAI21X1 U21189 ( .A(n26217), .B(n26218), .C(n26045), .Y(n26201) );
  NAND3X1 U21190 ( .A(n26219), .B(n26220), .C(n26221), .Y(n26218) );
  AOI21X1 U21191 ( .A(reg_A[93]), .B(n25434), .C(n26222), .Y(n26221) );
  OAI22X1 U21192 ( .A(n25437), .B(n25973), .C(n25438), .D(n25929), .Y(n26222)
         );
  AOI22X1 U21193 ( .A(reg_A[87]), .B(n25440), .C(n26223), .D(n25610), .Y(
        n26220) );
  AOI22X1 U21194 ( .A(reg_A[92]), .B(n25441), .C(reg_A[90]), .D(n25442), .Y(
        n26219) );
  NAND3X1 U21195 ( .A(n26224), .B(n26225), .C(n26226), .Y(n26217) );
  NOR2X1 U21196 ( .A(n26227), .B(n26228), .Y(n26226) );
  OAI22X1 U21197 ( .A(n26229), .B(n26230), .C(n25449), .D(n26195), .Y(n26228)
         );
  OAI21X1 U21198 ( .A(n25451), .B(n26094), .C(n26231), .Y(n26227) );
  OAI21X1 U21199 ( .A(n26232), .B(n26233), .C(n25044), .Y(n26231) );
  NAND3X1 U21200 ( .A(n26234), .B(n26235), .C(n26236), .Y(n26233) );
  NOR2X1 U21201 ( .A(n26237), .B(n26238), .Y(n26236) );
  OAI21X1 U21202 ( .A(n25043), .B(n25881), .C(n26239), .Y(n26238) );
  AOI22X1 U21203 ( .A(reg_A[92]), .B(n25135), .C(reg_A[91]), .D(n25252), .Y(
        n26239) );
  NAND2X1 U21204 ( .A(n26240), .B(n26241), .Y(n26237) );
  AOI22X1 U21205 ( .A(reg_A[90]), .B(n25136), .C(reg_A[87]), .D(n25253), .Y(
        n26241) );
  AOI22X1 U21206 ( .A(reg_A[89]), .B(n25071), .C(reg_A[88]), .D(n25123), .Y(
        n26240) );
  NOR2X1 U21207 ( .A(n26242), .B(n26243), .Y(n26235) );
  OAI22X1 U21208 ( .A(n25034), .B(n26215), .C(n25129), .D(n26039), .Y(n26243)
         );
  OAI22X1 U21209 ( .A(n25036), .B(n25875), .C(n25223), .D(n26230), .Y(n26242)
         );
  NOR2X1 U21210 ( .A(n26244), .B(n26245), .Y(n26234) );
  OAI22X1 U21211 ( .A(n25064), .B(n26094), .C(n25473), .D(n25874), .Y(n26245)
         );
  OAI22X1 U21212 ( .A(n25039), .B(n25584), .C(n25035), .D(n25864), .Y(n26244)
         );
  NAND3X1 U21213 ( .A(n26246), .B(n26247), .C(n26248), .Y(n26232) );
  NOR2X1 U21214 ( .A(n26249), .B(n26250), .Y(n26248) );
  OAI21X1 U21215 ( .A(n25065), .B(n25865), .C(n26251), .Y(n26250) );
  AOI22X1 U21216 ( .A(reg_A[76]), .B(n25246), .C(reg_A[77]), .D(n25247), .Y(
        n26251) );
  NAND2X1 U21217 ( .A(n26252), .B(n26253), .Y(n26249) );
  AOI22X1 U21218 ( .A(reg_A[74]), .B(n25487), .C(reg_A[75]), .D(n25241), .Y(
        n26253) );
  AOI22X1 U21219 ( .A(reg_A[73]), .B(n25339), .C(reg_A[72]), .D(n25257), .Y(
        n26252) );
  NOR2X1 U21220 ( .A(n26254), .B(n26255), .Y(n26247) );
  OAI22X1 U21221 ( .A(n25491), .B(n26256), .C(n25492), .D(n26101), .Y(n26255)
         );
  OAI22X1 U21222 ( .A(n25057), .B(n25856), .C(n25322), .D(n26107), .Y(n26254)
         );
  NOR2X1 U21223 ( .A(n26257), .B(n26258), .Y(n26246) );
  OAI22X1 U21224 ( .A(n25316), .B(n25851), .C(n25318), .D(n25884), .Y(n26258)
         );
  OAI22X1 U21225 ( .A(n25498), .B(n25853), .C(n25499), .D(n25855), .Y(n26257)
         );
  AOI22X1 U21226 ( .A(reg_A[85]), .B(n25501), .C(reg_A[86]), .D(n25502), .Y(
        n26225) );
  AOI22X1 U21227 ( .A(reg_A[82]), .B(n25503), .C(reg_A[83]), .D(n25439), .Y(
        n26224) );
  AOI22X1 U21228 ( .A(n26259), .B(n26260), .C(n26261), .D(n26262), .Y(n26200)
         );
  NOR2X1 U21229 ( .A(n26263), .B(n26264), .Y(n26172) );
  OAI21X1 U21230 ( .A(n26265), .B(n26195), .C(n26266), .Y(n26264) );
  AOI22X1 U21231 ( .A(n26267), .B(n26268), .C(n26269), .D(reg_A[89]), .Y(
        n26266) );
  NAND2X1 U21232 ( .A(n26270), .B(n26271), .Y(n26268) );
  AOI22X1 U21233 ( .A(n25984), .B(n25990), .C(n26148), .D(n26066), .Y(n26271)
         );
  NAND2X1 U21234 ( .A(n26272), .B(n26273), .Y(n25990) );
  AOI22X1 U21235 ( .A(n25989), .B(reg_A[81]), .C(reg_A[85]), .D(n25988), .Y(
        n26273) );
  AOI22X1 U21236 ( .A(n26274), .B(reg_A[89]), .C(reg_A[93]), .D(n26275), .Y(
        n26272) );
  AOI22X1 U21237 ( .A(n26276), .B(n26150), .C(n26149), .D(n26277), .Y(n26270)
         );
  OAI21X1 U21238 ( .A(n25944), .B(n26278), .C(n26279), .Y(n26263) );
  AOI22X1 U21239 ( .A(n26280), .B(n26160), .C(n26281), .D(n26115), .Y(n26279)
         );
  OAI21X1 U21240 ( .A(n26282), .B(n26112), .C(n26283), .Y(n26115) );
  AOI22X1 U21241 ( .A(n25930), .B(n25950), .C(n26160), .D(n25970), .Y(n26283)
         );
  OR2X1 U21242 ( .A(n26284), .B(n26285), .Y(n25930) );
  OAI22X1 U21243 ( .A(n25964), .B(n26215), .C(n25966), .D(n25881), .Y(n26285)
         );
  OAI21X1 U21244 ( .A(n25967), .B(n26286), .C(n26287), .Y(n26284) );
  AOI22X1 U21245 ( .A(reg_A[69]), .B(n25969), .C(reg_B[93]), .D(n26288), .Y(
        n26287) );
  INVX1 U21246 ( .A(n26289), .Y(n26282) );
  NOR2X1 U21247 ( .A(n25907), .B(n25031), .Y(n26280) );
  MUX2X1 U21248 ( .B(reg_A[91]), .A(reg_A[90]), .S(reg_B[95]), .Y(n25907) );
  NAND2X1 U21249 ( .A(n26290), .B(n26291), .Y(n25944) );
  AOI22X1 U21250 ( .A(n26292), .B(n25929), .C(n26293), .D(n25881), .Y(n26291)
         );
  AOI22X1 U21251 ( .A(n26294), .B(n26195), .C(n26295), .D(n25882), .Y(n26290)
         );
  NOR2X1 U21252 ( .A(n26296), .B(n26297), .Y(n26171) );
  OAI22X1 U21253 ( .A(n25886), .B(n26135), .C(n26298), .D(n26299), .Y(n26297)
         );
  OAI21X1 U21254 ( .A(n26300), .B(n26112), .C(n26301), .Y(n26135) );
  AOI22X1 U21255 ( .A(n25933), .B(n25950), .C(n26160), .D(n25906), .Y(n26301)
         );
  NAND2X1 U21256 ( .A(n26302), .B(n26303), .Y(n25933) );
  MUX2X1 U21257 ( .B(n26304), .A(n26305), .S(reg_B[93]), .Y(n26303) );
  NOR2X1 U21258 ( .A(n26306), .B(n25895), .Y(n26304) );
  AOI22X1 U21259 ( .A(n26057), .B(n25881), .C(n26307), .D(n26215), .Y(n26302)
         );
  OAI21X1 U21260 ( .A(n25883), .B(n26136), .C(n26308), .Y(n26296) );
  AOI22X1 U21261 ( .A(n26309), .B(n25150), .C(n26310), .D(reg_A[95]), .Y(
        n26308) );
  INVX1 U21262 ( .A(n25995), .Y(n26309) );
  NAND2X1 U21263 ( .A(n26311), .B(n26312), .Y(n25995) );
  AOI22X1 U21264 ( .A(n26313), .B(n25882), .C(n26314), .D(n25881), .Y(n26312)
         );
  AOI22X1 U21265 ( .A(reg_B[1]), .B(n26315), .C(reg_B[2]), .D(n26316), .Y(
        n26311) );
  INVX1 U21266 ( .A(n26317), .Y(n26315) );
  NAND3X1 U21267 ( .A(n26318), .B(n26319), .C(n26320), .Y(result[92]) );
  NOR2X1 U21268 ( .A(n26321), .B(n26322), .Y(n26320) );
  NAND3X1 U21269 ( .A(n26323), .B(n26324), .C(n26325), .Y(n26322) );
  NOR2X1 U21270 ( .A(n26326), .B(n26327), .Y(n26325) );
  OAI22X1 U21271 ( .A(n26328), .B(n26215), .C(n26181), .D(n26329), .Y(n26327)
         );
  MUX2X1 U21272 ( .B(n26330), .A(n26331), .S(reg_B[95]), .Y(n26326) );
  INVX1 U21273 ( .A(n26332), .Y(n26331) );
  NAND2X1 U21274 ( .A(n25170), .B(n26185), .Y(n26330) );
  OAI21X1 U21275 ( .A(n26333), .B(n25403), .C(n26334), .Y(n26185) );
  OAI21X1 U21276 ( .A(n26335), .B(n26336), .C(n25589), .Y(n26334) );
  OAI22X1 U21277 ( .A(n25882), .B(n26337), .C(n26068), .D(n26338), .Y(n26336)
         );
  NOR2X1 U21278 ( .A(n26195), .B(n25898), .Y(n26335) );
  AOI21X1 U21279 ( .A(n26159), .B(n26339), .C(n26340), .Y(n26333) );
  INVX1 U21280 ( .A(n26341), .Y(n26340) );
  AOI22X1 U21281 ( .A(n26060), .B(n26160), .C(n25950), .D(n26054), .Y(n26341)
         );
  OR2X1 U21282 ( .A(n26342), .B(n26343), .Y(n26054) );
  OAI22X1 U21283 ( .A(n25964), .B(n26230), .C(n25966), .D(n25882), .Y(n26343)
         );
  OAI21X1 U21284 ( .A(n25967), .B(n25863), .C(n26344), .Y(n26342) );
  AOI22X1 U21285 ( .A(reg_A[68]), .B(n25969), .C(reg_B[93]), .D(n26345), .Y(
        n26344) );
  NOR2X1 U21286 ( .A(n25895), .B(n26199), .Y(n25969) );
  AOI22X1 U21287 ( .A(reg_A[83]), .B(n26346), .C(reg_A[86]), .D(n26347), .Y(
        n26324) );
  AOI22X1 U21288 ( .A(reg_A[88]), .B(n26348), .C(n26349), .D(reg_A[77]), .Y(
        n26323) );
  NAND3X1 U21289 ( .A(n26350), .B(n26351), .C(n26352), .Y(n26321) );
  AOI21X1 U21290 ( .A(reg_A[87]), .B(n26353), .C(n26354), .Y(n26352) );
  OAI22X1 U21291 ( .A(n26355), .B(n26230), .C(n26012), .D(n26356), .Y(n26354)
         );
  AOI22X1 U21292 ( .A(reg_A[81]), .B(n26357), .C(reg_A[91]), .D(n26358), .Y(
        n26351) );
  AOI22X1 U21293 ( .A(reg_A[82]), .B(n26359), .C(n26259), .D(n26028), .Y(
        n26350) );
  INVX1 U21294 ( .A(n26360), .Y(n26259) );
  OAI21X1 U21295 ( .A(n26361), .B(n26208), .C(n26362), .Y(n26360) );
  AOI22X1 U21296 ( .A(n25026), .B(n26035), .C(n26363), .D(n26030), .Y(n26362)
         );
  INVX1 U21297 ( .A(n26029), .Y(n26363) );
  MUX2X1 U21298 ( .B(n26364), .A(n26365), .S(reg_B[2]), .Y(n26029) );
  OAI21X1 U21299 ( .A(reg_A[92]), .B(n25063), .C(n26366), .Y(n26364) );
  AOI22X1 U21300 ( .A(n26038), .B(n26230), .C(reg_B[0]), .D(n26367), .Y(n26366) );
  NOR2X1 U21301 ( .A(n26368), .B(n26369), .Y(n26319) );
  OAI21X1 U21302 ( .A(n26370), .B(n25584), .C(n26371), .Y(n26369) );
  INVX1 U21303 ( .A(n26372), .Y(n26371) );
  OAI21X1 U21304 ( .A(n25929), .B(n26373), .C(n26374), .Y(n26372) );
  OAI21X1 U21305 ( .A(n26375), .B(n26376), .C(n25188), .Y(n26374) );
  OAI21X1 U21306 ( .A(n26377), .B(n25882), .C(n26378), .Y(n26376) );
  AOI22X1 U21307 ( .A(n26379), .B(n25988), .C(n26380), .D(n26274), .Y(n26378)
         );
  OAI21X1 U21308 ( .A(n25973), .B(n26381), .C(n26382), .Y(n26375) );
  AOI21X1 U21309 ( .A(n26383), .B(n26149), .C(n26384), .Y(n26382) );
  INVX1 U21310 ( .A(n26385), .Y(n26384) );
  NOR2X1 U21311 ( .A(n26067), .B(n25929), .Y(n26383) );
  NAND3X1 U21312 ( .A(n26386), .B(n26387), .C(n26388), .Y(n26368) );
  AOI21X1 U21313 ( .A(reg_A[90]), .B(n26389), .C(n26390), .Y(n26388) );
  INVX1 U21314 ( .A(n26391), .Y(n26390) );
  OAI21X1 U21315 ( .A(n26392), .B(n25914), .C(n26393), .Y(n26389) );
  INVX1 U21316 ( .A(n26167), .Y(n26392) );
  NAND2X1 U21317 ( .A(n26394), .B(n26395), .Y(n26167) );
  INVX1 U21318 ( .A(n26396), .Y(n26395) );
  OAI21X1 U21319 ( .A(n26397), .B(n26398), .C(reg_A[92]), .Y(n26387) );
  INVX1 U21320 ( .A(n26399), .Y(n26386) );
  AOI21X1 U21321 ( .A(n26400), .B(n26401), .C(n26147), .Y(n26399) );
  AOI22X1 U21322 ( .A(n26402), .B(n26149), .C(n26277), .D(n26276), .Y(n26401)
         );
  AOI22X1 U21323 ( .A(n26150), .B(n26148), .C(n26066), .D(n25984), .Y(n26400)
         );
  OR2X1 U21324 ( .A(n26403), .B(n26404), .Y(n26066) );
  OAI22X1 U21325 ( .A(n26195), .B(n26069), .C(n26067), .D(n25882), .Y(n26404)
         );
  OAI21X1 U21326 ( .A(n26199), .B(n26230), .C(n26385), .Y(n26403) );
  NOR2X1 U21327 ( .A(n26405), .B(n26406), .Y(n26318) );
  OAI21X1 U21328 ( .A(n25886), .B(n26299), .C(n26407), .Y(n26406) );
  AOI22X1 U21329 ( .A(n26310), .B(reg_A[94]), .C(n26408), .D(reg_A[93]), .Y(
        n26407) );
  OAI21X1 U21330 ( .A(n26409), .B(n26112), .C(n26410), .Y(n26299) );
  AOI22X1 U21331 ( .A(n26130), .B(n25950), .C(n26160), .D(n26126), .Y(n26410)
         );
  NAND2X1 U21332 ( .A(n26411), .B(n26412), .Y(n26130) );
  MUX2X1 U21333 ( .B(n26413), .A(n26414), .S(reg_B[93]), .Y(n26412) );
  NOR2X1 U21334 ( .A(n26415), .B(n25895), .Y(n26413) );
  AOI22X1 U21335 ( .A(n26057), .B(n25882), .C(n26307), .D(n26230), .Y(n26411)
         );
  OR2X1 U21336 ( .A(n26416), .B(n26417), .Y(n26405) );
  OAI22X1 U21337 ( .A(n25873), .B(n26418), .C(n26419), .D(n26420), .Y(n26417)
         );
  OAI21X1 U21338 ( .A(n26421), .B(n26422), .C(n26423), .Y(n26416) );
  OAI21X1 U21339 ( .A(n26424), .B(n26425), .C(n25840), .Y(n26423) );
  NAND3X1 U21340 ( .A(n26426), .B(n26427), .C(n26428), .Y(n26425) );
  NOR2X1 U21341 ( .A(n26429), .B(n26430), .Y(n26428) );
  OAI22X1 U21342 ( .A(n25039), .B(n25864), .C(n25475), .D(n25865), .Y(n26430)
         );
  OAI22X1 U21343 ( .A(n26431), .B(n26195), .C(n25784), .D(n25973), .Y(n26429)
         );
  AOI22X1 U21344 ( .A(reg_A[68]), .B(n25647), .C(reg_A[65]), .D(n25648), .Y(
        n26427) );
  AOI22X1 U21345 ( .A(reg_A[66]), .B(n26432), .C(reg_A[64]), .D(n25324), .Y(
        n26426) );
  NAND3X1 U21346 ( .A(n26433), .B(n26434), .C(n26435), .Y(n26424) );
  NOR2X1 U21347 ( .A(n26436), .B(n26437), .Y(n26435) );
  OAI22X1 U21348 ( .A(n25492), .B(n26256), .C(n25331), .D(n26438), .Y(n26437)
         );
  OAI21X1 U21349 ( .A(n25038), .B(n26439), .C(n26440), .Y(n26436) );
  AOI22X1 U21350 ( .A(reg_A[75]), .B(n25246), .C(reg_A[76]), .D(n25247), .Y(
        n26440) );
  AOI22X1 U21351 ( .A(reg_A[69]), .B(n25338), .C(reg_A[72]), .D(n25339), .Y(
        n26434) );
  AOI22X1 U21352 ( .A(reg_A[71]), .B(n25257), .C(reg_A[67]), .D(n25857), .Y(
        n26433) );
  NAND2X1 U21353 ( .A(n26441), .B(n26442), .Y(result[91]) );
  NOR2X1 U21354 ( .A(n26443), .B(n26444), .Y(n26442) );
  NAND3X1 U21355 ( .A(n26445), .B(n26446), .C(n26447), .Y(n26444) );
  AOI21X1 U21356 ( .A(reg_A[80]), .B(n26357), .C(n26448), .Y(n26447) );
  OAI22X1 U21357 ( .A(n26298), .B(n26449), .C(n25882), .D(n26136), .Y(n26448)
         );
  AOI22X1 U21358 ( .A(reg_A[91]), .B(n26450), .C(n26451), .D(reg_A[94]), .Y(
        n26446) );
  AOI22X1 U21359 ( .A(n26261), .B(n25150), .C(n26310), .D(reg_A[93]), .Y(
        n26445) );
  AOI21X1 U21360 ( .A(n26452), .B(n25940), .C(n26453), .Y(n26261) );
  INVX1 U21361 ( .A(n26454), .Y(n26453) );
  AOI22X1 U21362 ( .A(n26455), .B(n25584), .C(n26456), .D(n26457), .Y(n26454)
         );
  NAND2X1 U21363 ( .A(n26458), .B(n26459), .Y(n25940) );
  AOI22X1 U21364 ( .A(n26460), .B(n25875), .C(n26461), .D(n25973), .Y(n26459)
         );
  AOI22X1 U21365 ( .A(n26462), .B(n26068), .C(n26463), .D(n25874), .Y(n26458)
         );
  NAND3X1 U21366 ( .A(n26464), .B(n26465), .C(n26466), .Y(n26443) );
  NOR2X1 U21367 ( .A(n26467), .B(n26468), .Y(n26466) );
  OAI21X1 U21368 ( .A(n25032), .B(n26469), .C(n26470), .Y(n26468) );
  OAI21X1 U21369 ( .A(n26471), .B(n26472), .C(reg_A[88]), .Y(n26470) );
  INVX1 U21370 ( .A(n26473), .Y(n26471) );
  MUX2X1 U21371 ( .B(n26189), .A(n26474), .S(reg_B[94]), .Y(n26469) );
  AOI21X1 U21372 ( .A(n25584), .B(n25989), .C(n26475), .Y(n26189) );
  OAI22X1 U21373 ( .A(n25904), .B(reg_B[93]), .C(n26069), .D(n25891), .Y(
        n26475) );
  MUX2X1 U21374 ( .B(n26476), .A(n26477), .S(reg_B[95]), .Y(n25904) );
  MUX2X1 U21375 ( .B(reg_A[91]), .A(reg_A[83]), .S(reg_B[92]), .Y(n26476) );
  OAI21X1 U21376 ( .A(n26478), .B(n26479), .C(n26391), .Y(n26467) );
  AOI22X1 U21377 ( .A(n25382), .B(n25974), .C(n26480), .D(n26134), .Y(n26478)
         );
  AOI22X1 U21378 ( .A(reg_A[90]), .B(n26481), .C(n26482), .D(reg_A[95]), .Y(
        n26465) );
  OAI21X1 U21379 ( .A(n26168), .B(n26394), .C(n26483), .Y(n26481) );
  AOI21X1 U21380 ( .A(reg_A[89]), .B(n26484), .C(n26485), .Y(n26464) );
  AOI21X1 U21381 ( .A(n26486), .B(n26487), .C(n26147), .Y(n26485) );
  AOI22X1 U21382 ( .A(n25984), .B(n26150), .C(n26148), .D(n26277), .Y(n26487)
         );
  OAI21X1 U21383 ( .A(n26067), .B(n25973), .C(n26488), .Y(n26150) );
  AOI22X1 U21384 ( .A(reg_A[83]), .B(n25988), .C(n26274), .D(reg_A[87]), .Y(
        n26488) );
  AOI22X1 U21385 ( .A(n26276), .B(n26402), .C(n26149), .D(n26489), .Y(n26486)
         );
  INVX1 U21386 ( .A(n26490), .Y(n26484) );
  NOR2X1 U21387 ( .A(n26491), .B(n26492), .Y(n26441) );
  NAND3X1 U21388 ( .A(n26493), .B(n26494), .C(n26495), .Y(n26492) );
  NOR2X1 U21389 ( .A(n26496), .B(n26497), .Y(n26495) );
  OAI22X1 U21390 ( .A(n26328), .B(n26230), .C(n26169), .D(n26111), .Y(n26497)
         );
  INVX1 U21391 ( .A(n26498), .Y(n26496) );
  MUX2X1 U21392 ( .B(n26332), .A(n26499), .S(reg_B[95]), .Y(n26498) );
  OAI21X1 U21393 ( .A(n26500), .B(n26501), .C(n26502), .Y(n26332) );
  AOI22X1 U21394 ( .A(n25170), .B(n26503), .C(n26504), .D(n26505), .Y(n26502)
         );
  INVX1 U21395 ( .A(n26506), .Y(n26503) );
  AOI21X1 U21396 ( .A(n26505), .B(n25589), .C(n26507), .Y(n26506) );
  AOI21X1 U21397 ( .A(n26508), .B(n26509), .C(n25403), .Y(n26507) );
  AOI22X1 U21398 ( .A(n26510), .B(n26159), .C(n26289), .D(n26059), .Y(n26509)
         );
  AOI22X1 U21399 ( .A(n26288), .B(n26160), .C(n25970), .D(n25838), .Y(n26508)
         );
  NAND2X1 U21400 ( .A(n26511), .B(n26512), .Y(n25970) );
  AOI22X1 U21401 ( .A(reg_A[67]), .B(n26061), .C(reg_A[75]), .D(n26513), .Y(
        n26512) );
  AOI22X1 U21402 ( .A(reg_A[91]), .B(n26134), .C(reg_A[83]), .D(n25892), .Y(
        n26511) );
  OAI22X1 U21403 ( .A(n25973), .B(n26337), .C(n25929), .D(n26338), .Y(n26505)
         );
  OAI21X1 U21404 ( .A(n26514), .B(n26112), .C(n25932), .Y(n26501) );
  OAI21X1 U21405 ( .A(n26300), .B(n25898), .C(n26515), .Y(n26500) );
  AOI22X1 U21406 ( .A(n25838), .B(n25906), .C(n26160), .D(n26305), .Y(n26515)
         );
  OAI21X1 U21407 ( .A(reg_A[83]), .B(n26131), .C(n26516), .Y(n25906) );
  AOI22X1 U21408 ( .A(reg_B[91]), .B(n26517), .C(n26134), .D(n25973), .Y(
        n26516) );
  INVX1 U21409 ( .A(n26518), .Y(n26517) );
  AOI22X1 U21410 ( .A(reg_A[82]), .B(n26346), .C(reg_A[85]), .D(n26347), .Y(
        n26494) );
  AOI22X1 U21411 ( .A(n26519), .B(reg_A[79]), .C(n26349), .D(reg_A[76]), .Y(
        n26493) );
  NAND3X1 U21412 ( .A(n26520), .B(n26521), .C(n26522), .Y(n26491) );
  NOR2X1 U21413 ( .A(n26523), .B(n26524), .Y(n26522) );
  OAI22X1 U21414 ( .A(n26525), .B(n26356), .C(n26526), .D(n26094), .Y(n26524)
         );
  NAND2X1 U21415 ( .A(n26527), .B(n26528), .Y(n26356) );
  AOI22X1 U21416 ( .A(n25025), .B(n26529), .C(n25026), .D(n26213), .Y(n26528)
         );
  AOI22X1 U21417 ( .A(n26032), .B(n25934), .C(n26530), .D(n26531), .Y(n26527)
         );
  OAI21X1 U21418 ( .A(reg_A[91]), .B(n25063), .C(n26532), .Y(n25934) );
  AOI22X1 U21419 ( .A(n26038), .B(n25875), .C(reg_B[0]), .D(n26533), .Y(n26532) );
  OAI21X1 U21420 ( .A(n26534), .B(n25965), .C(n26535), .Y(n26523) );
  OAI21X1 U21421 ( .A(n26536), .B(n26537), .C(n25840), .Y(n26535) );
  NAND3X1 U21422 ( .A(n26538), .B(n26539), .C(n26540), .Y(n26537) );
  AOI21X1 U21423 ( .A(reg_A[78]), .B(n25325), .C(n26541), .Y(n26540) );
  OAI22X1 U21424 ( .A(n25035), .B(n26286), .C(n25042), .D(n26068), .Y(n26541)
         );
  AOI22X1 U21425 ( .A(reg_A[66]), .B(n25857), .C(reg_A[67]), .D(n25647), .Y(
        n26539) );
  AOI22X1 U21426 ( .A(reg_A[64]), .B(n25648), .C(reg_A[65]), .D(n26432), .Y(
        n26538) );
  NAND3X1 U21427 ( .A(n26542), .B(n26543), .C(n26544), .Y(n26536) );
  NOR2X1 U21428 ( .A(n26545), .B(n26546), .Y(n26544) );
  OAI22X1 U21429 ( .A(n25051), .B(n26439), .C(n25038), .D(n26547), .Y(n26546)
         );
  OAI22X1 U21430 ( .A(n25334), .B(n26103), .C(n25336), .D(n26438), .Y(n26545)
         );
  AOI22X1 U21431 ( .A(reg_A[69]), .B(n25242), .C(reg_A[68]), .D(n25338), .Y(
        n26543) );
  AOI22X1 U21432 ( .A(reg_A[71]), .B(n25339), .C(reg_A[70]), .D(n25257), .Y(
        n26542) );
  AOI22X1 U21433 ( .A(n26548), .B(n26260), .C(n26549), .D(n26262), .Y(n26521)
         );
  INVX1 U21434 ( .A(n26550), .Y(n26549) );
  AOI22X1 U21435 ( .A(reg_A[83]), .B(n26551), .C(reg_A[86]), .D(n26353), .Y(
        n26520) );
  NAND2X1 U21436 ( .A(n26552), .B(n26553), .Y(result[90]) );
  NOR2X1 U21437 ( .A(n26554), .B(n26555), .Y(n26553) );
  NAND3X1 U21438 ( .A(n26556), .B(n26557), .C(n26558), .Y(n26555) );
  NOR2X1 U21439 ( .A(n26559), .B(n26560), .Y(n26558) );
  OAI22X1 U21440 ( .A(n26141), .B(n26420), .C(reg_B[93]), .D(n26561), .Y(
        n26560) );
  INVX1 U21441 ( .A(n26138), .Y(n26561) );
  OAI21X1 U21442 ( .A(n26562), .B(n25342), .C(n26563), .Y(n26138) );
  NAND3X1 U21443 ( .A(n26564), .B(n25188), .C(n26565), .Y(n26563) );
  AOI22X1 U21444 ( .A(n25984), .B(n26477), .C(n26148), .D(n26566), .Y(n26565)
         );
  MUX2X1 U21445 ( .B(reg_A[82]), .A(reg_A[90]), .S(n26063), .Y(n26477) );
  MUX2X1 U21446 ( .B(n26567), .A(n26568), .S(reg_B[92]), .Y(n26564) );
  NOR2X1 U21447 ( .A(reg_A[80]), .B(n25950), .Y(n26568) );
  OAI22X1 U21448 ( .A(reg_A[87]), .B(n26169), .C(reg_A[88]), .D(n25914), .Y(
        n26567) );
  AOI22X1 U21449 ( .A(n26148), .B(reg_A[89]), .C(reg_A[90]), .D(n25984), .Y(
        n26562) );
  OAI21X1 U21450 ( .A(n26569), .B(n26068), .C(n26570), .Y(n26559) );
  AOI22X1 U21451 ( .A(reg_A[88]), .B(n26571), .C(reg_A[80]), .D(n26572), .Y(
        n26570) );
  INVX1 U21452 ( .A(n26573), .Y(n26571) );
  AOI22X1 U21453 ( .A(n26451), .B(reg_A[93]), .C(n26310), .D(reg_A[92]), .Y(
        n26557) );
  AOI22X1 U21454 ( .A(n26408), .B(reg_A[91]), .C(n26574), .D(n26014), .Y(
        n26556) );
  INVX1 U21455 ( .A(n26575), .Y(n26574) );
  NAND3X1 U21456 ( .A(n26576), .B(n26577), .C(n26578), .Y(n26554) );
  NOR2X1 U21457 ( .A(n26579), .B(n26580), .Y(n26578) );
  OAI22X1 U21458 ( .A(n25873), .B(n26581), .C(n26582), .D(n26583), .Y(n26580)
         );
  OAI21X1 U21459 ( .A(n26144), .B(n26584), .C(n26585), .Y(n26579) );
  AOI22X1 U21460 ( .A(n26586), .B(n26148), .C(n25188), .D(n26587), .Y(n26585)
         );
  OAI21X1 U21461 ( .A(n26069), .B(n26155), .C(n26385), .Y(n26587) );
  NAND2X1 U21462 ( .A(n25989), .B(reg_A[80]), .Y(n26385) );
  NAND2X1 U21463 ( .A(n26588), .B(n26589), .Y(n26155) );
  AOI22X1 U21464 ( .A(n26276), .B(n26230), .C(n26149), .D(n25875), .Y(n26589)
         );
  AOI22X1 U21465 ( .A(n26148), .B(n26215), .C(n25984), .D(n26039), .Y(n26588)
         );
  AND2X1 U21466 ( .A(n26590), .B(n25170), .Y(n26586) );
  NAND2X1 U21467 ( .A(n26591), .B(n26592), .Y(n26144) );
  AOI22X1 U21468 ( .A(n26593), .B(n25874), .C(n26594), .D(n25584), .Y(n26592)
         );
  AOI22X1 U21469 ( .A(n26595), .B(n26596), .C(n26597), .D(n26598), .Y(n26591)
         );
  OAI21X1 U21470 ( .A(reg_A[90]), .B(n26599), .C(n26600), .Y(n26595) );
  AOI22X1 U21471 ( .A(n26601), .B(n26195), .C(n26602), .D(n25965), .Y(n26600)
         );
  AOI22X1 U21472 ( .A(n26482), .B(reg_A[94]), .C(n26603), .D(n26114), .Y(
        n26577) );
  AOI22X1 U21473 ( .A(n26267), .B(n26604), .C(n26499), .D(n25976), .Y(n26576)
         );
  OAI21X1 U21474 ( .A(n26605), .B(n26151), .C(n26606), .Y(n26499) );
  INVX1 U21475 ( .A(n26607), .Y(n26606) );
  AOI21X1 U21476 ( .A(n26608), .B(n26609), .C(n26610), .Y(n26607) );
  AOI22X1 U21477 ( .A(n26611), .B(n26159), .C(n26339), .D(n26059), .Y(n26609)
         );
  AOI22X1 U21478 ( .A(n26345), .B(n26160), .C(n26060), .D(n25838), .Y(n26608)
         );
  NAND2X1 U21479 ( .A(n26612), .B(n26613), .Y(n26060) );
  AOI22X1 U21480 ( .A(reg_A[66]), .B(n26061), .C(reg_A[74]), .D(n26513), .Y(
        n26613) );
  AOI22X1 U21481 ( .A(reg_A[90]), .B(n26134), .C(reg_A[82]), .D(n25892), .Y(
        n26612) );
  AOI22X1 U21482 ( .A(n26160), .B(reg_A[88]), .C(n25838), .D(reg_A[90]), .Y(
        n26605) );
  OAI21X1 U21483 ( .A(n26614), .B(n26169), .C(n26615), .Y(n26604) );
  AOI22X1 U21484 ( .A(n25984), .B(n26277), .C(n26276), .D(n26489), .Y(n26615)
         );
  OAI21X1 U21485 ( .A(n26067), .B(n26068), .C(n26616), .Y(n26277) );
  AOI22X1 U21486 ( .A(reg_A[82]), .B(n25988), .C(n26274), .D(reg_A[86]), .Y(
        n26616) );
  NOR2X1 U21487 ( .A(n26617), .B(n26618), .Y(n26552) );
  NAND3X1 U21488 ( .A(n26619), .B(n26620), .C(n26621), .Y(n26618) );
  NOR2X1 U21489 ( .A(n26622), .B(n26623), .Y(n26621) );
  OAI22X1 U21490 ( .A(n26328), .B(n25875), .C(n25838), .D(n26111), .Y(n26623)
         );
  OAI22X1 U21491 ( .A(n26181), .B(n26624), .C(n26103), .D(n26625), .Y(n26622)
         );
  AOI22X1 U21492 ( .A(reg_A[84]), .B(n26347), .C(reg_A[89]), .D(n26626), .Y(
        n26620) );
  AOI22X1 U21493 ( .A(n26627), .B(reg_A[79]), .C(n26519), .D(reg_A[78]), .Y(
        n26619) );
  NAND3X1 U21494 ( .A(n26628), .B(n26629), .C(n26630), .Y(n26617) );
  NOR2X1 U21495 ( .A(n26631), .B(n26632), .Y(n26630) );
  OAI22X1 U21496 ( .A(n26633), .B(n26094), .C(n26634), .D(n25965), .Y(n26632)
         );
  OAI22X1 U21497 ( .A(n26635), .B(n26215), .C(n26355), .D(n25874), .Y(n26631)
         );
  INVX1 U21498 ( .A(n26353), .Y(n26635) );
  AOI21X1 U21499 ( .A(reg_A[86]), .B(n26636), .C(n26637), .Y(n26629) );
  OAI21X1 U21500 ( .A(n25886), .B(n26449), .C(n26638), .Y(n26637) );
  OAI21X1 U21501 ( .A(n26639), .B(n26640), .C(n25840), .Y(n26638) );
  NAND3X1 U21502 ( .A(n26641), .B(n26642), .C(n26643), .Y(n26640) );
  AOI21X1 U21503 ( .A(reg_A[77]), .B(n25325), .C(n26644), .Y(n26643) );
  OAI22X1 U21504 ( .A(n25035), .B(n25863), .C(n25042), .D(n25929), .Y(n26644)
         );
  AOI22X1 U21505 ( .A(reg_A[69]), .B(n25257), .C(reg_A[65]), .D(n25857), .Y(
        n26642) );
  AOI22X1 U21506 ( .A(reg_A[66]), .B(n25647), .C(reg_A[64]), .D(n26432), .Y(
        n26641) );
  NAND3X1 U21507 ( .A(n26645), .B(n26646), .C(n26647), .Y(n26639) );
  AOI21X1 U21508 ( .A(reg_A[70]), .B(n25339), .C(n26648), .Y(n26647) );
  OAI22X1 U21509 ( .A(n25491), .B(n25851), .C(n25492), .D(n26107), .Y(n26648)
         );
  AOI22X1 U21510 ( .A(reg_A[73]), .B(n25246), .C(reg_A[74]), .D(n25247), .Y(
        n26646) );
  AOI22X1 U21511 ( .A(reg_A[71]), .B(n25487), .C(reg_A[72]), .D(n25241), .Y(
        n26645) );
  NAND2X1 U21512 ( .A(n26649), .B(n26650), .Y(n26449) );
  AOI22X1 U21513 ( .A(n25838), .B(n26126), .C(n26160), .D(n26414), .Y(n26650)
         );
  NAND2X1 U21514 ( .A(n26651), .B(n26652), .Y(n26126) );
  AOI22X1 U21515 ( .A(n26061), .B(n25884), .C(n26513), .D(n26438), .Y(n26652)
         );
  AOI22X1 U21516 ( .A(n26134), .B(n26068), .C(n25892), .D(n25874), .Y(n26651)
         );
  AOI22X1 U21517 ( .A(n26059), .B(n26653), .C(n26159), .D(n26654), .Y(n26649)
         );
  AOI22X1 U21518 ( .A(n26548), .B(n26028), .C(n26655), .D(n26260), .Y(n26628)
         );
  AND2X1 U21519 ( .A(n26656), .B(n26657), .Y(n26548) );
  AOI22X1 U21520 ( .A(n25025), .B(n26658), .C(n25026), .D(n26365), .Y(n26657)
         );
  AOI22X1 U21521 ( .A(n26032), .B(n26035), .C(n26530), .D(n26659), .Y(n26656)
         );
  NAND2X1 U21522 ( .A(n26660), .B(n26661), .Y(n26035) );
  AOI22X1 U21523 ( .A(n26662), .B(n25884), .C(n26663), .D(n26438), .Y(n26661)
         );
  AOI22X1 U21524 ( .A(n26038), .B(n25874), .C(n26664), .D(n26068), .Y(n26660)
         );
  NAND3X1 U21525 ( .A(n26665), .B(n26666), .C(n26667), .Y(result[8]) );
  NOR2X1 U21526 ( .A(n26668), .B(n26669), .Y(n26667) );
  NAND3X1 U21527 ( .A(n26670), .B(n26671), .C(n26672), .Y(n26669) );
  AOI21X1 U21528 ( .A(reg_A[1]), .B(n26673), .C(n26674), .Y(n26672) );
  OAI22X1 U21529 ( .A(n26675), .B(n25255), .C(n26676), .D(n26677), .Y(n26674)
         );
  AOI22X1 U21530 ( .A(reg_A[2]), .B(n26678), .C(reg_A[3]), .D(n26679), .Y(
        n26671) );
  AOI22X1 U21531 ( .A(reg_A[4]), .B(n26680), .C(reg_A[5]), .D(n26681), .Y(
        n26670) );
  NAND2X1 U21532 ( .A(n26682), .B(n26683), .Y(n26668) );
  NOR2X1 U21533 ( .A(n26684), .B(n26685), .Y(n26683) );
  OAI21X1 U21534 ( .A(n26686), .B(n26687), .C(n26688), .Y(n26685) );
  OAI21X1 U21535 ( .A(n26689), .B(n26690), .C(reg_A[8]), .Y(n26688) );
  NAND2X1 U21536 ( .A(n25188), .B(n26691), .Y(n26687) );
  OAI21X1 U21537 ( .A(n26692), .B(n26693), .C(n26694), .Y(n26684) );
  OAI21X1 U21538 ( .A(n26695), .B(n26696), .C(n25310), .Y(n26694) );
  NAND2X1 U21539 ( .A(n26697), .B(n26698), .Y(n26696) );
  NOR2X1 U21540 ( .A(n26699), .B(n26700), .Y(n26698) );
  OAI21X1 U21541 ( .A(n26701), .B(n25043), .C(n26702), .Y(n26700) );
  AOI22X1 U21542 ( .A(n25135), .B(reg_A[9]), .C(n25252), .D(reg_A[10]), .Y(
        n26702) );
  OAI21X1 U21543 ( .A(n25206), .B(n26703), .C(n26704), .Y(n26699) );
  AOI22X1 U21544 ( .A(reg_A[11]), .B(n25136), .C(n25069), .D(reg_A[12]), .Y(
        n26704) );
  NOR2X1 U21545 ( .A(n26705), .B(n26706), .Y(n26697) );
  OAI21X1 U21546 ( .A(n25250), .B(n25467), .C(n26707), .Y(n26706) );
  AOI22X1 U21547 ( .A(reg_A[14]), .B(n25253), .C(n25628), .D(reg_A[15]), .Y(
        n26707) );
  OAI21X1 U21548 ( .A(n25224), .B(n25219), .C(n26708), .Y(n26705) );
  AOI22X1 U21549 ( .A(reg_A[17]), .B(n25629), .C(reg_A[19]), .D(n25222), .Y(
        n26708) );
  NAND2X1 U21550 ( .A(n26709), .B(n26710), .Y(n26695) );
  NOR2X1 U21551 ( .A(n26711), .B(n26712), .Y(n26710) );
  OAI21X1 U21552 ( .A(n25232), .B(n25229), .C(n26713), .Y(n26712) );
  AOI22X1 U21553 ( .A(reg_A[22]), .B(n25234), .C(n25635), .D(reg_A[20]), .Y(
        n26713) );
  OAI21X1 U21554 ( .A(n26714), .B(n25482), .C(n26715), .Y(n26711) );
  AOI22X1 U21555 ( .A(reg_A[25]), .B(n25246), .C(reg_A[24]), .D(n25247), .Y(
        n26715) );
  NOR2X1 U21556 ( .A(n26716), .B(n26717), .Y(n26709) );
  OAI21X1 U21557 ( .A(n25244), .B(n25238), .C(n26718), .Y(n26717) );
  AOI22X1 U21558 ( .A(reg_A[27]), .B(n25487), .C(n25241), .D(reg_A[26]), .Y(
        n26718) );
  OAI21X1 U21559 ( .A(n25239), .B(n26719), .C(n26720), .Y(n26716) );
  AOI22X1 U21560 ( .A(reg_A[30]), .B(n25242), .C(n25338), .D(reg_A[31]), .Y(
        n26720) );
  NAND2X1 U21561 ( .A(n25170), .B(n25171), .Y(n26693) );
  OAI21X1 U21562 ( .A(n26721), .B(n25415), .C(n26722), .Y(n25171) );
  NAND3X1 U21563 ( .A(n25589), .B(n26723), .C(reg_A[8]), .Y(n26722) );
  AOI21X1 U21564 ( .A(n26267), .B(n26724), .C(n26725), .Y(n26682) );
  OAI22X1 U21565 ( .A(n26726), .B(n26727), .C(n26728), .D(n26729), .Y(n26725)
         );
  OAI21X1 U21566 ( .A(n26730), .B(n26731), .C(n26732), .Y(n26724) );
  AOI22X1 U21567 ( .A(n26733), .B(n25160), .C(n26734), .D(n26735), .Y(n26732)
         );
  NOR2X1 U21568 ( .A(n26736), .B(n26737), .Y(n26666) );
  INVX1 U21569 ( .A(n26738), .Y(n26737) );
  AOI21X1 U21570 ( .A(n26739), .B(reg_A[11]), .C(n26740), .Y(n26738) );
  OAI22X1 U21571 ( .A(n26741), .B(n26420), .C(n26742), .D(n26743), .Y(n26740)
         );
  NAND2X1 U21572 ( .A(n26744), .B(n26745), .Y(n26736) );
  AOI22X1 U21573 ( .A(reg_A[13]), .B(n26746), .C(reg_A[14]), .D(n26747), .Y(
        n26745) );
  AOI22X1 U21574 ( .A(reg_A[15]), .B(n26748), .C(reg_A[7]), .D(n26749), .Y(
        n26744) );
  NOR2X1 U21575 ( .A(n26750), .B(n26751), .Y(n26665) );
  NAND3X1 U21576 ( .A(n26752), .B(n26753), .C(n26754), .Y(n26751) );
  NAND2X1 U21577 ( .A(n26755), .B(n26756), .Y(n26753) );
  OAI21X1 U21578 ( .A(n26757), .B(n26758), .C(n26759), .Y(n26755) );
  AOI22X1 U21579 ( .A(n25258), .B(n26760), .C(n26761), .D(n26762), .Y(n26759)
         );
  OAI21X1 U21580 ( .A(n26763), .B(n26764), .C(n25382), .Y(n26752) );
  OAI21X1 U21581 ( .A(n26765), .B(n25093), .C(n26766), .Y(n26764) );
  OAI21X1 U21582 ( .A(n26767), .B(n26768), .C(n25044), .Y(n26766) );
  OAI21X1 U21583 ( .A(n26769), .B(n25099), .C(n26770), .Y(n26768) );
  AOI22X1 U21584 ( .A(n25101), .B(n26771), .C(n26772), .D(n26773), .Y(n26770)
         );
  OAI21X1 U21585 ( .A(n26774), .B(n26775), .C(n26776), .Y(n26767) );
  AOI22X1 U21586 ( .A(n25108), .B(n26777), .C(n25103), .D(n26778), .Y(n26776)
         );
  INVX1 U21587 ( .A(n26779), .Y(n26765) );
  NOR2X1 U21588 ( .A(n26780), .B(n25112), .Y(n26763) );
  OAI21X1 U21589 ( .A(n26781), .B(n25146), .C(n26782), .Y(n26750) );
  AOI22X1 U21590 ( .A(n25156), .B(n25143), .C(reg_A[10]), .D(n26783), .Y(
        n26782) );
  OR2X1 U21591 ( .A(n26784), .B(n26785), .Y(result[89]) );
  NAND3X1 U21592 ( .A(n26786), .B(n26787), .C(n26788), .Y(n26785) );
  NOR2X1 U21593 ( .A(n26789), .B(n26790), .Y(n26788) );
  OAI21X1 U21594 ( .A(n26195), .B(n26791), .C(n26792), .Y(n26790) );
  AOI22X1 U21595 ( .A(n26793), .B(n25972), .C(n25918), .D(n26794), .Y(n26792)
         );
  NAND3X1 U21596 ( .A(n26795), .B(n26796), .C(n26797), .Y(n26794) );
  NOR2X1 U21597 ( .A(n26798), .B(n26799), .Y(n26797) );
  OAI22X1 U21598 ( .A(n26800), .B(n26230), .C(n26801), .D(n26215), .Y(n26799)
         );
  OAI21X1 U21599 ( .A(n25062), .B(n25965), .C(n26802), .Y(n26798) );
  AOI22X1 U21600 ( .A(reg_A[88]), .B(n26803), .C(reg_A[86]), .D(n26804), .Y(
        n26802) );
  AOI22X1 U21601 ( .A(reg_A[80]), .B(n25614), .C(reg_A[81]), .D(n25615), .Y(
        n26796) );
  INVX1 U21602 ( .A(n26805), .Y(n26795) );
  OAI21X1 U21603 ( .A(n25929), .B(n25736), .C(n26806), .Y(n26805) );
  OAI21X1 U21604 ( .A(n26181), .B(n26807), .C(n26808), .Y(n26789) );
  AOI22X1 U21605 ( .A(n26809), .B(n26260), .C(n26349), .D(reg_A[74]), .Y(
        n26808) );
  INVX1 U21606 ( .A(n25903), .Y(n26181) );
  AOI21X1 U21607 ( .A(n26810), .B(n26014), .C(n26811), .Y(n26787) );
  OAI22X1 U21608 ( .A(n26068), .B(n26136), .C(n25973), .D(n26812), .Y(n26811)
         );
  AOI21X1 U21609 ( .A(n26655), .B(n26028), .C(n26813), .Y(n26786) );
  OAI21X1 U21610 ( .A(n25886), .B(n26575), .C(n26814), .Y(n26813) );
  OAI21X1 U21611 ( .A(n26815), .B(n26816), .C(n25840), .Y(n26814) );
  NAND2X1 U21612 ( .A(n26817), .B(n26818), .Y(n26816) );
  NOR2X1 U21613 ( .A(n26819), .B(n26820), .Y(n26818) );
  OAI21X1 U21614 ( .A(n25034), .B(n26094), .C(n26821), .Y(n26820) );
  AOI22X1 U21615 ( .A(reg_A[84]), .B(n25123), .C(reg_A[80]), .D(n25629), .Y(
        n26821) );
  OAI21X1 U21616 ( .A(n25056), .B(n26215), .C(n26822), .Y(n26819) );
  AOI22X1 U21617 ( .A(reg_A[83]), .B(n25253), .C(reg_A[82]), .D(n25628), .Y(
        n26822) );
  NOR2X1 U21618 ( .A(n26823), .B(n26824), .Y(n26817) );
  OAI21X1 U21619 ( .A(n25043), .B(n25929), .C(n26825), .Y(n26824) );
  AOI22X1 U21620 ( .A(reg_A[77]), .B(n25635), .C(reg_A[76]), .D(n25325), .Y(
        n26825) );
  OAI21X1 U21621 ( .A(n25035), .B(n26103), .C(n26826), .Y(n26823) );
  AOI22X1 U21622 ( .A(reg_A[78]), .B(n25222), .C(reg_A[79]), .D(n25637), .Y(
        n26826) );
  NAND3X1 U21623 ( .A(n26827), .B(n26828), .C(n26829), .Y(n26815) );
  NOR2X1 U21624 ( .A(n26830), .B(n26831), .Y(n26829) );
  OAI21X1 U21625 ( .A(n25040), .B(n25965), .C(n26832), .Y(n26831) );
  AOI22X1 U21626 ( .A(reg_A[88]), .B(n25135), .C(reg_A[86]), .D(n25136), .Y(
        n26832) );
  OAI21X1 U21627 ( .A(n25057), .B(n25855), .C(n26833), .Y(n26830) );
  AOI22X1 U21628 ( .A(reg_A[68]), .B(n25257), .C(reg_A[64]), .D(n25857), .Y(
        n26833) );
  NOR2X1 U21629 ( .A(n26834), .B(n26835), .Y(n26828) );
  OAI22X1 U21630 ( .A(n25051), .B(n26101), .C(n25243), .D(n26256), .Y(n26835)
         );
  OAI22X1 U21631 ( .A(n25334), .B(n26439), .C(n25336), .D(n26547), .Y(n26834)
         );
  AOI21X1 U21632 ( .A(reg_A[69]), .B(n25339), .C(n26836), .Y(n26827) );
  OAI22X1 U21633 ( .A(n25491), .B(n25884), .C(n25492), .D(n25851), .Y(n26836)
         );
  NAND2X1 U21634 ( .A(n26837), .B(n26838), .Y(n26575) );
  AOI22X1 U21635 ( .A(n25838), .B(n26305), .C(n26160), .D(n26839), .Y(n26838)
         );
  INVX1 U21636 ( .A(n26300), .Y(n26839) );
  NAND2X1 U21637 ( .A(n26840), .B(n26841), .Y(n26305) );
  AOI22X1 U21638 ( .A(n26061), .B(n25855), .C(n26513), .D(n26439), .Y(n26841)
         );
  AOI22X1 U21639 ( .A(n26134), .B(n25929), .C(n25892), .D(n26094), .Y(n26840)
         );
  INVX1 U21640 ( .A(n26842), .Y(n26837) );
  OAI22X1 U21641 ( .A(n25898), .B(n26514), .C(n26112), .D(n26843), .Y(n26842)
         );
  AND2X1 U21642 ( .A(n26844), .B(n26845), .Y(n26655) );
  AOI22X1 U21643 ( .A(n25025), .B(n26531), .C(n25026), .D(n26529), .Y(n26845)
         );
  AOI22X1 U21644 ( .A(n26032), .B(n26213), .C(n26530), .D(n26846), .Y(n26844)
         );
  NAND2X1 U21645 ( .A(n26847), .B(n26848), .Y(n26213) );
  AOI22X1 U21646 ( .A(n26662), .B(n25855), .C(n26663), .D(n26439), .Y(n26848)
         );
  AOI22X1 U21647 ( .A(n26038), .B(n26094), .C(n26664), .D(n25929), .Y(n26847)
         );
  NAND3X1 U21648 ( .A(n26849), .B(n26850), .C(n26851), .Y(n26784) );
  NOR2X1 U21649 ( .A(n26852), .B(n26853), .Y(n26851) );
  OAI21X1 U21650 ( .A(n26854), .B(n26550), .C(n26855), .Y(n26853) );
  AOI22X1 U21651 ( .A(n26148), .B(n26856), .C(n26451), .D(reg_A[92]), .Y(
        n26855) );
  NAND2X1 U21652 ( .A(n26857), .B(n26858), .Y(n26550) );
  AOI22X1 U21653 ( .A(n26859), .B(n26230), .C(n26860), .D(n26215), .Y(n26858)
         );
  AOI22X1 U21654 ( .A(n26455), .B(n25584), .C(n26316), .D(n26452), .Y(n26857)
         );
  OAI21X1 U21655 ( .A(reg_A[80]), .B(n26861), .C(n26862), .Y(n26316) );
  AOI22X1 U21656 ( .A(n26598), .B(n26863), .C(n26462), .D(n26195), .Y(n26862)
         );
  MUX2X1 U21657 ( .B(reg_A[81]), .A(reg_A[89]), .S(n26596), .Y(n26598) );
  OAI21X1 U21658 ( .A(n26806), .B(n26864), .C(n26865), .Y(n26852) );
  AOI22X1 U21659 ( .A(n26866), .B(reg_A[80]), .C(n25188), .D(n26867), .Y(
        n26865) );
  NAND2X1 U21660 ( .A(n26868), .B(n26869), .Y(n26867) );
  AOI22X1 U21661 ( .A(n26870), .B(n25891), .C(n26871), .D(n26276), .Y(n26869)
         );
  MUX2X1 U21662 ( .B(n25965), .A(n26039), .S(reg_B[95]), .Y(n25891) );
  INVX1 U21663 ( .A(n26872), .Y(n26870) );
  AOI21X1 U21664 ( .A(n26474), .B(n25950), .C(n26873), .Y(n26868) );
  MUX2X1 U21665 ( .B(n26874), .A(n26875), .S(reg_B[92]), .Y(n26873) );
  NAND2X1 U21666 ( .A(reg_B[94]), .B(reg_A[80]), .Y(n26875) );
  NAND3X1 U21667 ( .A(reg_B[95]), .B(reg_A[82]), .C(n26159), .Y(n26874) );
  AOI21X1 U21668 ( .A(n25584), .B(n25989), .C(n26876), .Y(n26474) );
  OAI22X1 U21669 ( .A(n26069), .B(n26198), .C(n26196), .D(reg_B[93]), .Y(
        n26876) );
  MUX2X1 U21670 ( .B(n26566), .A(n26877), .S(reg_B[95]), .Y(n26196) );
  MUX2X1 U21671 ( .B(reg_A[88]), .A(reg_A[80]), .S(reg_B[92]), .Y(n26877) );
  MUX2X1 U21672 ( .B(reg_A[81]), .A(reg_A[89]), .S(n26063), .Y(n26566) );
  MUX2X1 U21673 ( .B(n26215), .A(n26230), .S(reg_B[95]), .Y(n26198) );
  AOI22X1 U21674 ( .A(n25613), .B(reg_A[82]), .C(n26878), .D(reg_A[83]), .Y(
        n26806) );
  NOR2X1 U21675 ( .A(n26879), .B(n26880), .Y(n26850) );
  OAI21X1 U21676 ( .A(n26881), .B(n26457), .C(n26882), .Y(n26880) );
  OAI21X1 U21677 ( .A(n26397), .B(n26883), .C(reg_A[89]), .Y(n26882) );
  NOR2X1 U21678 ( .A(n26394), .B(n25972), .Y(n26397) );
  NAND2X1 U21679 ( .A(n26504), .B(n26197), .Y(n26394) );
  INVX1 U21680 ( .A(n25936), .Y(n26457) );
  OAI21X1 U21681 ( .A(n26884), .B(n26147), .C(n26391), .Y(n26879) );
  NAND2X1 U21682 ( .A(n26793), .B(reg_B[93]), .Y(n26391) );
  INVX1 U21683 ( .A(n26111), .Y(n26793) );
  NAND2X1 U21684 ( .A(reg_A[88]), .B(n26504), .Y(n26111) );
  AOI22X1 U21685 ( .A(n26276), .B(n26885), .C(n26149), .D(n26886), .Y(n26884)
         );
  AOI21X1 U21686 ( .A(n25170), .B(n26887), .C(n26888), .Y(n26849) );
  OAI21X1 U21687 ( .A(n26182), .B(n26889), .C(n26890), .Y(n26888) );
  OAI21X1 U21688 ( .A(n26891), .B(n26892), .C(n25203), .Y(n26890) );
  OAI22X1 U21689 ( .A(n26893), .B(n25883), .C(n26894), .D(n25873), .Y(n26892)
         );
  NOR2X1 U21690 ( .A(n26895), .B(n25881), .Y(n26891) );
  INVX1 U21691 ( .A(n26603), .Y(n26889) );
  OAI21X1 U21692 ( .A(n26582), .B(n26896), .C(n26897), .Y(n26887) );
  AOI22X1 U21693 ( .A(n25980), .B(n26898), .C(n25984), .D(n26590), .Y(n26897)
         );
  OAI21X1 U21694 ( .A(n26899), .B(n25415), .C(n26900), .Y(n26590) );
  NAND3X1 U21695 ( .A(n25589), .B(n26197), .C(reg_A[89]), .Y(n26900) );
  INVX1 U21696 ( .A(n26402), .Y(n26899) );
  OAI21X1 U21697 ( .A(n26067), .B(n25929), .C(n26901), .Y(n26402) );
  AOI22X1 U21698 ( .A(reg_A[81]), .B(n25988), .C(n26274), .D(reg_A[85]), .Y(
        n26901) );
  AND2X1 U21699 ( .A(n26902), .B(n26903), .Y(n26582) );
  AOI22X1 U21700 ( .A(n25838), .B(n26288), .C(n26160), .D(n26289), .Y(n26903)
         );
  NAND2X1 U21701 ( .A(n26904), .B(n26905), .Y(n26288) );
  AOI22X1 U21702 ( .A(reg_A[65]), .B(n26061), .C(reg_A[73]), .D(n26513), .Y(
        n26905) );
  AOI22X1 U21703 ( .A(reg_A[89]), .B(n26134), .C(reg_A[81]), .D(n25892), .Y(
        n26904) );
  AOI22X1 U21704 ( .A(n26059), .B(n26510), .C(n26159), .D(n26906), .Y(n26902)
         );
  NAND3X1 U21705 ( .A(n26907), .B(n26908), .C(n26909), .Y(result[88]) );
  NOR2X1 U21706 ( .A(n26910), .B(n26911), .Y(n26909) );
  NAND3X1 U21707 ( .A(n26912), .B(n26913), .C(n26914), .Y(n26911) );
  AOI21X1 U21708 ( .A(n26915), .B(n25903), .C(n26916), .Y(n26914) );
  OAI22X1 U21709 ( .A(n26439), .B(n26625), .C(n25863), .D(n26917), .Y(n26916)
         );
  OAI21X1 U21710 ( .A(n25087), .B(n26918), .C(n26919), .Y(n25903) );
  NAND2X1 U21711 ( .A(n25974), .B(n26197), .Y(n26918) );
  OAI21X1 U21712 ( .A(n26920), .B(n26921), .C(n25730), .Y(n26913) );
  NAND2X1 U21713 ( .A(n26922), .B(n26923), .Y(n26921) );
  AOI22X1 U21714 ( .A(reg_A[95]), .B(n25613), .C(reg_A[92]), .D(n25749), .Y(
        n26923) );
  AOI22X1 U21715 ( .A(reg_A[93]), .B(n25750), .C(reg_A[88]), .D(n26924), .Y(
        n26922) );
  NAND2X1 U21716 ( .A(n26925), .B(n26926), .Y(n26920) );
  AOI22X1 U21717 ( .A(reg_A[89]), .B(n26803), .C(reg_A[91]), .D(n26804), .Y(
        n26926) );
  AOI22X1 U21718 ( .A(reg_A[90]), .B(n26927), .C(reg_A[94]), .D(n26878), .Y(
        n26925) );
  AOI22X1 U21719 ( .A(n26928), .B(n26929), .C(n25918), .D(n26930), .Y(n26912)
         );
  NAND3X1 U21720 ( .A(n26931), .B(n26932), .C(n26933), .Y(n26930) );
  NOR2X1 U21721 ( .A(n26934), .B(n26935), .Y(n26933) );
  OAI22X1 U21722 ( .A(n26936), .B(n26094), .C(n25745), .D(n25874), .Y(n26935)
         );
  OAI21X1 U21723 ( .A(n25062), .B(n26039), .C(n26937), .Y(n26934) );
  AOI22X1 U21724 ( .A(reg_A[87]), .B(n26803), .C(reg_A[85]), .D(n26804), .Y(
        n26937) );
  AOI22X1 U21725 ( .A(reg_A[84]), .B(n25749), .C(reg_A[83]), .D(n25750), .Y(
        n26932) );
  AOI22X1 U21726 ( .A(reg_A[80]), .B(n25615), .C(reg_A[88]), .D(n26924), .Y(
        n26931) );
  NAND3X1 U21727 ( .A(n26938), .B(n26939), .C(n26940), .Y(n26929) );
  NOR2X1 U21728 ( .A(n26941), .B(n26942), .Y(n26940) );
  OAI22X1 U21729 ( .A(n26943), .B(n26195), .C(n26944), .D(n25881), .Y(n26942)
         );
  OAI22X1 U21730 ( .A(n26945), .B(n25882), .C(n25753), .D(n25873), .Y(n26941)
         );
  AOI22X1 U21731 ( .A(reg_A[89]), .B(n26007), .C(reg_A[91]), .D(n26008), .Y(
        n26939) );
  AOI22X1 U21732 ( .A(reg_A[90]), .B(n26009), .C(reg_A[94]), .D(n26010), .Y(
        n26938) );
  NAND2X1 U21733 ( .A(n26946), .B(n26947), .Y(n26910) );
  AOI21X1 U21734 ( .A(n26809), .B(n26028), .C(n26948), .Y(n26947) );
  OAI21X1 U21735 ( .A(n26949), .B(n26950), .C(n26951), .Y(n26948) );
  OAI21X1 U21736 ( .A(n26952), .B(n26953), .C(n25840), .Y(n26951) );
  NAND3X1 U21737 ( .A(n26954), .B(n26955), .C(n26956), .Y(n26953) );
  NOR2X1 U21738 ( .A(n26957), .B(n26958), .Y(n26956) );
  OAI21X1 U21739 ( .A(n25037), .B(n25864), .C(n26959), .Y(n26958) );
  AOI22X1 U21740 ( .A(reg_A[84]), .B(n25071), .C(reg_A[83]), .D(n25123), .Y(
        n26959) );
  OAI21X1 U21741 ( .A(n25030), .B(n26094), .C(n26960), .Y(n26957) );
  AOI22X1 U21742 ( .A(reg_A[86]), .B(n25252), .C(reg_A[82]), .D(n25253), .Y(
        n26960) );
  AOI21X1 U21743 ( .A(reg_A[74]), .B(n25234), .C(n26961), .Y(n26955) );
  OAI22X1 U21744 ( .A(n25036), .B(n25865), .C(n25467), .D(n25584), .Y(n26961)
         );
  AOI22X1 U21745 ( .A(reg_A[75]), .B(n25325), .C(reg_A[88]), .D(n25125), .Y(
        n26954) );
  NAND3X1 U21746 ( .A(n26962), .B(n26963), .C(n26964), .Y(n26952) );
  NOR2X1 U21747 ( .A(n26965), .B(n26966), .Y(n26964) );
  OAI21X1 U21748 ( .A(n25491), .B(n25855), .C(n26967), .Y(n26966) );
  AOI22X1 U21749 ( .A(reg_A[70]), .B(n25241), .C(reg_A[66]), .D(n25242), .Y(
        n26967) );
  OAI21X1 U21750 ( .A(n25038), .B(n25856), .C(n26968), .Y(n26965) );
  AOI22X1 U21751 ( .A(reg_A[71]), .B(n25246), .C(reg_A[72]), .D(n25247), .Y(
        n26968) );
  AOI21X1 U21752 ( .A(reg_A[64]), .B(n25647), .C(n26969), .Y(n26963) );
  OAI22X1 U21753 ( .A(n26719), .B(n25851), .C(n25238), .D(n26107), .Y(n26969)
         );
  AOI22X1 U21754 ( .A(reg_A[87]), .B(n25135), .C(reg_A[85]), .D(n25136), .Y(
        n26962) );
  INVX1 U21755 ( .A(n26898), .Y(n26949) );
  NAND2X1 U21756 ( .A(n26970), .B(n26971), .Y(n26898) );
  AOI22X1 U21757 ( .A(n25838), .B(n26345), .C(n26160), .D(n26339), .Y(n26971)
         );
  NAND2X1 U21758 ( .A(n26972), .B(n26973), .Y(n26345) );
  AOI22X1 U21759 ( .A(reg_A[72]), .B(n26513), .C(reg_A[88]), .D(n26134), .Y(
        n26973) );
  AOI22X1 U21760 ( .A(n26974), .B(reg_B[91]), .C(n25892), .D(reg_A[80]), .Y(
        n26972) );
  AOI22X1 U21761 ( .A(n26059), .B(n26611), .C(n26159), .D(n26975), .Y(n26970)
         );
  AND2X1 U21762 ( .A(n26976), .B(n26977), .Y(n26809) );
  AOI22X1 U21763 ( .A(n25025), .B(n26659), .C(n25026), .D(n26658), .Y(n26977)
         );
  AOI22X1 U21764 ( .A(n26032), .B(n26365), .C(n26530), .D(n26978), .Y(n26976)
         );
  OR2X1 U21765 ( .A(n26979), .B(n26980), .Y(n26365) );
  OAI22X1 U21766 ( .A(reg_A[88]), .B(n26036), .C(reg_A[80]), .D(n26981), .Y(
        n26980) );
  OAI21X1 U21767 ( .A(reg_A[72]), .B(n26982), .C(n26983), .Y(n26979) );
  AOI21X1 U21768 ( .A(n26627), .B(reg_A[77]), .C(n26984), .Y(n26946) );
  OAI22X1 U21769 ( .A(n26985), .B(n25584), .C(n26012), .D(n26986), .Y(n26984)
         );
  NOR2X1 U21770 ( .A(n26987), .B(n26988), .Y(n26908) );
  OAI21X1 U21771 ( .A(n26989), .B(n26990), .C(n26991), .Y(n26988) );
  AOI22X1 U21772 ( .A(n26603), .B(n26992), .C(n26267), .D(n26993), .Y(n26991)
         );
  OAI21X1 U21773 ( .A(n26994), .B(n26169), .C(n26995), .Y(n26993) );
  AOI22X1 U21774 ( .A(n26148), .B(n26885), .C(n26276), .D(n26886), .Y(n26995)
         );
  OAI21X1 U21775 ( .A(n26996), .B(n26997), .C(n26998), .Y(n26603) );
  NAND3X1 U21776 ( .A(n25382), .B(n25974), .C(reg_B[93]), .Y(n26998) );
  OAI21X1 U21777 ( .A(reg_B[92]), .B(n25415), .C(n26999), .Y(n25974) );
  NOR2X1 U21778 ( .A(n27000), .B(n27001), .Y(n26989) );
  OAI21X1 U21779 ( .A(n25028), .B(n25881), .C(n27002), .Y(n27001) );
  AOI22X1 U21780 ( .A(reg_A[95]), .B(n25628), .C(reg_A[92]), .D(n25066), .Y(
        n27002) );
  NAND2X1 U21781 ( .A(n27003), .B(n27004), .Y(n27000) );
  AOI22X1 U21782 ( .A(reg_A[89]), .B(n25135), .C(reg_A[91]), .D(n25136), .Y(
        n27004) );
  AOI22X1 U21783 ( .A(reg_A[90]), .B(n25252), .C(reg_A[94]), .D(n25253), .Y(
        n27003) );
  NAND3X1 U21784 ( .A(n27005), .B(n27006), .C(n27007), .Y(n26987) );
  AOI22X1 U21785 ( .A(n26396), .B(n26380), .C(n27008), .D(n27009), .Y(n27007)
         );
  INVX1 U21786 ( .A(n26419), .Y(n27009) );
  NAND2X1 U21787 ( .A(n27010), .B(n27011), .Y(n26419) );
  AOI22X1 U21788 ( .A(n26601), .B(n26039), .C(n26602), .D(n26215), .Y(n27011)
         );
  AOI22X1 U21789 ( .A(n27012), .B(n26195), .C(n26597), .D(n25965), .Y(n27010)
         );
  AND2X1 U21790 ( .A(n27013), .B(n27014), .Y(n26380) );
  AOI22X1 U21791 ( .A(n26276), .B(n26039), .C(n26149), .D(n26215), .Y(n27014)
         );
  AOI22X1 U21792 ( .A(n26148), .B(n25965), .C(n25984), .D(n26195), .Y(n27013)
         );
  NAND3X1 U21793 ( .A(n26274), .B(n25188), .C(n26379), .Y(n27005) );
  AND2X1 U21794 ( .A(n27015), .B(n27016), .Y(n26379) );
  AOI22X1 U21795 ( .A(n26276), .B(n25874), .C(n26149), .D(n26094), .Y(n27016)
         );
  AOI22X1 U21796 ( .A(n26148), .B(n25875), .C(n25984), .D(n26230), .Y(n27015)
         );
  NOR2X1 U21797 ( .A(n27017), .B(n27018), .Y(n26907) );
  OAI21X1 U21798 ( .A(n27019), .B(n27020), .C(n27021), .Y(n27018) );
  AOI22X1 U21799 ( .A(n27022), .B(n26014), .C(n26810), .D(n26125), .Y(n27021)
         );
  AND2X1 U21800 ( .A(n27023), .B(n27024), .Y(n26810) );
  AOI22X1 U21801 ( .A(n25838), .B(n26414), .C(n26160), .D(n26653), .Y(n27024)
         );
  OR2X1 U21802 ( .A(n27025), .B(n27026), .Y(n26414) );
  OAI22X1 U21803 ( .A(reg_A[80]), .B(n26131), .C(reg_A[88]), .D(n25894), .Y(
        n27026) );
  OAI21X1 U21804 ( .A(reg_A[72]), .B(n27027), .C(n27028), .Y(n27025) );
  AOI22X1 U21805 ( .A(n26059), .B(n26654), .C(n26159), .D(n27029), .Y(n27023)
         );
  INVX1 U21806 ( .A(n27030), .Y(n27019) );
  OAI21X1 U21807 ( .A(n26422), .B(n26420), .C(n27031), .Y(n27017) );
  AOI22X1 U21808 ( .A(n25984), .B(n26856), .C(reg_A[88]), .D(n27032), .Y(
        n27031) );
  OAI21X1 U21809 ( .A(n27033), .B(n26147), .C(n27034), .Y(n26856) );
  NAND3X1 U21810 ( .A(n26186), .B(n26197), .C(reg_A[88]), .Y(n27034) );
  INVX1 U21811 ( .A(n26489), .Y(n27033) );
  OAI21X1 U21812 ( .A(n26067), .B(n26195), .C(n27035), .Y(n26489) );
  AOI22X1 U21813 ( .A(n25988), .B(reg_A[80]), .C(n26274), .D(reg_A[84]), .Y(
        n27035) );
  NAND3X1 U21814 ( .A(n27036), .B(n27037), .C(n27038), .Y(result[87]) );
  AND2X1 U21815 ( .A(n27039), .B(n27040), .Y(n27038) );
  NOR2X1 U21816 ( .A(n27041), .B(n27042), .Y(n27040) );
  NAND2X1 U21817 ( .A(n27043), .B(n27044), .Y(n27042) );
  OAI21X1 U21818 ( .A(n27045), .B(n27046), .C(reg_A[87]), .Y(n27044) );
  AOI22X1 U21819 ( .A(n25170), .B(n27047), .C(reg_A[80]), .D(n27048), .Y(
        n27043) );
  OAI21X1 U21820 ( .A(n26169), .B(n27049), .C(n27050), .Y(n27048) );
  INVX1 U21821 ( .A(n27051), .Y(n27050) );
  NAND2X1 U21822 ( .A(reg_B[93]), .B(n25188), .Y(n27049) );
  OAI21X1 U21823 ( .A(n27052), .B(n27053), .C(n27054), .Y(n27047) );
  OAI21X1 U21824 ( .A(n27055), .B(n27056), .C(n27057), .Y(n27054) );
  OAI22X1 U21825 ( .A(n25965), .B(n27058), .C(n27059), .D(n27060), .Y(n27056)
         );
  MUX2X1 U21826 ( .B(reg_A[83]), .A(reg_A[81]), .S(reg_B[86]), .Y(n27060) );
  NOR2X1 U21827 ( .A(n26215), .B(n27061), .Y(n27055) );
  INVX1 U21828 ( .A(n27062), .Y(n27052) );
  NAND3X1 U21829 ( .A(n27063), .B(n27006), .C(n27064), .Y(n27041) );
  OAI21X1 U21830 ( .A(n27065), .B(n27066), .C(n27067), .Y(n27064) );
  OAI21X1 U21831 ( .A(n25060), .B(n25965), .C(n27068), .Y(n27066) );
  AOI22X1 U21832 ( .A(reg_A[83]), .B(n25749), .C(reg_A[82]), .D(n25750), .Y(
        n27068) );
  NAND2X1 U21833 ( .A(n27069), .B(n27070), .Y(n27065) );
  AOI22X1 U21834 ( .A(reg_A[86]), .B(n26803), .C(reg_A[84]), .D(n26804), .Y(
        n27070) );
  AOI22X1 U21835 ( .A(reg_A[85]), .B(n26927), .C(reg_A[81]), .D(n26878), .Y(
        n27069) );
  NAND2X1 U21836 ( .A(n25890), .B(reg_A[80]), .Y(n27006) );
  OAI21X1 U21837 ( .A(n27071), .B(n27072), .C(n25840), .Y(n27063) );
  NAND2X1 U21838 ( .A(n27073), .B(n27074), .Y(n27072) );
  NOR2X1 U21839 ( .A(n27075), .B(n27076), .Y(n27074) );
  OAI21X1 U21840 ( .A(n25043), .B(n25965), .C(n27077), .Y(n27076) );
  AOI22X1 U21841 ( .A(reg_A[86]), .B(n25135), .C(reg_A[85]), .D(n25252), .Y(
        n27077) );
  OAI21X1 U21842 ( .A(n25028), .B(n25874), .C(n27078), .Y(n27075) );
  AOI22X1 U21843 ( .A(reg_A[84]), .B(n25136), .C(reg_A[83]), .D(n25066), .Y(
        n27078) );
  NOR2X1 U21844 ( .A(n27079), .B(n27080), .Y(n27073) );
  OAI21X1 U21845 ( .A(n25034), .B(n25864), .C(n27081), .Y(n27080) );
  AOI22X1 U21846 ( .A(reg_A[81]), .B(n25253), .C(reg_A[80]), .D(n25628), .Y(
        n27081) );
  OAI21X1 U21847 ( .A(n25036), .B(n26286), .C(n27082), .Y(n27079) );
  AOI22X1 U21848 ( .A(reg_A[78]), .B(n25629), .C(reg_A[76]), .D(n25222), .Y(
        n27082) );
  NAND2X1 U21849 ( .A(n27083), .B(n27084), .Y(n27071) );
  NOR2X1 U21850 ( .A(n27085), .B(n27086), .Y(n27084) );
  OAI21X1 U21851 ( .A(n25039), .B(n26438), .C(n27087), .Y(n27086) );
  AOI22X1 U21852 ( .A(reg_A[73]), .B(n25234), .C(reg_A[75]), .D(n25635), .Y(
        n27087) );
  OAI21X1 U21853 ( .A(n25065), .B(n26547), .C(n27088), .Y(n27085) );
  AOI22X1 U21854 ( .A(reg_A[70]), .B(n25246), .C(reg_A[71]), .D(n25247), .Y(
        n27088) );
  NOR2X1 U21855 ( .A(n27089), .B(n27090), .Y(n27083) );
  OAI21X1 U21856 ( .A(n25238), .B(n25851), .C(n27091), .Y(n27090) );
  AOI22X1 U21857 ( .A(reg_A[68]), .B(n25487), .C(reg_A[69]), .D(n25241), .Y(
        n27091) );
  OAI21X1 U21858 ( .A(n26719), .B(n25884), .C(n27092), .Y(n27089) );
  AOI22X1 U21859 ( .A(reg_A[65]), .B(n25242), .C(reg_A[64]), .D(n25338), .Y(
        n27092) );
  NOR2X1 U21860 ( .A(n27093), .B(n27094), .Y(n27039) );
  OAI21X1 U21861 ( .A(n26230), .B(n27095), .C(n27096), .Y(n27094) );
  AOI22X1 U21862 ( .A(n25999), .B(n27097), .C(n26504), .D(n27098), .Y(n27096)
         );
  NAND2X1 U21863 ( .A(n27099), .B(n27100), .Y(n27098) );
  AOI22X1 U21864 ( .A(n27101), .B(n27102), .C(n27103), .D(n27104), .Y(n27100)
         );
  AOI22X1 U21865 ( .A(reg_B[87]), .B(n27105), .C(n27106), .D(reg_B[86]), .Y(
        n27099) );
  OAI21X1 U21866 ( .A(n25754), .B(n26094), .C(n27107), .Y(n27097) );
  AOI22X1 U21867 ( .A(reg_A[86]), .B(n26007), .C(reg_A[85]), .D(n26009), .Y(
        n27107) );
  OAI21X1 U21868 ( .A(n25874), .B(n27108), .C(n27109), .Y(n27093) );
  AOI22X1 U21869 ( .A(n26281), .B(n27030), .C(n27110), .D(n25936), .Y(n27109)
         );
  MUX2X1 U21870 ( .B(n25965), .A(n26039), .S(reg_B[4]), .Y(n25936) );
  NAND2X1 U21871 ( .A(n27111), .B(n27112), .Y(n27030) );
  AOI22X1 U21872 ( .A(n25838), .B(n26289), .C(n26160), .D(n26510), .Y(n27112)
         );
  OAI21X1 U21873 ( .A(n26131), .B(n25864), .C(n27113), .Y(n26289) );
  AOI22X1 U21874 ( .A(reg_A[71]), .B(n26513), .C(reg_A[87]), .D(n26134), .Y(
        n27113) );
  AOI22X1 U21875 ( .A(n26059), .B(n26906), .C(n26159), .D(n27114), .Y(n27111)
         );
  NOR2X1 U21876 ( .A(n27115), .B(n27116), .Y(n27037) );
  OAI21X1 U21877 ( .A(n26525), .B(n26986), .C(n27117), .Y(n27116) );
  AOI22X1 U21878 ( .A(n27118), .B(n26014), .C(n27022), .D(n26125), .Y(n27117)
         );
  NOR2X1 U21879 ( .A(n27119), .B(n27120), .Y(n27022) );
  OAI22X1 U21880 ( .A(n26337), .B(n26300), .C(n26338), .D(n26514), .Y(n27120)
         );
  NOR2X1 U21881 ( .A(n27121), .B(n27122), .Y(n26300) );
  OAI22X1 U21882 ( .A(reg_A[79]), .B(n26131), .C(reg_A[87]), .D(n25894), .Y(
        n27122) );
  OAI21X1 U21883 ( .A(reg_A[71]), .B(n27027), .C(n27028), .Y(n27121) );
  OAI22X1 U21884 ( .A(n25898), .B(n26843), .C(n26112), .D(n27123), .Y(n27119)
         );
  NAND2X1 U21885 ( .A(n27124), .B(n27125), .Y(n26986) );
  AOI22X1 U21886 ( .A(n25025), .B(n26846), .C(n25026), .D(n26531), .Y(n27125)
         );
  INVX1 U21887 ( .A(n27126), .Y(n26846) );
  AOI22X1 U21888 ( .A(n26032), .B(n26529), .C(n26530), .D(n27127), .Y(n27124)
         );
  INVX1 U21889 ( .A(n26207), .Y(n26529) );
  NOR2X1 U21890 ( .A(n27128), .B(n27129), .Y(n26207) );
  OAI22X1 U21891 ( .A(reg_A[87]), .B(n26036), .C(reg_A[79]), .D(n26981), .Y(
        n27129) );
  OAI21X1 U21892 ( .A(reg_A[71]), .B(n26982), .C(n26983), .Y(n27128) );
  OAI21X1 U21893 ( .A(n25945), .B(n27130), .C(n27131), .Y(n27115) );
  AOI22X1 U21894 ( .A(n27132), .B(reg_A[83]), .C(n26149), .D(n27133), .Y(
        n27131) );
  INVX1 U21895 ( .A(n27134), .Y(n27133) );
  NOR2X1 U21896 ( .A(n27135), .B(n27136), .Y(n27036) );
  OAI21X1 U21897 ( .A(n27137), .B(n27138), .C(n27139), .Y(n27136) );
  AOI22X1 U21898 ( .A(n25310), .B(n27140), .C(n27141), .D(n27142), .Y(n27139)
         );
  NAND3X1 U21899 ( .A(n27143), .B(n27144), .C(n27145), .Y(n27140) );
  NOR2X1 U21900 ( .A(n27146), .B(n27147), .Y(n27145) );
  OAI22X1 U21901 ( .A(n25030), .B(n25883), .C(n25131), .D(n25881), .Y(n27147)
         );
  OAI21X1 U21902 ( .A(n25040), .B(n25929), .C(n27148), .Y(n27146) );
  AOI22X1 U21903 ( .A(reg_A[88]), .B(n25135), .C(reg_A[90]), .D(n25136), .Y(
        n27148) );
  AOI22X1 U21904 ( .A(reg_A[91]), .B(n25070), .C(reg_A[92]), .D(n25123), .Y(
        n27144) );
  AOI22X1 U21905 ( .A(reg_A[95]), .B(n25124), .C(reg_A[87]), .D(n25125), .Y(
        n27143) );
  INVX1 U21906 ( .A(n27149), .Y(n27138) );
  INVX1 U21907 ( .A(n27150), .Y(n27137) );
  OAI21X1 U21908 ( .A(n27151), .B(n27152), .C(n27153), .Y(n27135) );
  AOI22X1 U21909 ( .A(n27154), .B(n26260), .C(n27155), .D(n27156), .Y(n27153)
         );
  OAI21X1 U21910 ( .A(n26994), .B(n25914), .C(n27157), .Y(n27156) );
  AOI22X1 U21911 ( .A(n25984), .B(n26885), .C(n26148), .D(n26886), .Y(n27157)
         );
  INVX1 U21912 ( .A(n26614), .Y(n26885) );
  AOI21X1 U21913 ( .A(n26275), .B(reg_A[87]), .C(n26871), .Y(n26614) );
  NOR2X1 U21914 ( .A(n26069), .B(n25875), .Y(n26871) );
  INVX1 U21915 ( .A(n27158), .Y(n27154) );
  INVX1 U21916 ( .A(n27159), .Y(n27151) );
  NAND3X1 U21917 ( .A(n27160), .B(n27161), .C(n27162), .Y(n27159) );
  NOR2X1 U21918 ( .A(n27163), .B(n27164), .Y(n27162) );
  OAI22X1 U21919 ( .A(n26936), .B(n25883), .C(n25745), .D(n25881), .Y(n27164)
         );
  OAI21X1 U21920 ( .A(n25062), .B(n25929), .C(n27165), .Y(n27163) );
  AOI22X1 U21921 ( .A(reg_A[88]), .B(n26803), .C(reg_A[90]), .D(n26804), .Y(
        n27165) );
  AOI22X1 U21922 ( .A(reg_A[91]), .B(n25749), .C(reg_A[92]), .D(n25750), .Y(
        n27161) );
  AOI22X1 U21923 ( .A(reg_A[95]), .B(n25615), .C(reg_A[87]), .D(n26924), .Y(
        n27160) );
  NAND3X1 U21924 ( .A(n27166), .B(n27167), .C(n27168), .Y(result[86]) );
  NOR2X1 U21925 ( .A(n27169), .B(n27170), .Y(n27168) );
  OR2X1 U21926 ( .A(n27171), .B(n27172), .Y(n27170) );
  OAI21X1 U21927 ( .A(n27173), .B(n25874), .C(n27174), .Y(n27172) );
  AOI22X1 U21928 ( .A(n27175), .B(n26014), .C(n27118), .D(n26125), .Y(n27174)
         );
  AND2X1 U21929 ( .A(n27176), .B(n27177), .Y(n27118) );
  AOI22X1 U21930 ( .A(n25838), .B(n26653), .C(n26160), .D(n26654), .Y(n27177)
         );
  INVX1 U21931 ( .A(n26409), .Y(n26653) );
  NOR2X1 U21932 ( .A(n27178), .B(n27179), .Y(n26409) );
  OAI22X1 U21933 ( .A(reg_A[78]), .B(n26131), .C(reg_A[86]), .D(n25894), .Y(
        n27179) );
  OAI21X1 U21934 ( .A(reg_A[70]), .B(n27027), .C(n27028), .Y(n27178) );
  AOI22X1 U21935 ( .A(n26159), .B(n27180), .C(n26059), .D(n27029), .Y(n27176)
         );
  INVX1 U21936 ( .A(n27181), .Y(n27029) );
  OAI21X1 U21937 ( .A(n27134), .B(n25914), .C(n27182), .Y(n27171) );
  AOI22X1 U21938 ( .A(n27183), .B(reg_A[84]), .C(reg_A[86]), .D(n27184), .Y(
        n27182) );
  NAND3X1 U21939 ( .A(n27185), .B(n27186), .C(n27187), .Y(n27169) );
  AOI21X1 U21940 ( .A(n27188), .B(reg_A[85]), .C(n27189), .Y(n27187) );
  OAI21X1 U21941 ( .A(n26141), .B(n27190), .C(n27191), .Y(n27189) );
  OAI21X1 U21942 ( .A(n27192), .B(n27193), .C(reg_A[80]), .Y(n27191) );
  OAI21X1 U21943 ( .A(n25032), .B(n26112), .C(n27194), .Y(n27193) );
  NAND2X1 U21944 ( .A(n27195), .B(n27196), .Y(n26141) );
  AOI22X1 U21945 ( .A(n26601), .B(n26230), .C(n26602), .D(n25875), .Y(n27196)
         );
  AOI22X1 U21946 ( .A(n27012), .B(n26039), .C(n26597), .D(n26215), .Y(n27195)
         );
  AOI22X1 U21947 ( .A(n27197), .B(n27155), .C(n27198), .D(n26504), .Y(n27186)
         );
  MUX2X1 U21948 ( .B(n27199), .A(n27200), .S(reg_B[87]), .Y(n27198) );
  INVX1 U21949 ( .A(n27201), .Y(n27200) );
  INVX1 U21950 ( .A(n27202), .Y(n27197) );
  AOI22X1 U21951 ( .A(n27203), .B(reg_B[95]), .C(n26886), .D(n25984), .Y(
        n27202) );
  OAI22X1 U21952 ( .A(n26067), .B(n26039), .C(n25874), .D(n26069), .Y(n26886)
         );
  AOI22X1 U21953 ( .A(n27204), .B(reg_A[83]), .C(n27205), .D(n27206), .Y(
        n27185) );
  NOR2X1 U21954 ( .A(n27207), .B(n27208), .Y(n27167) );
  OAI21X1 U21955 ( .A(n27209), .B(n27152), .C(n27210), .Y(n27208) );
  AOI22X1 U21956 ( .A(n27211), .B(n26260), .C(n26045), .D(n27212), .Y(n27210)
         );
  NAND3X1 U21957 ( .A(n27213), .B(n27214), .C(n27215), .Y(n27212) );
  NOR2X1 U21958 ( .A(n27216), .B(n27217), .Y(n27215) );
  OAI22X1 U21959 ( .A(n27218), .B(n26215), .C(n25207), .D(n26094), .Y(n27217)
         );
  OAI21X1 U21960 ( .A(n27219), .B(n25584), .C(n27220), .Y(n27216) );
  OAI21X1 U21961 ( .A(n27221), .B(n27222), .C(n25044), .Y(n27220) );
  NAND3X1 U21962 ( .A(n27223), .B(n27224), .C(n27225), .Y(n27222) );
  NOR2X1 U21963 ( .A(n27226), .B(n27227), .Y(n27225) );
  OAI21X1 U21964 ( .A(n25036), .B(n25863), .C(n27228), .Y(n27227) );
  AOI22X1 U21965 ( .A(reg_A[78]), .B(n25124), .C(reg_A[75]), .D(n25222), .Y(
        n27228) );
  OAI21X1 U21966 ( .A(n25037), .B(n26286), .C(n27229), .Y(n27226) );
  AOI22X1 U21967 ( .A(reg_A[82]), .B(n25070), .C(reg_A[81]), .D(n25123), .Y(
        n27229) );
  AOI21X1 U21968 ( .A(reg_A[74]), .B(n25635), .C(n27230), .Y(n27224) );
  OAI22X1 U21969 ( .A(n25065), .B(n26101), .C(n25035), .D(n26547), .Y(n27230)
         );
  AOI22X1 U21970 ( .A(reg_A[73]), .B(n25325), .C(reg_A[86]), .D(n25125), .Y(
        n27223) );
  NAND2X1 U21971 ( .A(n27231), .B(n27232), .Y(n27221) );
  NOR2X1 U21972 ( .A(n27233), .B(n27234), .Y(n27232) );
  OAI21X1 U21973 ( .A(n25238), .B(n25884), .C(n27235), .Y(n27234) );
  AOI22X1 U21974 ( .A(reg_A[68]), .B(n25241), .C(reg_A[64]), .D(n25242), .Y(
        n27235) );
  OAI21X1 U21975 ( .A(n25038), .B(n25851), .C(n27236), .Y(n27233) );
  AOI22X1 U21976 ( .A(reg_A[69]), .B(n25246), .C(reg_A[70]), .D(n25247), .Y(
        n27236) );
  NOR2X1 U21977 ( .A(n27237), .B(n27238), .Y(n27231) );
  OAI21X1 U21978 ( .A(n25030), .B(n25864), .C(n27239), .Y(n27238) );
  AOI22X1 U21979 ( .A(reg_A[84]), .B(n25252), .C(reg_A[80]), .D(n25253), .Y(
        n27239) );
  OAI21X1 U21980 ( .A(n25041), .B(n25875), .C(n27240), .Y(n27237) );
  AOI22X1 U21981 ( .A(reg_A[65]), .B(n25257), .C(reg_A[85]), .D(n25135), .Y(
        n27240) );
  AOI22X1 U21982 ( .A(reg_A[83]), .B(n27241), .C(reg_A[82]), .D(n27242), .Y(
        n27214) );
  AOI22X1 U21983 ( .A(reg_A[84]), .B(n27243), .C(reg_A[86]), .D(n25434), .Y(
        n27213) );
  INVX1 U21984 ( .A(n27244), .Y(n27211) );
  AND2X1 U21985 ( .A(n27245), .B(n27246), .Y(n27209) );
  NOR2X1 U21986 ( .A(n27247), .B(n27248), .Y(n27246) );
  OAI22X1 U21987 ( .A(n26936), .B(n25881), .C(n25745), .D(n25882), .Y(n27248)
         );
  OAI21X1 U21988 ( .A(n25062), .B(n26195), .C(n27249), .Y(n27247) );
  AOI22X1 U21989 ( .A(reg_A[87]), .B(n26803), .C(reg_A[89]), .D(n26804), .Y(
        n27249) );
  NOR2X1 U21990 ( .A(n27250), .B(n27251), .Y(n27245) );
  OAI22X1 U21991 ( .A(n25736), .B(n26039), .C(n27252), .D(n25883), .Y(n27251)
         );
  OAI21X1 U21992 ( .A(n27253), .B(n25873), .C(n27254), .Y(n27250) );
  AOI22X1 U21993 ( .A(reg_A[90]), .B(n25749), .C(reg_A[91]), .D(n25750), .Y(
        n27254) );
  OAI21X1 U21994 ( .A(n26525), .B(n27158), .C(n27255), .Y(n27207) );
  AOI22X1 U21995 ( .A(n26050), .B(n27062), .C(reg_A[81]), .D(n27256), .Y(
        n27255) );
  NAND2X1 U21996 ( .A(n27257), .B(n27258), .Y(n27062) );
  AOI22X1 U21997 ( .A(n25838), .B(n26339), .C(n26160), .D(n26611), .Y(n27258)
         );
  OAI21X1 U21998 ( .A(n26131), .B(n25865), .C(n27259), .Y(n26339) );
  AOI22X1 U21999 ( .A(reg_A[70]), .B(n26513), .C(reg_A[86]), .D(n26134), .Y(
        n27259) );
  AOI22X1 U22000 ( .A(n26059), .B(n26975), .C(n26159), .D(n27260), .Y(n27257)
         );
  NAND2X1 U22001 ( .A(n27261), .B(n27262), .Y(n27158) );
  AOI22X1 U22002 ( .A(n25025), .B(n26978), .C(n25026), .D(n26659), .Y(n27262)
         );
  INVX1 U22003 ( .A(n27263), .Y(n26978) );
  AOI22X1 U22004 ( .A(n26032), .B(n26658), .C(n26530), .D(n27264), .Y(n27261)
         );
  INVX1 U22005 ( .A(n26361), .Y(n26658) );
  NOR2X1 U22006 ( .A(n27265), .B(n27266), .Y(n26361) );
  OAI22X1 U22007 ( .A(reg_A[86]), .B(n25063), .C(reg_A[78]), .D(n26981), .Y(
        n27266) );
  OAI21X1 U22008 ( .A(reg_A[70]), .B(n26982), .C(n26983), .Y(n27265) );
  NOR2X1 U22009 ( .A(n27267), .B(n27268), .Y(n27166) );
  OAI21X1 U22010 ( .A(n25719), .B(n25965), .C(n27269), .Y(n27268) );
  AOI22X1 U22011 ( .A(n27141), .B(n27201), .C(n27270), .D(n27149), .Y(n27269)
         );
  OAI21X1 U22012 ( .A(n27271), .B(n27020), .C(n27272), .Y(n27267) );
  AOI22X1 U22013 ( .A(n25310), .B(n27273), .C(n27274), .D(n27142), .Y(n27272)
         );
  OAI21X1 U22014 ( .A(n27275), .B(n27276), .C(n27199), .Y(n27142) );
  AOI21X1 U22015 ( .A(reg_A[84]), .B(n27277), .C(n27105), .Y(n27199) );
  OAI22X1 U22016 ( .A(n26039), .B(n27278), .C(n25874), .D(n27279), .Y(n27105)
         );
  NAND2X1 U22017 ( .A(reg_B[85]), .B(reg_A[80]), .Y(n27276) );
  NAND3X1 U22018 ( .A(n27280), .B(n27281), .C(n27282), .Y(n27273) );
  NOR2X1 U22019 ( .A(n27283), .B(n27284), .Y(n27282) );
  OAI22X1 U22020 ( .A(n25043), .B(n26039), .C(n25467), .D(n25883), .Y(n27284)
         );
  OAI21X1 U22021 ( .A(n25037), .B(n25873), .C(n27285), .Y(n27283) );
  AOI22X1 U22022 ( .A(reg_A[90]), .B(n25070), .C(reg_A[91]), .D(n25123), .Y(
        n27285) );
  AOI21X1 U22023 ( .A(reg_A[88]), .B(n25252), .C(n27286), .Y(n27281) );
  OAI22X1 U22024 ( .A(n25041), .B(n25929), .C(n25784), .D(n25965), .Y(n27286)
         );
  AOI22X1 U22025 ( .A(reg_A[92]), .B(n25253), .C(reg_A[93]), .D(n25628), .Y(
        n27280) );
  NAND3X1 U22026 ( .A(n27287), .B(n27288), .C(n27289), .Y(result[85]) );
  NOR2X1 U22027 ( .A(n27290), .B(n27291), .Y(n27289) );
  OR2X1 U22028 ( .A(n27292), .B(n27293), .Y(n27291) );
  OAI21X1 U22029 ( .A(n27294), .B(n26215), .C(n27295), .Y(n27293) );
  AOI22X1 U22030 ( .A(n27296), .B(n26014), .C(n27175), .D(n26125), .Y(n27295)
         );
  INVX1 U22031 ( .A(n27297), .Y(n27175) );
  OAI21X1 U22032 ( .A(n27123), .B(n25898), .C(n27298), .Y(n27297) );
  AOI22X1 U22033 ( .A(n25838), .B(n27299), .C(reg_B[94]), .D(n27300), .Y(
        n27298) );
  INVX1 U22034 ( .A(n26514), .Y(n27299) );
  NOR2X1 U22035 ( .A(n27301), .B(n27302), .Y(n26514) );
  OAI22X1 U22036 ( .A(reg_A[77]), .B(n26131), .C(reg_A[85]), .D(n25894), .Y(
        n27302) );
  OAI21X1 U22037 ( .A(reg_A[69]), .B(n27027), .C(n27028), .Y(n27301) );
  INVX1 U22038 ( .A(n27303), .Y(n27294) );
  OAI21X1 U22039 ( .A(n27134), .B(n26168), .C(n27304), .Y(n27292) );
  AOI22X1 U22040 ( .A(reg_A[80]), .B(n27305), .C(n25310), .D(n27306), .Y(
        n27304) );
  NAND3X1 U22041 ( .A(n27307), .B(n27308), .C(n27309), .Y(n27306) );
  NOR2X1 U22042 ( .A(n27310), .B(n27311), .Y(n27309) );
  OAI22X1 U22043 ( .A(n25036), .B(n25873), .C(n25467), .D(n25881), .Y(n27311)
         );
  OAI21X1 U22044 ( .A(n25037), .B(n25883), .C(n27312), .Y(n27310) );
  AOI22X1 U22045 ( .A(reg_A[89]), .B(n25071), .C(reg_A[90]), .D(n25123), .Y(
        n27312) );
  AOI21X1 U22046 ( .A(reg_A[87]), .B(n25252), .C(n27313), .Y(n27308) );
  OAI22X1 U22047 ( .A(n25041), .B(n26195), .C(n25042), .D(n26039), .Y(n27313)
         );
  AOI22X1 U22048 ( .A(reg_A[91]), .B(n25253), .C(reg_A[92]), .D(n25628), .Y(
        n27307) );
  NAND3X1 U22049 ( .A(n27194), .B(n27314), .C(n27315), .Y(n27305) );
  INVX1 U22050 ( .A(n27316), .Y(n27315) );
  NAND3X1 U22051 ( .A(n25188), .B(n25972), .C(reg_B[93]), .Y(n27314) );
  AOI21X1 U22052 ( .A(reg_B[86]), .B(n27317), .C(n25890), .Y(n27194) );
  NOR2X1 U22053 ( .A(n26063), .B(n25032), .Y(n25890) );
  NOR2X1 U22054 ( .A(n27318), .B(n25031), .Y(n27317) );
  AOI22X1 U22055 ( .A(n27319), .B(n26267), .C(reg_A[84]), .D(n26396), .Y(
        n27134) );
  NOR2X1 U22056 ( .A(n26067), .B(n25032), .Y(n26396) );
  NAND3X1 U22057 ( .A(n27320), .B(n27321), .C(n27322), .Y(n27290) );
  AOI21X1 U22058 ( .A(n27323), .B(reg_A[81]), .C(n27324), .Y(n27322) );
  OAI22X1 U22059 ( .A(n27325), .B(n27326), .C(n27327), .D(n25342), .Y(n27324)
         );
  AOI22X1 U22060 ( .A(n27277), .B(n27328), .C(n27106), .D(n27275), .Y(n27327)
         );
  MUX2X1 U22061 ( .B(n27329), .A(n27330), .S(reg_B[87]), .Y(n27106) );
  MUX2X1 U22062 ( .B(reg_A[84]), .A(reg_A[80]), .S(reg_B[85]), .Y(n27330) );
  MUX2X1 U22063 ( .B(reg_A[85]), .A(reg_A[81]), .S(reg_B[85]), .Y(n27329) );
  OAI21X1 U22064 ( .A(n25874), .B(n27057), .C(n27331), .Y(n27328) );
  INVX1 U22065 ( .A(n27206), .Y(n27326) );
  OAI21X1 U22066 ( .A(n27332), .B(n27333), .C(n25840), .Y(n27321) );
  NAND3X1 U22067 ( .A(n27334), .B(n27335), .C(n27336), .Y(n27333) );
  NOR2X1 U22068 ( .A(n27337), .B(n27338), .Y(n27336) );
  OAI21X1 U22069 ( .A(n25036), .B(n26103), .C(n27339), .Y(n27338) );
  AOI22X1 U22070 ( .A(reg_A[77]), .B(n25124), .C(reg_A[74]), .D(n25222), .Y(
        n27339) );
  OAI21X1 U22071 ( .A(n25037), .B(n25863), .C(n27340), .Y(n27337) );
  AOI22X1 U22072 ( .A(reg_A[81]), .B(n25071), .C(reg_A[80]), .D(n25123), .Y(
        n27340) );
  AOI21X1 U22073 ( .A(reg_A[73]), .B(n25635), .C(n27341), .Y(n27335) );
  OAI22X1 U22074 ( .A(n25065), .B(n26256), .C(n25035), .D(n26101), .Y(n27341)
         );
  AOI22X1 U22075 ( .A(reg_A[72]), .B(n25325), .C(reg_A[85]), .D(n25125), .Y(
        n27334) );
  NAND3X1 U22076 ( .A(n27342), .B(n27343), .C(n27344), .Y(n27332) );
  NOR2X1 U22077 ( .A(n27345), .B(n27346), .Y(n27344) );
  OAI21X1 U22078 ( .A(n26719), .B(n25853), .C(n27347), .Y(n27346) );
  AOI22X1 U22079 ( .A(reg_A[67]), .B(n25241), .C(reg_A[65]), .D(n25339), .Y(
        n27347) );
  OAI21X1 U22080 ( .A(n25038), .B(n25884), .C(n27348), .Y(n27345) );
  AOI22X1 U22081 ( .A(reg_A[68]), .B(n25246), .C(reg_A[69]), .D(n25247), .Y(
        n27348) );
  AOI21X1 U22082 ( .A(reg_A[83]), .B(n25252), .C(n27349), .Y(n27343) );
  OAI22X1 U22083 ( .A(n25041), .B(n25874), .C(n25042), .D(n26230), .Y(n27349)
         );
  AOI22X1 U22084 ( .A(reg_A[79]), .B(n25253), .C(reg_A[78]), .D(n25628), .Y(
        n27342) );
  AOI22X1 U22085 ( .A(n27350), .B(n27351), .C(n27352), .D(n27203), .Y(n27320)
         );
  OAI22X1 U22086 ( .A(reg_B[94]), .B(n26994), .C(n25875), .D(n26872), .Y(
        n27203) );
  AOI22X1 U22087 ( .A(n26275), .B(reg_A[85]), .C(reg_A[81]), .D(n26274), .Y(
        n26994) );
  OAI21X1 U22088 ( .A(reg_B[95]), .B(n25794), .C(n27353), .Y(n27352) );
  NOR2X1 U22089 ( .A(n27354), .B(n26169), .Y(n27350) );
  NOR2X1 U22090 ( .A(n27355), .B(n27356), .Y(n27288) );
  OAI21X1 U22091 ( .A(n27271), .B(n26950), .C(n27357), .Y(n27356) );
  AOI22X1 U22092 ( .A(n27358), .B(n27359), .C(n25730), .D(n27360), .Y(n27357)
         );
  NAND3X1 U22093 ( .A(n27361), .B(n27362), .C(n27363), .Y(n27360) );
  NOR2X1 U22094 ( .A(n27364), .B(n27365), .Y(n27363) );
  OAI21X1 U22095 ( .A(n26801), .B(n25929), .C(n27366), .Y(n27365) );
  AOI22X1 U22096 ( .A(reg_A[91]), .B(n26878), .C(reg_A[92]), .D(n25613), .Y(
        n27366) );
  OAI21X1 U22097 ( .A(n25062), .B(n25965), .C(n27367), .Y(n27364) );
  AOI22X1 U22098 ( .A(reg_A[86]), .B(n26803), .C(reg_A[88]), .D(n26804), .Y(
        n27367) );
  AOI21X1 U22099 ( .A(reg_A[93]), .B(n25615), .C(n27368), .Y(n27362) );
  OAI22X1 U22100 ( .A(n27253), .B(n25883), .C(n26800), .D(n26068), .Y(n27368)
         );
  AOI22X1 U22101 ( .A(reg_A[95]), .B(n25607), .C(reg_A[85]), .D(n26924), .Y(
        n27361) );
  NAND3X1 U22102 ( .A(n27369), .B(n27370), .C(n27371), .Y(n27359) );
  NOR2X1 U22103 ( .A(n27372), .B(n27373), .Y(n27371) );
  OAI22X1 U22104 ( .A(n27130), .B(n27374), .C(n25584), .D(n27375), .Y(n27373)
         );
  NAND2X1 U22105 ( .A(n27376), .B(n26317), .Y(n27130) );
  AOI22X1 U22106 ( .A(n26230), .B(n26295), .C(n26215), .D(n26293), .Y(n26317)
         );
  AOI22X1 U22107 ( .A(n26292), .B(n26094), .C(n26294), .D(n25584), .Y(n27376)
         );
  OAI22X1 U22108 ( .A(n27244), .B(n27377), .C(n27378), .D(n27379), .Y(n27372)
         );
  OAI21X1 U22109 ( .A(n27380), .B(n26030), .C(n27381), .Y(n27244) );
  AOI22X1 U22110 ( .A(n25025), .B(n27127), .C(n26032), .D(n26531), .Y(n27381)
         );
  OR2X1 U22111 ( .A(n27382), .B(n27383), .Y(n26531) );
  OAI22X1 U22112 ( .A(reg_A[85]), .B(n26036), .C(reg_A[77]), .D(n26981), .Y(
        n27383) );
  OAI21X1 U22113 ( .A(reg_A[69]), .B(n26982), .C(n26983), .Y(n27382) );
  INVX1 U22114 ( .A(n27384), .Y(n27127) );
  INVX1 U22115 ( .A(n27385), .Y(n27380) );
  AOI22X1 U22116 ( .A(reg_A[82]), .B(n27386), .C(reg_A[81]), .D(n27387), .Y(
        n27370) );
  AOI22X1 U22117 ( .A(reg_A[83]), .B(n27388), .C(n27389), .D(reg_A[85]), .Y(
        n27369) );
  AND2X1 U22118 ( .A(n27390), .B(n27391), .Y(n27271) );
  AOI22X1 U22119 ( .A(n25838), .B(n26510), .C(n26160), .D(n26906), .Y(n27391)
         );
  OAI21X1 U22120 ( .A(n26131), .B(n26286), .C(n27392), .Y(n26510) );
  AOI22X1 U22121 ( .A(n26513), .B(reg_A[69]), .C(reg_A[85]), .D(n26134), .Y(
        n27392) );
  AOI22X1 U22122 ( .A(n26059), .B(n27114), .C(n26159), .D(n27393), .Y(n27390)
         );
  OAI21X1 U22123 ( .A(n27394), .B(n26230), .C(n27395), .Y(n27355) );
  AOI22X1 U22124 ( .A(reg_A[82]), .B(n27396), .C(reg_A[83]), .D(n27397), .Y(
        n27395) );
  NOR2X1 U22125 ( .A(n27398), .B(n27399), .Y(n27287) );
  OAI21X1 U22126 ( .A(n25717), .B(n25965), .C(n27400), .Y(n27399) );
  AOI22X1 U22127 ( .A(n27401), .B(n27149), .C(reg_A[86]), .D(n27402), .Y(
        n27400) );
  OAI21X1 U22128 ( .A(n27403), .B(n27404), .C(n27405), .Y(n27398) );
  AOI22X1 U22129 ( .A(n27274), .B(n27201), .C(n26116), .D(n27406), .Y(n27405)
         );
  OAI21X1 U22130 ( .A(n26215), .B(n27278), .C(n27407), .Y(n27201) );
  AOI22X1 U22131 ( .A(n27101), .B(reg_A[81]), .C(n27277), .D(reg_A[83]), .Y(
        n27407) );
  INVX1 U22132 ( .A(n27408), .Y(n27403) );
  NAND2X1 U22133 ( .A(n27409), .B(n27410), .Y(result[84]) );
  NOR2X1 U22134 ( .A(n27411), .B(n27412), .Y(n27410) );
  NAND3X1 U22135 ( .A(n27413), .B(n27414), .C(n27415), .Y(n27412) );
  NOR2X1 U22136 ( .A(n27416), .B(n27417), .Y(n27415) );
  OAI22X1 U22137 ( .A(n27418), .B(n25874), .C(n27419), .D(n26094), .Y(n27417)
         );
  OAI22X1 U22138 ( .A(n25360), .B(n25965), .C(n27420), .D(n26039), .Y(n27416)
         );
  AOI22X1 U22139 ( .A(reg_A[84]), .B(n27421), .C(n27206), .D(n27422), .Y(
        n27414) );
  NOR2X1 U22140 ( .A(n25523), .B(reg_B[85]), .Y(n27206) );
  OAI21X1 U22141 ( .A(n25032), .B(n26377), .C(n27423), .Y(n27421) );
  AOI22X1 U22142 ( .A(reg_A[80]), .B(n27424), .C(n27296), .D(n26125), .Y(
        n27413) );
  AOI21X1 U22143 ( .A(n27425), .B(reg_B[94]), .C(n27426), .Y(n27296) );
  INVX1 U22144 ( .A(n27427), .Y(n27426) );
  AOI22X1 U22145 ( .A(n25838), .B(n26654), .C(n26059), .D(n27180), .Y(n27427)
         );
  OR2X1 U22146 ( .A(n27428), .B(n27429), .Y(n26654) );
  OAI22X1 U22147 ( .A(reg_A[76]), .B(n26131), .C(reg_A[84]), .D(n25894), .Y(
        n27429) );
  OAI21X1 U22148 ( .A(reg_A[68]), .B(n27027), .C(n27028), .Y(n27428) );
  OAI21X1 U22149 ( .A(n26275), .B(n25794), .C(n27430), .Y(n27424) );
  AOI21X1 U22150 ( .A(reg_B[85]), .B(n26504), .C(n27323), .Y(n27430) );
  INVX1 U22151 ( .A(n27431), .Y(n27323) );
  NAND3X1 U22152 ( .A(n27432), .B(n27433), .C(n27434), .Y(n27411) );
  NOR2X1 U22153 ( .A(n27435), .B(n27436), .Y(n27434) );
  OAI21X1 U22154 ( .A(n27437), .B(n27438), .C(n27439), .Y(n27436) );
  OAI21X1 U22155 ( .A(n27440), .B(n27441), .C(n27358), .Y(n27439) );
  OAI22X1 U22156 ( .A(n26230), .B(n27442), .C(n27443), .D(n27444), .Y(n27441)
         );
  OAI21X1 U22157 ( .A(n27445), .B(n25403), .C(n27446), .Y(n27440) );
  INVX1 U22158 ( .A(n27447), .Y(n27446) );
  OAI22X1 U22159 ( .A(n27448), .B(n25584), .C(n27449), .D(n26422), .Y(n27447)
         );
  NAND2X1 U22160 ( .A(n27450), .B(n27451), .Y(n26422) );
  AOI22X1 U22161 ( .A(n26601), .B(n25874), .C(n26602), .D(n26094), .Y(n27451)
         );
  AOI22X1 U22162 ( .A(n27012), .B(n26230), .C(n26597), .D(n25875), .Y(n27450)
         );
  AOI21X1 U22163 ( .A(n27452), .B(n26863), .C(n27453), .Y(n27445) );
  OAI22X1 U22164 ( .A(n27454), .B(n27385), .C(n27455), .D(n27456), .Y(n27453)
         );
  INVX1 U22165 ( .A(n27378), .Y(n27452) );
  OAI21X1 U22166 ( .A(n27457), .B(n26030), .C(n27458), .Y(n27378) );
  AOI22X1 U22167 ( .A(n25025), .B(n27264), .C(n26032), .D(n26659), .Y(n27458)
         );
  OR2X1 U22168 ( .A(n27459), .B(n27460), .Y(n26659) );
  OAI22X1 U22169 ( .A(reg_A[84]), .B(n26036), .C(reg_A[76]), .D(n26981), .Y(
        n27460) );
  OAI21X1 U22170 ( .A(reg_A[68]), .B(n26982), .C(n26983), .Y(n27459) );
  INVX1 U22171 ( .A(n27461), .Y(n27437) );
  OAI22X1 U22172 ( .A(n27300), .B(n26168), .C(n27462), .D(n26169), .Y(n27461)
         );
  OAI21X1 U22173 ( .A(n27353), .B(n27463), .C(n27464), .Y(n27435) );
  OAI21X1 U22174 ( .A(n27465), .B(n27466), .C(n25840), .Y(n27464) );
  NAND3X1 U22175 ( .A(n27467), .B(n27468), .C(n27469), .Y(n27466) );
  NOR2X1 U22176 ( .A(n27470), .B(n27471), .Y(n27469) );
  OAI22X1 U22177 ( .A(n25043), .B(n26230), .C(n25039), .D(n26101), .Y(n27471)
         );
  OAI21X1 U22178 ( .A(n25064), .B(n26547), .C(n27472), .Y(n27470) );
  AOI22X1 U22179 ( .A(reg_A[70]), .B(n25234), .C(reg_A[69]), .D(n25235), .Y(
        n27472) );
  AOI21X1 U22180 ( .A(reg_A[76]), .B(n25124), .C(n27473), .Y(n27468) );
  OAI22X1 U22181 ( .A(n25037), .B(n26103), .C(n26703), .D(n25864), .Y(n27473)
         );
  AOI22X1 U22182 ( .A(reg_A[73]), .B(n25222), .C(reg_A[74]), .D(n25637), .Y(
        n27467) );
  NAND3X1 U22183 ( .A(n27474), .B(n27475), .C(n27476), .Y(n27465) );
  NOR2X1 U22184 ( .A(n27477), .B(n27478), .Y(n27476) );
  OAI21X1 U22185 ( .A(n25042), .B(n25875), .C(n27479), .Y(n27478) );
  AOI22X1 U22186 ( .A(reg_A[66]), .B(n25241), .C(reg_A[64]), .D(n25339), .Y(
        n27479) );
  OAI21X1 U22187 ( .A(n25038), .B(n25855), .C(n27480), .Y(n27477) );
  AOI22X1 U22188 ( .A(reg_A[67]), .B(n25246), .C(reg_A[68]), .D(n25247), .Y(
        n27480) );
  AOI21X1 U22189 ( .A(reg_A[78]), .B(n25253), .C(n27481), .Y(n27475) );
  OAI22X1 U22190 ( .A(n25040), .B(n25874), .C(n25041), .D(n26094), .Y(n27481)
         );
  AOI22X1 U22191 ( .A(reg_A[77]), .B(n25628), .C(reg_A[80]), .D(n25067), .Y(
        n27474) );
  MUX2X1 U22192 ( .B(n27319), .A(n27351), .S(reg_B[94]), .Y(n27463) );
  OAI22X1 U22193 ( .A(n26067), .B(n26230), .C(n25584), .D(n26069), .Y(n27319)
         );
  AOI22X1 U22194 ( .A(n27482), .B(n27483), .C(n27484), .D(n27485), .Y(n27433)
         );
  MUX2X1 U22195 ( .B(n25874), .A(n26094), .S(reg_B[87]), .Y(n27485) );
  NOR2X1 U22196 ( .A(n25517), .B(n27061), .Y(n27484) );
  MUX2X1 U22197 ( .B(n26230), .A(n25875), .S(reg_B[87]), .Y(n27483) );
  NOR2X1 U22198 ( .A(n25031), .B(n27278), .Y(n27482) );
  AOI22X1 U22199 ( .A(n27486), .B(reg_B[95]), .C(n27487), .D(n27351), .Y(
        n27432) );
  INVX1 U22200 ( .A(n27488), .Y(n27351) );
  NOR2X1 U22201 ( .A(n25032), .B(n25914), .Y(n27487) );
  NOR2X1 U22202 ( .A(n27354), .B(n27489), .Y(n27486) );
  NOR2X1 U22203 ( .A(n27490), .B(n27491), .Y(n27409) );
  NAND3X1 U22204 ( .A(n27492), .B(n27493), .C(n27494), .Y(n27491) );
  INVX1 U22205 ( .A(n27495), .Y(n27494) );
  OAI21X1 U22206 ( .A(n27404), .B(n27496), .C(n27497), .Y(n27495) );
  AOI22X1 U22207 ( .A(n27498), .B(n26116), .C(n27149), .D(n27499), .Y(n27497)
         );
  OAI21X1 U22208 ( .A(reg_B[91]), .B(n26996), .C(n27500), .Y(n27149) );
  AOI22X1 U22209 ( .A(reg_A[91]), .B(n25293), .C(reg_A[85]), .D(n25282), .Y(
        n27493) );
  AOI22X1 U22210 ( .A(n26050), .B(n27406), .C(n27274), .D(n27408), .Y(n27492)
         );
  OAI21X1 U22211 ( .A(n26230), .B(n27278), .C(n27501), .Y(n27408) );
  AOI22X1 U22212 ( .A(n27101), .B(reg_A[80]), .C(n27277), .D(reg_A[82]), .Y(
        n27501) );
  INVX1 U22213 ( .A(n27279), .Y(n27101) );
  NAND2X1 U22214 ( .A(reg_B[85]), .B(n27275), .Y(n27279) );
  NAND2X1 U22215 ( .A(n27502), .B(n27503), .Y(n27406) );
  AOI22X1 U22216 ( .A(n25838), .B(n26611), .C(n26160), .D(n26975), .Y(n27503)
         );
  OAI21X1 U22217 ( .A(n26131), .B(n25863), .C(n27504), .Y(n26611) );
  AOI22X1 U22218 ( .A(reg_A[68]), .B(n26513), .C(reg_A[84]), .D(n26134), .Y(
        n27504) );
  AOI22X1 U22219 ( .A(n26059), .B(n27260), .C(n26159), .D(n27505), .Y(n27502)
         );
  NAND3X1 U22220 ( .A(n27506), .B(n27507), .C(n27508), .Y(n27490) );
  NOR2X1 U22221 ( .A(n27509), .B(n27510), .Y(n27508) );
  OAI22X1 U22222 ( .A(n25295), .B(n26068), .C(n25297), .D(n25929), .Y(n27510)
         );
  OAI22X1 U22223 ( .A(n27511), .B(n26195), .C(n27512), .D(n25882), .Y(n27509)
         );
  AOI22X1 U22224 ( .A(reg_A[83]), .B(n27513), .C(reg_A[94]), .D(n25299), .Y(
        n27507) );
  AOI22X1 U22225 ( .A(reg_A[95]), .B(n25300), .C(reg_A[93]), .D(n25301), .Y(
        n27506) );
  NAND3X1 U22226 ( .A(n27514), .B(n27515), .C(n27516), .Y(result[83]) );
  NOR2X1 U22227 ( .A(n27517), .B(n27518), .Y(n27516) );
  NAND2X1 U22228 ( .A(n27519), .B(n27520), .Y(n27518) );
  AOI21X1 U22229 ( .A(n26050), .B(n27498), .C(n27521), .Y(n27520) );
  OAI21X1 U22230 ( .A(n27522), .B(n27523), .C(n27524), .Y(n27521) );
  OAI21X1 U22231 ( .A(n27525), .B(n27526), .C(n25372), .Y(n27524) );
  NAND3X1 U22232 ( .A(n27527), .B(n27528), .C(n27529), .Y(n27526) );
  MUX2X1 U22233 ( .B(n27530), .A(n27531), .S(reg_B[87]), .Y(n27529) );
  INVX1 U22234 ( .A(n27532), .Y(n27531) );
  NOR2X1 U22235 ( .A(n27496), .B(n26999), .Y(n27530) );
  MUX2X1 U22236 ( .B(n27533), .A(n27534), .S(reg_B[94]), .Y(n27527) );
  OAI21X1 U22237 ( .A(n26896), .B(n27462), .C(n27535), .Y(n27534) );
  OAI21X1 U22238 ( .A(n27536), .B(n27537), .C(n25980), .Y(n27535) );
  AND2X1 U22239 ( .A(n25895), .B(n27538), .Y(n27536) );
  OAI22X1 U22240 ( .A(n27053), .B(n27425), .C(n26896), .D(n27300), .Y(n27533)
         );
  OAI21X1 U22241 ( .A(reg_B[93]), .B(n26843), .C(n27539), .Y(n27300) );
  AOI21X1 U22242 ( .A(n27540), .B(n25896), .C(n27541), .Y(n27539) );
  NOR2X1 U22243 ( .A(n27542), .B(n27543), .Y(n26843) );
  OAI22X1 U22244 ( .A(reg_A[75]), .B(n26131), .C(reg_A[83]), .D(n25894), .Y(
        n27543) );
  OAI21X1 U22245 ( .A(reg_A[67]), .B(n27027), .C(n27028), .Y(n27542) );
  OAI21X1 U22246 ( .A(n26169), .B(n27444), .C(n27544), .Y(n27525) );
  AOI22X1 U22247 ( .A(n27545), .B(n25604), .C(reg_A[82]), .D(n27546), .Y(
        n27544) );
  NOR2X1 U22248 ( .A(reg_B[95]), .B(n27489), .Y(n27545) );
  NAND2X1 U22249 ( .A(n27547), .B(n27548), .Y(n27498) );
  AOI22X1 U22250 ( .A(n25838), .B(n26906), .C(n26160), .D(n27114), .Y(n27548)
         );
  OAI21X1 U22251 ( .A(n26131), .B(n26103), .C(n27549), .Y(n26906) );
  AOI22X1 U22252 ( .A(reg_A[67]), .B(n26513), .C(reg_A[83]), .D(n26134), .Y(
        n27549) );
  AOI22X1 U22253 ( .A(n26059), .B(n27393), .C(n26159), .D(n27550), .Y(n27547)
         );
  AOI21X1 U22254 ( .A(n27141), .B(n27551), .C(n27552), .Y(n27519) );
  OAI22X1 U22255 ( .A(n27489), .B(n27353), .C(n27496), .D(n27553), .Y(n27552)
         );
  AOI22X1 U22256 ( .A(reg_A[83]), .B(n27104), .C(reg_A[81]), .D(n27277), .Y(
        n27496) );
  INVX1 U22257 ( .A(n27554), .Y(n27489) );
  OAI21X1 U22258 ( .A(n26094), .B(n26872), .C(n27555), .Y(n27554) );
  NAND3X1 U22259 ( .A(n26275), .B(n25950), .C(reg_A[83]), .Y(n27555) );
  INVX1 U22260 ( .A(n27404), .Y(n27141) );
  NAND3X1 U22261 ( .A(n27556), .B(n27557), .C(n27558), .Y(n27517) );
  AOI21X1 U22262 ( .A(reg_A[90]), .B(n25293), .C(n27559), .Y(n27558) );
  OAI22X1 U22263 ( .A(n25295), .B(n25929), .C(n25297), .D(n26195), .Y(n27559)
         );
  OAI21X1 U22264 ( .A(n27560), .B(n27561), .C(n27358), .Y(n27557) );
  OAI21X1 U22265 ( .A(n25438), .B(n25853), .C(n27522), .Y(n27561) );
  INVX1 U22266 ( .A(n27562), .Y(n27522) );
  OAI21X1 U22267 ( .A(n25204), .B(n25875), .C(n27563), .Y(n27562) );
  AOI22X1 U22268 ( .A(reg_A[82]), .B(n25441), .C(reg_A[81]), .D(n27243), .Y(
        n27563) );
  OAI21X1 U22269 ( .A(n27564), .B(n25584), .C(n27565), .Y(n27560) );
  OAI21X1 U22270 ( .A(n27566), .B(n27567), .C(n25044), .Y(n27565) );
  OAI22X1 U22271 ( .A(n27454), .B(n27568), .C(n26599), .D(n27385), .Y(n27567)
         );
  OAI21X1 U22272 ( .A(reg_B[2]), .B(n27126), .C(n27569), .Y(n27385) );
  AOI21X1 U22273 ( .A(n27570), .B(n27571), .C(n27572), .Y(n27569) );
  NOR2X1 U22274 ( .A(n27573), .B(n27574), .Y(n27126) );
  OAI22X1 U22275 ( .A(reg_A[83]), .B(n25063), .C(reg_A[75]), .D(n26981), .Y(
        n27574) );
  OAI21X1 U22276 ( .A(reg_A[67]), .B(n26982), .C(n26983), .Y(n27573) );
  OAI21X1 U22277 ( .A(n27575), .B(n27456), .C(n27576), .Y(n27566) );
  AOI22X1 U22278 ( .A(n27577), .B(n27578), .C(n27579), .D(reg_A[64]), .Y(
        n27576) );
  AOI22X1 U22279 ( .A(reg_A[84]), .B(n25282), .C(reg_A[83]), .D(n25283), .Y(
        n27556) );
  NOR2X1 U22280 ( .A(n27580), .B(n27581), .Y(n27515) );
  OAI21X1 U22281 ( .A(n27582), .B(n25873), .C(n27583), .Y(n27581) );
  AOI22X1 U22282 ( .A(reg_A[87]), .B(n25368), .C(n26116), .D(n27584), .Y(
        n27583) );
  OR2X1 U22283 ( .A(n27585), .B(n27586), .Y(n27580) );
  OAI21X1 U22284 ( .A(n25584), .B(n27587), .C(n27588), .Y(n27586) );
  OAI21X1 U22285 ( .A(n27589), .B(n27590), .C(n25382), .Y(n27588) );
  OAI22X1 U22286 ( .A(n27591), .B(n27592), .C(n27593), .D(n27058), .Y(n27590)
         );
  INVX1 U22287 ( .A(n27594), .Y(n27591) );
  OAI21X1 U22288 ( .A(n27595), .B(n27061), .C(n27596), .Y(n27589) );
  NAND3X1 U22289 ( .A(n27597), .B(n27275), .C(n27103), .Y(n27596) );
  OAI21X1 U22290 ( .A(n25976), .B(n27598), .C(n27599), .Y(n27585) );
  OAI21X1 U22291 ( .A(n27600), .B(n27601), .C(n25840), .Y(n27599) );
  NAND3X1 U22292 ( .A(n27602), .B(n27603), .C(n27604), .Y(n27601) );
  NOR2X1 U22293 ( .A(n27605), .B(n27606), .Y(n27604) );
  OAI22X1 U22294 ( .A(n25043), .B(n25875), .C(n25039), .D(n26256), .Y(n27606)
         );
  OAI21X1 U22295 ( .A(n25064), .B(n26101), .C(n27607), .Y(n27605) );
  AOI22X1 U22296 ( .A(reg_A[69]), .B(n25234), .C(reg_A[68]), .D(n25235), .Y(
        n27607) );
  AOI21X1 U22297 ( .A(reg_A[75]), .B(n25124), .C(n27608), .Y(n27603) );
  OAI22X1 U22298 ( .A(n25037), .B(n26438), .C(n26703), .D(n25865), .Y(n27608)
         );
  AOI22X1 U22299 ( .A(reg_A[72]), .B(n25222), .C(reg_A[73]), .D(n25637), .Y(
        n27602) );
  NAND3X1 U22300 ( .A(n27609), .B(n27610), .C(n27611), .Y(n27600) );
  NOR2X1 U22301 ( .A(n27612), .B(n27613), .Y(n27611) );
  OAI22X1 U22302 ( .A(n25042), .B(n25874), .C(n25331), .D(n25855), .Y(n27613)
         );
  OAI21X1 U22303 ( .A(n25038), .B(n25853), .C(n27614), .Y(n27612) );
  AOI22X1 U22304 ( .A(reg_A[66]), .B(n25246), .C(reg_A[67]), .D(n25247), .Y(
        n27614) );
  AOI21X1 U22305 ( .A(reg_A[77]), .B(n25253), .C(n27615), .Y(n27610) );
  OAI22X1 U22306 ( .A(n25040), .B(n26094), .C(n25041), .D(n25584), .Y(n27615)
         );
  AOI22X1 U22307 ( .A(reg_A[76]), .B(n25628), .C(reg_A[79]), .D(n25067), .Y(
        n27609) );
  NAND2X1 U22308 ( .A(n26267), .B(n27616), .Y(n27598) );
  NOR2X1 U22309 ( .A(n27617), .B(n27618), .Y(n27514) );
  OAI21X1 U22310 ( .A(n27512), .B(n25973), .C(n27619), .Y(n27618) );
  AOI22X1 U22311 ( .A(reg_A[94]), .B(n25300), .C(reg_A[92]), .D(n25301), .Y(
        n27619) );
  OAI21X1 U22312 ( .A(n27620), .B(n25881), .C(n27621), .Y(n27617) );
  AOI22X1 U22313 ( .A(reg_A[85]), .B(n25364), .C(reg_A[86]), .D(n27622), .Y(
        n27621) );
  OR2X1 U22314 ( .A(n27623), .B(n27624), .Y(result[82]) );
  NAND3X1 U22315 ( .A(n27625), .B(n27626), .C(n27627), .Y(n27624) );
  NOR2X1 U22316 ( .A(n27628), .B(n27629), .Y(n27627) );
  OAI21X1 U22317 ( .A(n27630), .B(n27020), .C(n27631), .Y(n27629) );
  OAI21X1 U22318 ( .A(n27632), .B(n27633), .C(n25203), .Y(n27631) );
  NAND3X1 U22319 ( .A(n27634), .B(n27635), .C(n27636), .Y(n27633) );
  AOI21X1 U22320 ( .A(reg_A[84]), .B(n27637), .C(n27638), .Y(n27636) );
  OAI22X1 U22321 ( .A(n25599), .B(n26215), .C(n25600), .D(n25965), .Y(n27638)
         );
  AOI22X1 U22322 ( .A(reg_A[82]), .B(n27639), .C(reg_A[83]), .D(n25617), .Y(
        n27635) );
  AOI22X1 U22323 ( .A(reg_A[86]), .B(n25650), .C(reg_A[88]), .D(n25651), .Y(
        n27634) );
  NAND3X1 U22324 ( .A(n27640), .B(n27641), .C(n27642), .Y(n27632) );
  AOI21X1 U22325 ( .A(reg_A[93]), .B(n27643), .C(n27644), .Y(n27642) );
  OAI22X1 U22326 ( .A(n27645), .B(n25882), .C(n27646), .D(n25973), .Y(n27644)
         );
  AOI22X1 U22327 ( .A(reg_A[94]), .B(n27647), .C(reg_A[95]), .D(n27648), .Y(
        n27641) );
  AOI22X1 U22328 ( .A(reg_A[89]), .B(n27649), .C(reg_A[90]), .D(n27650), .Y(
        n27640) );
  OAI21X1 U22329 ( .A(n27651), .B(n27652), .C(n27653), .Y(n27628) );
  OAI21X1 U22330 ( .A(n27654), .B(n27655), .C(n25372), .Y(n27653) );
  NAND2X1 U22331 ( .A(n27656), .B(n27528), .Y(n27655) );
  AOI22X1 U22332 ( .A(reg_A[81]), .B(n27546), .C(n26223), .D(reg_B[94]), .Y(
        n27656) );
  OAI21X1 U22333 ( .A(n25415), .B(n26381), .C(n27657), .Y(n27546) );
  OAI21X1 U22334 ( .A(n27658), .B(n25403), .C(n27659), .Y(n27654) );
  INVX1 U22335 ( .A(n27660), .Y(n27659) );
  OAI21X1 U22336 ( .A(n25874), .B(n27661), .C(n27532), .Y(n27660) );
  NAND3X1 U22337 ( .A(reg_A[80]), .B(n25589), .C(reg_B[86]), .Y(n27532) );
  NOR2X1 U22338 ( .A(n27662), .B(n27663), .Y(n27658) );
  OAI21X1 U22339 ( .A(n26169), .B(n27664), .C(n27665), .Y(n27663) );
  MUX2X1 U22340 ( .B(n27666), .A(n27667), .S(reg_B[93]), .Y(n27665) );
  OAI21X1 U22341 ( .A(reg_B[91]), .B(n27668), .C(n27664), .Y(n27667) );
  AOI22X1 U22342 ( .A(n26518), .B(n26149), .C(n26415), .D(n26276), .Y(n27668)
         );
  OAI21X1 U22343 ( .A(n25914), .B(n27180), .C(n27669), .Y(n27666) );
  NAND3X1 U22344 ( .A(n27670), .B(n25895), .C(n26149), .Y(n27669) );
  OAI21X1 U22345 ( .A(reg_A[64]), .B(n25895), .C(n27671), .Y(n27180) );
  AOI22X1 U22346 ( .A(n26134), .B(n25584), .C(n25892), .D(n26547), .Y(n27671)
         );
  OAI22X1 U22347 ( .A(n26168), .B(n27462), .C(n25972), .D(n27425), .Y(n27662)
         );
  OAI21X1 U22348 ( .A(reg_B[93]), .B(n27181), .C(n27672), .Y(n27425) );
  AOI21X1 U22349 ( .A(n27540), .B(n26133), .C(n27541), .Y(n27672) );
  NOR2X1 U22350 ( .A(n27673), .B(n27674), .Y(n27181) );
  OAI22X1 U22351 ( .A(reg_A[74]), .B(n26131), .C(reg_A[82]), .D(n25894), .Y(
        n27674) );
  OAI21X1 U22352 ( .A(reg_A[66]), .B(n27027), .C(n27028), .Y(n27673) );
  NAND2X1 U22353 ( .A(n27675), .B(n27676), .Y(n27652) );
  AOI22X1 U22354 ( .A(n26597), .B(n27456), .C(n26009), .D(n27264), .Y(n27675)
         );
  OAI21X1 U22355 ( .A(reg_A[64]), .B(n27677), .C(n27678), .Y(n27264) );
  AOI22X1 U22356 ( .A(n26038), .B(n26547), .C(n26664), .D(n25584), .Y(n27678)
         );
  OAI21X1 U22357 ( .A(n27457), .B(n26599), .C(n27679), .Y(n27651) );
  AOI22X1 U22358 ( .A(n27680), .B(n25853), .C(n27681), .D(n27677), .Y(n27679)
         );
  OAI21X1 U22359 ( .A(n27682), .B(n25754), .C(n27683), .Y(n27681) );
  AOI22X1 U22360 ( .A(n26002), .B(n26533), .C(n26008), .D(n27571), .Y(n27683)
         );
  INVX1 U22361 ( .A(n27568), .Y(n27457) );
  OAI21X1 U22362 ( .A(reg_B[2]), .B(n27263), .C(n27684), .Y(n27568) );
  AOI21X1 U22363 ( .A(n27570), .B(n26040), .C(n27572), .Y(n27684) );
  NOR2X1 U22364 ( .A(n27685), .B(n27686), .Y(n27263) );
  OAI22X1 U22365 ( .A(reg_A[82]), .B(n26036), .C(reg_A[74]), .D(n26981), .Y(
        n27686) );
  OAI21X1 U22366 ( .A(reg_A[66]), .B(n26982), .C(n26983), .Y(n27685) );
  AOI22X1 U22367 ( .A(n26050), .B(n27584), .C(reg_A[82]), .D(n27687), .Y(
        n27626) );
  NAND2X1 U22368 ( .A(n27688), .B(n27689), .Y(n27584) );
  AOI22X1 U22369 ( .A(n25838), .B(n26975), .C(n26160), .D(n27260), .Y(n27689)
         );
  OAI21X1 U22370 ( .A(n26131), .B(n26438), .C(n27690), .Y(n26975) );
  AOI22X1 U22371 ( .A(reg_A[66]), .B(n26513), .C(reg_A[82]), .D(n26134), .Y(
        n27690) );
  AOI22X1 U22372 ( .A(n26159), .B(n27691), .C(n26059), .D(n27505), .Y(n27688)
         );
  AOI22X1 U22373 ( .A(n26049), .B(n27616), .C(n27274), .D(n27551), .Y(n27625)
         );
  INVX1 U22374 ( .A(n27692), .Y(n27551) );
  AOI22X1 U22375 ( .A(reg_A[82]), .B(n27104), .C(reg_A[80]), .D(n27277), .Y(
        n27692) );
  OAI22X1 U22376 ( .A(reg_B[94]), .B(n27488), .C(n25584), .D(n26872), .Y(
        n27616) );
  NAND2X1 U22377 ( .A(reg_B[94]), .B(n26275), .Y(n26872) );
  NAND2X1 U22378 ( .A(reg_A[82]), .B(n26275), .Y(n27488) );
  INVX1 U22379 ( .A(n27353), .Y(n26049) );
  NAND2X1 U22380 ( .A(n26267), .B(n25976), .Y(n27353) );
  NAND3X1 U22381 ( .A(n27693), .B(n27694), .C(n27695), .Y(n27623) );
  NOR2X1 U22382 ( .A(n27696), .B(n27697), .Y(n27695) );
  OAI22X1 U22383 ( .A(n25583), .B(n25853), .C(n27698), .D(n25584), .Y(n27697)
         );
  NAND3X1 U22384 ( .A(n27699), .B(n27700), .C(n27701), .Y(n27696) );
  OAI21X1 U22385 ( .A(n27702), .B(n27703), .C(n25382), .Y(n27701) );
  INVX1 U22386 ( .A(n27704), .Y(n27703) );
  AOI22X1 U22387 ( .A(n27705), .B(n27706), .C(n27597), .D(n27205), .Y(n27704)
         );
  NOR2X1 U22388 ( .A(n27707), .B(reg_B[86]), .Y(n27205) );
  OAI22X1 U22389 ( .A(n27708), .B(n27058), .C(n27709), .D(n27061), .Y(n27702)
         );
  OAI21X1 U22390 ( .A(n27710), .B(n27711), .C(n25840), .Y(n27700) );
  NAND3X1 U22391 ( .A(n27712), .B(n27713), .C(n27714), .Y(n27711) );
  NOR2X1 U22392 ( .A(n27715), .B(n27716), .Y(n27714) );
  OAI22X1 U22393 ( .A(n25035), .B(n26107), .C(n25036), .D(n26547), .Y(n27716)
         );
  OAI21X1 U22394 ( .A(n25027), .B(n26101), .C(n27717), .Y(n27715) );
  AOI22X1 U22395 ( .A(reg_A[73]), .B(n25629), .C(reg_A[74]), .D(n25124), .Y(
        n27717) );
  AOI22X1 U22396 ( .A(reg_A[67]), .B(n25235), .C(reg_A[70]), .D(n25635), .Y(
        n27713) );
  AOI22X1 U22397 ( .A(reg_A[69]), .B(n25325), .C(reg_A[82]), .D(n25125), .Y(
        n27712) );
  NAND3X1 U22398 ( .A(n27718), .B(n27719), .C(n27720), .Y(n27710) );
  NOR2X1 U22399 ( .A(n27721), .B(n27722), .Y(n27720) );
  OAI22X1 U22400 ( .A(n25041), .B(n25864), .C(n25042), .D(n26094), .Y(n27722)
         );
  OAI21X1 U22401 ( .A(n25051), .B(n25853), .C(n27723), .Y(n27721) );
  AOI22X1 U22402 ( .A(reg_A[65]), .B(n25246), .C(reg_A[66]), .D(n25247), .Y(
        n27723) );
  AOI21X1 U22403 ( .A(reg_A[75]), .B(n25628), .C(n27724), .Y(n27719) );
  OAI22X1 U22404 ( .A(n25033), .B(n25863), .C(n25040), .D(n25584), .Y(n27724)
         );
  AOI22X1 U22405 ( .A(reg_A[78]), .B(n25071), .C(reg_A[77]), .D(n25123), .Y(
        n27718) );
  OAI21X1 U22406 ( .A(n27725), .B(n27726), .C(reg_A[81]), .Y(n27699) );
  AOI22X1 U22407 ( .A(reg_A[84]), .B(n25506), .C(reg_A[85]), .D(n25507), .Y(
        n27694) );
  AOI22X1 U22408 ( .A(reg_A[86]), .B(n25508), .C(reg_A[87]), .D(n25509), .Y(
        n27693) );
  OR2X1 U22409 ( .A(n27727), .B(n27728), .Y(result[81]) );
  NAND3X1 U22410 ( .A(n27729), .B(n27730), .C(n27731), .Y(n27728) );
  NOR2X1 U22411 ( .A(n27732), .B(n27733), .Y(n27731) );
  OAI21X1 U22412 ( .A(n27630), .B(n26950), .C(n27734), .Y(n27733) );
  OAI21X1 U22413 ( .A(n27735), .B(n27736), .C(n25203), .Y(n27734) );
  NAND3X1 U22414 ( .A(n27737), .B(n27738), .C(n27739), .Y(n27736) );
  AOI22X1 U22415 ( .A(reg_A[84]), .B(n27740), .C(reg_A[83]), .D(n27637), .Y(
        n27739) );
  OAI21X1 U22416 ( .A(n27741), .B(n27742), .C(n25044), .Y(n27738) );
  NAND2X1 U22417 ( .A(n27743), .B(n27744), .Y(n27742) );
  AOI22X1 U22418 ( .A(reg_A[91]), .B(n25637), .C(reg_A[95]), .D(n25234), .Y(
        n27744) );
  AOI22X1 U22419 ( .A(reg_A[93]), .B(n25635), .C(reg_A[94]), .D(n25325), .Y(
        n27743) );
  NAND2X1 U22420 ( .A(n27745), .B(n27746), .Y(n27741) );
  AOI22X1 U22421 ( .A(reg_A[88]), .B(n25628), .C(reg_A[90]), .D(n25629), .Y(
        n27746) );
  AOI22X1 U22422 ( .A(reg_A[89]), .B(n25124), .C(reg_A[92]), .D(n25222), .Y(
        n27745) );
  OAI21X1 U22423 ( .A(n27747), .B(n27748), .C(n25604), .Y(n27737) );
  NAND2X1 U22424 ( .A(n27749), .B(n27750), .Y(n27748) );
  AOI22X1 U22425 ( .A(reg_A[91]), .B(n25607), .C(reg_A[95]), .D(n25608), .Y(
        n27750) );
  AOI22X1 U22426 ( .A(reg_A[93]), .B(n25609), .C(reg_A[94]), .D(n25610), .Y(
        n27749) );
  NAND2X1 U22427 ( .A(n27751), .B(n27752), .Y(n27747) );
  AOI22X1 U22428 ( .A(reg_A[88]), .B(n25613), .C(reg_A[90]), .D(n25614), .Y(
        n27752) );
  AOI22X1 U22429 ( .A(reg_A[89]), .B(n25615), .C(reg_A[92]), .D(n25616), .Y(
        n27751) );
  OR2X1 U22430 ( .A(n27753), .B(n27754), .Y(n27735) );
  OAI22X1 U22431 ( .A(n25600), .B(n26039), .C(n27755), .D(n25965), .Y(n27754)
         );
  OAI21X1 U22432 ( .A(n27756), .B(n26215), .C(n27757), .Y(n27753) );
  AOI22X1 U22433 ( .A(reg_A[81]), .B(n27639), .C(reg_A[82]), .D(n25617), .Y(
        n27757) );
  AND2X1 U22434 ( .A(n27758), .B(n27759), .Y(n27630) );
  AOI22X1 U22435 ( .A(n25838), .B(n27114), .C(n26160), .D(n27393), .Y(n27759)
         );
  OAI21X1 U22436 ( .A(n26439), .B(n26131), .C(n27760), .Y(n27114) );
  AOI22X1 U22437 ( .A(n26513), .B(reg_A[65]), .C(reg_A[81]), .D(n26134), .Y(
        n27760) );
  AOI22X1 U22438 ( .A(n26159), .B(n27761), .C(n26059), .D(n27550), .Y(n27758)
         );
  OAI22X1 U22439 ( .A(n27762), .B(n27020), .C(n25652), .D(n26039), .Y(n27732)
         );
  AOI21X1 U22440 ( .A(reg_A[83]), .B(n25506), .C(n27763), .Y(n27730) );
  OAI21X1 U22441 ( .A(n25702), .B(n25965), .C(n27764), .Y(n27763) );
  OAI21X1 U22442 ( .A(n27726), .B(n27765), .C(reg_A[80]), .Y(n27764) );
  OAI21X1 U22443 ( .A(n27766), .B(n25342), .C(n27767), .Y(n27765) );
  NOR2X1 U22444 ( .A(reg_B[86]), .B(reg_B[87]), .Y(n27766) );
  OAI21X1 U22445 ( .A(n27278), .B(n27404), .C(n27768), .Y(n27726) );
  AOI21X1 U22446 ( .A(n27769), .B(n26267), .C(n27770), .Y(n27768) );
  INVX1 U22447 ( .A(n26381), .Y(n27769) );
  NAND2X1 U22448 ( .A(n26148), .B(n26275), .Y(n26381) );
  NAND2X1 U22449 ( .A(reg_B[87]), .B(n26186), .Y(n27404) );
  AOI22X1 U22450 ( .A(reg_A[84]), .B(n25507), .C(reg_A[85]), .D(n25508), .Y(
        n27729) );
  NAND3X1 U22451 ( .A(n27771), .B(n27772), .C(n27773), .Y(n27727) );
  NOR2X1 U22452 ( .A(n27774), .B(n27775), .Y(n27773) );
  OAI21X1 U22453 ( .A(n27776), .B(n26094), .C(n27777), .Y(n27775) );
  OAI21X1 U22454 ( .A(n25369), .B(n27778), .C(reg_A[64]), .Y(n27777) );
  NOR2X1 U22455 ( .A(n27779), .B(n27687), .Y(n27776) );
  NAND3X1 U22456 ( .A(n27780), .B(n27781), .C(n27782), .Y(n27774) );
  OAI21X1 U22457 ( .A(n27783), .B(n27784), .C(n25372), .Y(n27782) );
  OAI21X1 U22458 ( .A(n25984), .B(n27444), .C(n27528), .Y(n27784) );
  AOI22X1 U22459 ( .A(reg_A[80]), .B(n27597), .C(n26067), .D(n26223), .Y(
        n27528) );
  INVX1 U22460 ( .A(n27444), .Y(n26223) );
  NAND2X1 U22461 ( .A(reg_A[80]), .B(n25604), .Y(n27444) );
  OAI21X1 U22462 ( .A(n27661), .B(n26094), .C(n27785), .Y(n27783) );
  AOI22X1 U22463 ( .A(n25980), .B(n27786), .C(n27787), .D(n27788), .Y(n27785)
         );
  OAI21X1 U22464 ( .A(reg_B[91]), .B(n27789), .C(n27790), .Y(n27788) );
  INVX1 U22465 ( .A(n27791), .Y(n27790) );
  MUX2X1 U22466 ( .B(n27462), .A(n27664), .S(reg_B[94]), .Y(n27791) );
  OAI21X1 U22467 ( .A(reg_B[93]), .B(n27123), .C(n27792), .Y(n27462) );
  AOI21X1 U22468 ( .A(n27540), .B(n27793), .C(n27541), .Y(n27792) );
  INVX1 U22469 ( .A(n27794), .Y(n27541) );
  NAND3X1 U22470 ( .A(reg_B[91]), .B(n25853), .C(reg_B[93]), .Y(n27794) );
  INVX1 U22471 ( .A(n26306), .Y(n27793) );
  NOR2X1 U22472 ( .A(n26197), .B(reg_B[91]), .Y(n27540) );
  NOR2X1 U22473 ( .A(n27795), .B(n27796), .Y(n27123) );
  OAI22X1 U22474 ( .A(reg_A[73]), .B(n26131), .C(reg_A[81]), .D(n25894), .Y(
        n27796) );
  OAI21X1 U22475 ( .A(reg_A[65]), .B(n27027), .C(n27028), .Y(n27795) );
  NAND2X1 U22476 ( .A(n26061), .B(n25853), .Y(n27028) );
  NOR2X1 U22477 ( .A(n25895), .B(n26063), .Y(n26061) );
  AOI22X1 U22478 ( .A(n26518), .B(n26159), .C(n26160), .D(n27670), .Y(n27789)
         );
  OAI21X1 U22479 ( .A(reg_B[91]), .B(n27797), .C(n27664), .Y(n27786) );
  AOI22X1 U22480 ( .A(n25604), .B(n27798), .C(n27057), .D(n27799), .Y(n27661)
         );
  OAI21X1 U22481 ( .A(n27800), .B(n27801), .C(n25840), .Y(n27781) );
  NAND3X1 U22482 ( .A(n27802), .B(n27803), .C(n27804), .Y(n27801) );
  NOR2X1 U22483 ( .A(n27805), .B(n27806), .Y(n27804) );
  OAI22X1 U22484 ( .A(n25035), .B(n25851), .C(n25219), .D(n26101), .Y(n27806)
         );
  OAI21X1 U22485 ( .A(n25027), .B(n26256), .C(n27807), .Y(n27805) );
  AOI22X1 U22486 ( .A(reg_A[72]), .B(n25629), .C(reg_A[73]), .D(n25124), .Y(
        n27807) );
  AOI22X1 U22487 ( .A(reg_A[66]), .B(n25235), .C(reg_A[69]), .D(n25635), .Y(
        n27803) );
  AOI22X1 U22488 ( .A(reg_A[68]), .B(n25325), .C(reg_A[81]), .D(n25125), .Y(
        n27802) );
  NAND3X1 U22489 ( .A(n27808), .B(n27809), .C(n27810), .Y(n27800) );
  NOR2X1 U22490 ( .A(n27811), .B(n27812), .Y(n27810) );
  OAI22X1 U22491 ( .A(n25040), .B(n25864), .C(n25041), .D(n25865), .Y(n27812)
         );
  OAI21X1 U22492 ( .A(n25042), .B(n25584), .C(n27813), .Y(n27811) );
  AOI22X1 U22493 ( .A(reg_A[64]), .B(n25246), .C(reg_A[65]), .D(n25247), .Y(
        n27813) );
  AOI22X1 U22494 ( .A(reg_A[75]), .B(n25253), .C(reg_A[74]), .D(n25628), .Y(
        n27809) );
  AOI22X1 U22495 ( .A(reg_A[77]), .B(n25071), .C(reg_A[76]), .D(n25123), .Y(
        n27808) );
  OAI21X1 U22496 ( .A(n27814), .B(n27815), .C(n25382), .Y(n27780) );
  OAI22X1 U22497 ( .A(n27592), .B(n27816), .C(n27325), .D(n27059), .Y(n27815)
         );
  MUX2X1 U22498 ( .B(n27817), .A(n27103), .S(reg_B[86]), .Y(n27325) );
  NOR2X1 U22499 ( .A(n25965), .B(reg_B[87]), .Y(n27103) );
  INVX1 U22500 ( .A(n27595), .Y(n27817) );
  MUX2X1 U22501 ( .B(reg_A[85]), .A(reg_A[86]), .S(reg_B[87]), .Y(n27595) );
  INVX1 U22502 ( .A(n27818), .Y(n27816) );
  INVX1 U22503 ( .A(n27705), .Y(n27592) );
  OAI22X1 U22504 ( .A(n27593), .B(n27061), .C(n25874), .D(n27657), .Y(n27814)
         );
  AOI21X1 U22505 ( .A(reg_A[84]), .B(reg_B[87]), .C(n27102), .Y(n27593) );
  INVX1 U22506 ( .A(n27331), .Y(n27102) );
  NAND2X1 U22507 ( .A(reg_A[83]), .B(n27057), .Y(n27331) );
  INVX1 U22508 ( .A(n27819), .Y(n27772) );
  OAI22X1 U22509 ( .A(n27820), .B(n26533), .C(n27821), .D(n27822), .Y(n27819)
         );
  INVX1 U22510 ( .A(n27823), .Y(n26533) );
  INVX1 U22511 ( .A(n27824), .Y(n27771) );
  OAI22X1 U22512 ( .A(n27825), .B(n27456), .C(n27826), .D(n27571), .Y(n27824)
         );
  OAI21X1 U22513 ( .A(reg_B[2]), .B(n27384), .C(n27827), .Y(n27456) );
  AOI21X1 U22514 ( .A(n27570), .B(n26216), .C(n27572), .Y(n27827) );
  AND2X1 U22515 ( .A(n27828), .B(n25853), .Y(n27572) );
  NOR2X1 U22516 ( .A(n27829), .B(n27830), .Y(n27384) );
  OAI22X1 U22517 ( .A(reg_A[81]), .B(n25063), .C(reg_A[73]), .D(n26981), .Y(
        n27830) );
  OAI21X1 U22518 ( .A(reg_A[65]), .B(n26982), .C(n26983), .Y(n27829) );
  NAND2X1 U22519 ( .A(n26662), .B(n25853), .Y(n26983) );
  NAND3X1 U22520 ( .A(n27831), .B(n27832), .C(n27833), .Y(result[80]) );
  NOR2X1 U22521 ( .A(n27834), .B(n27835), .Y(n27833) );
  NAND2X1 U22522 ( .A(n27836), .B(n27837), .Y(n27835) );
  INVX1 U22523 ( .A(n27838), .Y(n27837) );
  OAI21X1 U22524 ( .A(n27839), .B(n27822), .C(n27840), .Y(n27838) );
  INVX1 U22525 ( .A(n27841), .Y(n27840) );
  OAI21X1 U22526 ( .A(reg_B[91]), .B(n27842), .C(n27843), .Y(n27841) );
  OAI21X1 U22527 ( .A(n27779), .B(n27844), .C(reg_A[80]), .Y(n27843) );
  OAI21X1 U22528 ( .A(n26147), .B(n26377), .C(n27845), .Y(n27779) );
  AOI21X1 U22529 ( .A(n27274), .B(n27104), .C(n27045), .Y(n27845) );
  INVX1 U22530 ( .A(n27846), .Y(n27045) );
  NAND3X1 U22531 ( .A(n25382), .B(n27057), .C(n27799), .Y(n27846) );
  INVX1 U22532 ( .A(n27553), .Y(n27274) );
  NAND2X1 U22533 ( .A(n26186), .B(n27057), .Y(n27553) );
  INVX1 U22534 ( .A(reg_B[87]), .Y(n27057) );
  AOI22X1 U22535 ( .A(n26014), .B(n27847), .C(n27848), .D(n26125), .Y(n27842)
         );
  INVX1 U22536 ( .A(n27797), .Y(n27848) );
  OAI21X1 U22537 ( .A(reg_B[94]), .B(n27538), .C(n27849), .Y(n27797) );
  AOI22X1 U22538 ( .A(n27850), .B(n26159), .C(n26160), .D(n26133), .Y(n27849)
         );
  MUX2X1 U22539 ( .B(reg_A[70]), .A(reg_A[78]), .S(n26063), .Y(n26133) );
  MUX2X1 U22540 ( .B(reg_A[74]), .A(reg_A[66]), .S(reg_B[92]), .Y(n27850) );
  AOI21X1 U22541 ( .A(n25584), .B(n26275), .C(n27851), .Y(n27538) );
  OAI22X1 U22542 ( .A(n26197), .B(n26415), .C(n26199), .D(reg_A[72]), .Y(
        n27851) );
  MUX2X1 U22543 ( .B(n25863), .A(n26107), .S(reg_B[92]), .Y(n26415) );
  OAI21X1 U22544 ( .A(n25896), .B(n26337), .C(n27852), .Y(n27847) );
  AOI22X1 U22545 ( .A(n26306), .B(n26160), .C(n26518), .D(n26059), .Y(n27852)
         );
  MUX2X1 U22546 ( .B(n26103), .A(n25851), .S(reg_B[92]), .Y(n26518) );
  MUX2X1 U22547 ( .B(n26286), .A(n25856), .S(reg_B[92]), .Y(n26306) );
  INVX1 U22548 ( .A(n27670), .Y(n25896) );
  MUX2X1 U22549 ( .B(n25864), .A(n26101), .S(reg_B[92]), .Y(n27670) );
  INVX1 U22550 ( .A(n26298), .Y(n26014) );
  OAI21X1 U22551 ( .A(reg_B[3]), .B(n27578), .C(n27853), .Y(n27822) );
  AOI22X1 U22552 ( .A(n26530), .B(n27854), .C(n25026), .D(n26040), .Y(n27853)
         );
  MUX2X1 U22553 ( .B(reg_A[70]), .A(reg_A[78]), .S(n26596), .Y(n26040) );
  INVX1 U22554 ( .A(n27855), .Y(n27854) );
  INVX1 U22555 ( .A(n27856), .Y(n27578) );
  OAI21X1 U22556 ( .A(reg_A[80]), .B(n27857), .C(n27858), .Y(n27856) );
  AOI22X1 U22557 ( .A(n27859), .B(n26547), .C(reg_B[2]), .D(n26367), .Y(n27858) );
  AOI22X1 U22558 ( .A(n27860), .B(reg_A[73]), .C(n27861), .D(reg_A[65]), .Y(
        n27836) );
  NAND3X1 U22559 ( .A(n27862), .B(n27863), .C(n27864), .Y(n27834) );
  AOI21X1 U22560 ( .A(n25382), .B(n27865), .C(n27866), .Y(n27864) );
  OAI21X1 U22561 ( .A(n26298), .B(n27867), .C(n27868), .Y(n27866) );
  OAI21X1 U22562 ( .A(n27869), .B(n27870), .C(n25840), .Y(n27868) );
  NAND3X1 U22563 ( .A(n27871), .B(n27872), .C(n27873), .Y(n27870) );
  NOR2X1 U22564 ( .A(n27874), .B(n27875), .Y(n27873) );
  OAI22X1 U22565 ( .A(n25043), .B(n25584), .C(n25039), .D(n25851), .Y(n27875)
         );
  OAI22X1 U22566 ( .A(n25064), .B(n26107), .C(n25065), .D(n25855), .Y(n27874)
         );
  AOI22X1 U22567 ( .A(reg_A[72]), .B(n25124), .C(reg_A[69]), .D(n25222), .Y(
        n27872) );
  AOI22X1 U22568 ( .A(reg_A[70]), .B(n25637), .C(reg_A[66]), .D(n25234), .Y(
        n27871) );
  NAND3X1 U22569 ( .A(n27876), .B(n27877), .C(n27878), .Y(n27869) );
  NOR2X1 U22570 ( .A(n27879), .B(n27880), .Y(n27878) );
  OAI22X1 U22571 ( .A(n25033), .B(n26438), .C(n25040), .D(n25865), .Y(n27880)
         );
  OAI21X1 U22572 ( .A(n25041), .B(n26286), .C(n27881), .Y(n27879) );
  AOI22X1 U22573 ( .A(reg_A[64]), .B(n25247), .C(reg_A[79]), .D(n25135), .Y(
        n27881) );
  AOI22X1 U22574 ( .A(reg_A[73]), .B(n25628), .C(reg_A[76]), .D(n25068), .Y(
        n27877) );
  AOI22X1 U22575 ( .A(reg_A[75]), .B(n25123), .C(reg_A[71]), .D(n25629), .Y(
        n27876) );
  NAND2X1 U22576 ( .A(n26159), .B(n27882), .Y(n27867) );
  NAND2X1 U22577 ( .A(n27883), .B(n27884), .Y(n27865) );
  INVX1 U22578 ( .A(n27885), .Y(n27884) );
  OAI22X1 U22579 ( .A(n27657), .B(n26094), .C(n27061), .D(n27708), .Y(n27885)
         );
  MUX2X1 U22580 ( .B(reg_A[82]), .A(reg_A[83]), .S(reg_B[87]), .Y(n27708) );
  NAND2X1 U22581 ( .A(n27277), .B(n25589), .Y(n27061) );
  NOR2X1 U22582 ( .A(n27275), .B(reg_B[85]), .Y(n27277) );
  NAND2X1 U22583 ( .A(reg_B[87]), .B(n27799), .Y(n27657) );
  INVX1 U22584 ( .A(n27058), .Y(n27799) );
  NAND2X1 U22585 ( .A(n27104), .B(n25029), .Y(n27058) );
  INVX1 U22586 ( .A(n27278), .Y(n27104) );
  NAND2X1 U22587 ( .A(n27318), .B(n27275), .Y(n27278) );
  INVX1 U22588 ( .A(reg_B[85]), .Y(n27318) );
  AOI22X1 U22589 ( .A(n27886), .B(n27705), .C(n27597), .D(n27422), .Y(n27883)
         );
  MUX2X1 U22590 ( .B(n27707), .A(n27709), .S(n27275), .Y(n27422) );
  INVX1 U22591 ( .A(reg_B[86]), .Y(n27275) );
  MUX2X1 U22592 ( .B(reg_A[84]), .A(reg_A[85]), .S(reg_B[87]), .Y(n27709) );
  MUX2X1 U22593 ( .B(reg_A[86]), .A(reg_A[87]), .S(reg_B[87]), .Y(n27707) );
  INVX1 U22594 ( .A(n27059), .Y(n27597) );
  NAND2X1 U22595 ( .A(reg_B[85]), .B(n25029), .Y(n27059) );
  OAI21X1 U22596 ( .A(reg_B[91]), .B(n25403), .C(n25052), .Y(n27705) );
  OAI21X1 U22597 ( .A(n27887), .B(n27888), .C(n25730), .Y(n27863) );
  NAND3X1 U22598 ( .A(n27889), .B(n27890), .C(n27891), .Y(n27888) );
  NOR2X1 U22599 ( .A(n27892), .B(n27893), .Y(n27891) );
  OAI22X1 U22600 ( .A(n25736), .B(n25584), .C(n25737), .D(n25881), .Y(n27893)
         );
  OAI22X1 U22601 ( .A(n25738), .B(n25882), .C(n25739), .D(n25873), .Y(n27892)
         );
  AOI22X1 U22602 ( .A(reg_A[88]), .B(n25615), .C(reg_A[91]), .D(n25616), .Y(
        n27890) );
  AOI22X1 U22603 ( .A(reg_A[90]), .B(n25607), .C(reg_A[94]), .D(n25608), .Y(
        n27889) );
  NAND3X1 U22604 ( .A(n27894), .B(n27895), .C(n27896), .Y(n27887) );
  NOR2X1 U22605 ( .A(n27897), .B(n27898), .Y(n27896) );
  OAI22X1 U22606 ( .A(n25061), .B(n26039), .C(n25746), .D(n25874), .Y(n27898)
         );
  OAI22X1 U22607 ( .A(n25747), .B(n25875), .C(n25748), .D(n26094), .Y(n27897)
         );
  AOI22X1 U22608 ( .A(reg_A[87]), .B(n25613), .C(reg_A[84]), .D(n25749), .Y(
        n27895) );
  AOI22X1 U22609 ( .A(reg_A[85]), .B(n25750), .C(reg_A[89]), .D(n25614), .Y(
        n27894) );
  OAI21X1 U22610 ( .A(n27899), .B(n27900), .C(n25310), .Y(n27862) );
  NAND3X1 U22611 ( .A(n27901), .B(n27902), .C(n27903), .Y(n27900) );
  NOR2X1 U22612 ( .A(n27904), .B(n27905), .Y(n27903) );
  OAI22X1 U22613 ( .A(n25043), .B(n25584), .C(n25229), .D(n25881), .Y(n27905)
         );
  OAI22X1 U22614 ( .A(n25064), .B(n25882), .C(n25482), .D(n25873), .Y(n27904)
         );
  AOI22X1 U22615 ( .A(reg_A[88]), .B(n25124), .C(reg_A[91]), .D(n25222), .Y(
        n27902) );
  AOI22X1 U22616 ( .A(reg_A[90]), .B(n25637), .C(reg_A[94]), .D(n25234), .Y(
        n27901) );
  NAND3X1 U22617 ( .A(n27906), .B(n27907), .C(n27908), .Y(n27899) );
  NOR2X1 U22618 ( .A(n27909), .B(n27910), .Y(n27908) );
  OAI22X1 U22619 ( .A(n25033), .B(n26039), .C(n25040), .D(n25874), .Y(n27910)
         );
  OAI22X1 U22620 ( .A(n25041), .B(n25875), .C(n25042), .D(n26094), .Y(n27909)
         );
  AOI22X1 U22621 ( .A(reg_A[87]), .B(n25628), .C(reg_A[84]), .D(n25068), .Y(
        n27907) );
  AOI22X1 U22622 ( .A(reg_A[85]), .B(n25123), .C(reg_A[89]), .D(n25629), .Y(
        n27906) );
  NOR2X1 U22623 ( .A(n27911), .B(n27912), .Y(n27832) );
  OAI22X1 U22624 ( .A(n27913), .B(n27020), .C(n27762), .D(n26950), .Y(n27912)
         );
  AND2X1 U22625 ( .A(n27914), .B(n27915), .Y(n27762) );
  AOI22X1 U22626 ( .A(n25838), .B(n27260), .C(n26159), .D(n27916), .Y(n27915)
         );
  OAI21X1 U22627 ( .A(n26131), .B(n26547), .C(n27917), .Y(n27260) );
  AOI22X1 U22628 ( .A(reg_A[64]), .B(n26513), .C(n26134), .D(reg_A[80]), .Y(
        n27917) );
  INVX1 U22629 ( .A(n27027), .Y(n26513) );
  AOI22X1 U22630 ( .A(n26160), .B(n27505), .C(n26059), .D(n27691), .Y(n27914)
         );
  INVX1 U22631 ( .A(n27918), .Y(n27913) );
  OAI21X1 U22632 ( .A(n27919), .B(n25853), .C(n27920), .Y(n27911) );
  AOI22X1 U22633 ( .A(n27921), .B(n27922), .C(n26928), .D(n27923), .Y(n27920)
         );
  OAI21X1 U22634 ( .A(n26944), .B(n26215), .C(n27924), .Y(n27923) );
  AOI22X1 U22635 ( .A(reg_A[86]), .B(n26010), .C(reg_A[87]), .D(n26002), .Y(
        n27924) );
  OAI21X1 U22636 ( .A(n27925), .B(n27571), .C(n27926), .Y(n27922) );
  AOI22X1 U22637 ( .A(n27927), .B(n26008), .C(n27823), .D(n25751), .Y(n27926)
         );
  INVX1 U22638 ( .A(n25901), .Y(n27571) );
  MUX2X1 U22639 ( .B(n25864), .A(n26101), .S(reg_B[1]), .Y(n25901) );
  NOR2X1 U22640 ( .A(n27928), .B(n27929), .Y(n27831) );
  OAI22X1 U22641 ( .A(n25717), .B(n25874), .C(n25718), .D(n25875), .Y(n27929)
         );
  OAI21X1 U22642 ( .A(n25719), .B(n26094), .C(n27930), .Y(n27928) );
  AOI22X1 U22643 ( .A(n27537), .B(n25932), .C(reg_A[84]), .D(n25722), .Y(
        n27930) );
  OR2X1 U22644 ( .A(n27931), .B(n27932), .Y(result[7]) );
  NAND3X1 U22645 ( .A(n27933), .B(n27934), .C(n27935), .Y(n27932) );
  NOR2X1 U22646 ( .A(n27936), .B(n27937), .Y(n27935) );
  OAI21X1 U22647 ( .A(n27938), .B(n25146), .C(n27939), .Y(n27937) );
  AOI22X1 U22648 ( .A(reg_A[8]), .B(n27940), .C(reg_A[15]), .D(n25302), .Y(
        n27939) );
  OR2X1 U22649 ( .A(n27941), .B(n27942), .Y(n27936) );
  OAI21X1 U22650 ( .A(n27943), .B(n27944), .C(n27945), .Y(n27942) );
  OAI21X1 U22651 ( .A(n27946), .B(n27947), .C(n25310), .Y(n27945) );
  NAND3X1 U22652 ( .A(n27948), .B(n27949), .C(n27950), .Y(n27947) );
  NOR2X1 U22653 ( .A(n27951), .B(n27952), .Y(n27950) );
  OAI22X1 U22654 ( .A(n27953), .B(n25219), .C(n25224), .D(n25473), .Y(n27952)
         );
  OAI22X1 U22655 ( .A(n25250), .B(n25223), .C(n27954), .D(n25320), .Y(n27951)
         );
  AOI22X1 U22656 ( .A(reg_A[21]), .B(n25234), .C(reg_A[22]), .D(n25235), .Y(
        n27949) );
  AOI22X1 U22657 ( .A(n25635), .B(reg_A[19]), .C(n25325), .D(reg_A[20]), .Y(
        n27948) );
  NAND3X1 U22658 ( .A(n27955), .B(n27956), .C(n27957), .Y(n27946) );
  NOR2X1 U22659 ( .A(n27958), .B(n27959), .Y(n27957) );
  OAI22X1 U22660 ( .A(n27960), .B(n25331), .C(n27961), .D(n25243), .Y(n27959)
         );
  OAI22X1 U22661 ( .A(n25048), .B(n26714), .C(n25047), .D(n27962), .Y(n27958)
         );
  AOI22X1 U22662 ( .A(reg_A[29]), .B(n25242), .C(n25338), .D(reg_A[30]), .Y(
        n27956) );
  AOI22X1 U22663 ( .A(n25339), .B(reg_A[27]), .C(n25257), .D(reg_A[28]), .Y(
        n27955) );
  OAI22X1 U22664 ( .A(n25945), .B(n27963), .C(n27964), .D(n25132), .Y(n27941)
         );
  NOR2X1 U22665 ( .A(n27965), .B(n27966), .Y(n27934) );
  OAI22X1 U22666 ( .A(n25295), .B(n25206), .C(n25297), .D(n25255), .Y(n27966)
         );
  OAI22X1 U22667 ( .A(n27511), .B(n27967), .C(n27968), .D(n25147), .Y(n27965)
         );
  NOR2X1 U22668 ( .A(n27969), .B(n27970), .Y(n27933) );
  OAI21X1 U22669 ( .A(n27971), .B(n25208), .C(n27972), .Y(n27970) );
  OAI21X1 U22670 ( .A(n27973), .B(n27974), .C(n25170), .Y(n27972) );
  OAI21X1 U22671 ( .A(n25132), .B(n27975), .C(n27976), .Y(n27974) );
  OAI21X1 U22672 ( .A(n27977), .B(n27978), .C(n25044), .Y(n27976) );
  NOR2X1 U22673 ( .A(n27979), .B(n25264), .Y(n27977) );
  INVX1 U22674 ( .A(n27980), .Y(n27975) );
  OAI21X1 U22675 ( .A(n27981), .B(n27982), .C(n27983), .Y(n27973) );
  NAND3X1 U22676 ( .A(n27984), .B(reg_A[5]), .C(n27985), .Y(n27983) );
  AOI22X1 U22677 ( .A(n27985), .B(reg_A[1]), .C(n27986), .D(reg_A[3]), .Y(
        n27981) );
  NAND3X1 U22678 ( .A(n27987), .B(n27988), .C(n27989), .Y(n27931) );
  NOR2X1 U22679 ( .A(n27990), .B(n27991), .Y(n27989) );
  INVX1 U22680 ( .A(n27992), .Y(n27991) );
  AOI21X1 U22681 ( .A(n27978), .B(n25932), .C(n27993), .Y(n27992) );
  OAI22X1 U22682 ( .A(n25194), .B(n27994), .C(n27995), .D(n25130), .Y(n27993)
         );
  OAI21X1 U22683 ( .A(n26757), .B(n25262), .C(n27996), .Y(n27978) );
  AOI22X1 U22684 ( .A(n25142), .B(n26760), .C(n25258), .D(n26762), .Y(n27996)
         );
  NAND2X1 U22685 ( .A(n27997), .B(n27998), .Y(n27990) );
  AOI22X1 U22686 ( .A(n27999), .B(n27155), .C(n25999), .D(n28000), .Y(n27998)
         );
  OAI21X1 U22687 ( .A(n25754), .B(n25177), .C(n28001), .Y(n28000) );
  AOI22X1 U22688 ( .A(reg_A[6]), .B(n26007), .C(n26009), .D(reg_A[5]), .Y(
        n28001) );
  OAI21X1 U22689 ( .A(n26730), .B(n26692), .C(n28002), .Y(n27999) );
  AOI22X1 U22690 ( .A(n25172), .B(n25160), .C(n26733), .D(n26735), .Y(n28002)
         );
  INVX1 U22691 ( .A(n25169), .Y(n26730) );
  AOI22X1 U22692 ( .A(n26504), .B(n28003), .C(n28004), .D(reg_A[4]), .Y(n27997) );
  OAI21X1 U22693 ( .A(n28005), .B(n28006), .C(n28007), .Y(n28003) );
  AOI22X1 U22694 ( .A(n28008), .B(n27986), .C(n28009), .D(n28010), .Y(n28007)
         );
  MUX2X1 U22695 ( .B(n25132), .A(n25130), .S(reg_B[5]), .Y(n28008) );
  INVX1 U22696 ( .A(n28011), .Y(n28006) );
  NOR2X1 U22697 ( .A(n28012), .B(n28013), .Y(n27988) );
  OAI21X1 U22698 ( .A(n28014), .B(n25087), .C(n28015), .Y(n28013) );
  OAI21X1 U22699 ( .A(n28016), .B(n28017), .C(n25119), .Y(n28015) );
  OAI21X1 U22700 ( .A(n25132), .B(n25228), .C(n28018), .Y(n28017) );
  AOI22X1 U22701 ( .A(n25075), .B(reg_A[3]), .C(n25123), .D(reg_A[2]), .Y(
        n28018) );
  NAND2X1 U22702 ( .A(n28019), .B(n28020), .Y(n28016) );
  AOI22X1 U22703 ( .A(n25135), .B(reg_A[6]), .C(n25136), .D(reg_A[4]), .Y(
        n28020) );
  AOI22X1 U22704 ( .A(n25252), .B(reg_A[5]), .C(n25253), .D(reg_A[1]), .Y(
        n28019) );
  AND2X1 U22705 ( .A(n28021), .B(n28022), .Y(n28014) );
  AOI21X1 U22706 ( .A(n28023), .B(n28024), .C(n28025), .Y(n28022) );
  OAI21X1 U22707 ( .A(n28026), .B(n28027), .C(n28028), .Y(n28025) );
  OAI21X1 U22708 ( .A(n28029), .B(n28030), .C(n25044), .Y(n28028) );
  OAI22X1 U22709 ( .A(n28031), .B(n25099), .C(n28032), .D(n28033), .Y(n28030)
         );
  OAI21X1 U22710 ( .A(n28034), .B(n25106), .C(n28035), .Y(n28029) );
  AOI22X1 U22711 ( .A(n25110), .B(n28036), .C(reg_B[27]), .D(n28037), .Y(
        n28035) );
  NAND2X1 U22712 ( .A(n25116), .B(reg_A[15]), .Y(n28027) );
  AOI22X1 U22713 ( .A(n28038), .B(n28039), .C(reg_A[7]), .D(n28040), .Y(n28021) );
  OAI21X1 U22714 ( .A(n28041), .B(n28042), .C(n28043), .Y(n28012) );
  OAI21X1 U22715 ( .A(n28044), .B(n28045), .C(n27067), .Y(n28043) );
  OAI21X1 U22716 ( .A(n25132), .B(n25736), .C(n28046), .Y(n28045) );
  AOI22X1 U22717 ( .A(n25749), .B(reg_A[3]), .C(n25750), .D(reg_A[2]), .Y(
        n28046) );
  NAND2X1 U22718 ( .A(n28047), .B(n28048), .Y(n28044) );
  AOI22X1 U22719 ( .A(reg_A[6]), .B(n26803), .C(n26804), .D(reg_A[4]), .Y(
        n28048) );
  AOI22X1 U22720 ( .A(n26927), .B(reg_A[5]), .C(reg_A[1]), .D(n26878), .Y(
        n28047) );
  OR2X1 U22721 ( .A(n26151), .B(n28049), .Y(n28042) );
  AOI21X1 U22722 ( .A(n28050), .B(reg_A[2]), .C(n28051), .Y(n27987) );
  OAI21X1 U22723 ( .A(n28052), .B(n28053), .C(n28054), .Y(n28051) );
  OAI21X1 U22724 ( .A(n28055), .B(n28056), .C(reg_A[0]), .Y(n28054) );
  OAI21X1 U22725 ( .A(n25194), .B(n28057), .C(n28058), .Y(n28056) );
  OR2X1 U22726 ( .A(n28059), .B(n28060), .Y(result[79]) );
  NAND3X1 U22727 ( .A(n28061), .B(n28062), .C(n28063), .Y(n28060) );
  NOR2X1 U22728 ( .A(n28064), .B(n28065), .Y(n28063) );
  OAI21X1 U22729 ( .A(n28066), .B(n25853), .C(n28067), .Y(n28065) );
  MUX2X1 U22730 ( .B(n28068), .A(n28069), .S(reg_B[78]), .Y(n28067) );
  NOR2X1 U22731 ( .A(n28070), .B(n25032), .Y(n28068) );
  AOI22X1 U22732 ( .A(n28071), .B(reg_B[77]), .C(n28072), .D(n28073), .Y(
        n28070) );
  NAND2X1 U22733 ( .A(n28074), .B(n28075), .Y(n28064) );
  OAI21X1 U22734 ( .A(n28076), .B(n28077), .C(n25999), .Y(n28075) );
  NAND2X1 U22735 ( .A(n28078), .B(n28079), .Y(n28077) );
  AOI22X1 U22736 ( .A(reg_A[72]), .B(n26002), .C(reg_A[75]), .D(n26003), .Y(
        n28079) );
  AOI22X1 U22737 ( .A(reg_A[74]), .B(n25751), .C(reg_A[79]), .D(n26004), .Y(
        n28078) );
  NAND2X1 U22738 ( .A(n28080), .B(n28081), .Y(n28076) );
  AOI22X1 U22739 ( .A(reg_A[78]), .B(n26007), .C(reg_A[76]), .D(n26008), .Y(
        n28081) );
  AOI22X1 U22740 ( .A(reg_A[77]), .B(n26009), .C(reg_A[73]), .D(n26010), .Y(
        n28080) );
  AOI22X1 U22741 ( .A(reg_A[79]), .B(n28082), .C(n28083), .D(n28084), .Y(
        n28074) );
  AOI21X1 U22742 ( .A(n25932), .B(n28085), .C(n28086), .Y(n28062) );
  OAI21X1 U22743 ( .A(n28087), .B(n28088), .C(n28089), .Y(n28086) );
  OAI21X1 U22744 ( .A(n28090), .B(n28091), .C(n26480), .Y(n28089) );
  OAI22X1 U22745 ( .A(n28092), .B(n28093), .C(n28094), .D(n25964), .Y(n28091)
         );
  OAI21X1 U22746 ( .A(n28095), .B(n26997), .C(n28096), .Y(n28090) );
  NAND3X1 U22747 ( .A(reg_B[91]), .B(n27798), .C(reg_A[95]), .Y(n28096) );
  INVX1 U22748 ( .A(n26377), .Y(n27798) );
  AOI21X1 U22749 ( .A(reg_A[79]), .B(n28097), .C(n28098), .Y(n28087) );
  OAI21X1 U22750 ( .A(n28099), .B(n25697), .C(n28100), .Y(n28098) );
  NAND3X1 U22751 ( .A(reg_A[75]), .B(n28101), .C(reg_B[77]), .Y(n28100) );
  OAI21X1 U22752 ( .A(n28102), .B(n25697), .C(n25031), .Y(n28101) );
  AOI22X1 U22753 ( .A(n28103), .B(reg_A[71]), .C(n28104), .D(reg_A[67]), .Y(
        n28099) );
  OAI21X1 U22754 ( .A(n28105), .B(n28106), .C(n28107), .Y(n28097) );
  INVX1 U22755 ( .A(n28108), .Y(n28106) );
  NAND2X1 U22756 ( .A(n28109), .B(n28110), .Y(n28085) );
  AOI21X1 U22757 ( .A(n25984), .B(n28111), .C(n28112), .Y(n28110) );
  OAI21X1 U22758 ( .A(n28113), .B(n26169), .C(n27664), .Y(n28112) );
  NOR2X1 U22759 ( .A(n28114), .B(n28115), .Y(n28113) );
  OAI21X1 U22760 ( .A(n25964), .B(n26101), .C(n28116), .Y(n28111) );
  AOI22X1 U22761 ( .A(reg_B[93]), .B(n27761), .C(reg_A[79]), .D(n26057), .Y(
        n28116) );
  AOI22X1 U22762 ( .A(n26148), .B(n28117), .C(n26276), .D(n28118), .Y(n28109)
         );
  AOI21X1 U22763 ( .A(n28119), .B(n26262), .C(n28120), .Y(n28061) );
  OAI22X1 U22764 ( .A(n25945), .B(n28121), .C(n26103), .D(n28122), .Y(n28120)
         );
  INVX1 U22765 ( .A(n28123), .Y(n28119) );
  NAND3X1 U22766 ( .A(n28124), .B(n28125), .C(n28126), .Y(n28059) );
  NOR2X1 U22767 ( .A(n28127), .B(n28128), .Y(n28126) );
  OAI21X1 U22768 ( .A(n28129), .B(n28130), .C(n28131), .Y(n28128) );
  AOI22X1 U22769 ( .A(n28132), .B(n28133), .C(n28134), .D(n25935), .Y(n28131)
         );
  OAI21X1 U22770 ( .A(n28135), .B(n26583), .C(n28136), .Y(n28127) );
  AOI22X1 U22771 ( .A(n26281), .B(n27918), .C(n28137), .D(n28138), .Y(n28136)
         );
  NAND2X1 U22772 ( .A(n28139), .B(n28140), .Y(n27918) );
  AOI22X1 U22773 ( .A(n25838), .B(n27393), .C(n26159), .D(n27882), .Y(n28140)
         );
  OAI22X1 U22774 ( .A(n26131), .B(n26101), .C(n25894), .D(n25864), .Y(n27393)
         );
  AOI22X1 U22775 ( .A(n26160), .B(n27550), .C(n26059), .D(n27761), .Y(n28139)
         );
  NOR2X1 U22776 ( .A(n26896), .B(n25697), .Y(n26281) );
  NOR2X1 U22777 ( .A(n28141), .B(n28142), .Y(n28125) );
  OAI21X1 U22778 ( .A(n28143), .B(n28144), .C(n28145), .Y(n28142) );
  OAI21X1 U22779 ( .A(n28146), .B(n28147), .C(n25119), .Y(n28145) );
  NAND3X1 U22780 ( .A(n28148), .B(n28149), .C(n28150), .Y(n28147) );
  AOI21X1 U22781 ( .A(reg_A[79]), .B(n25125), .C(n28151), .Y(n28150) );
  OAI22X1 U22782 ( .A(n25039), .B(n25884), .C(n25231), .D(n25851), .Y(n28151)
         );
  AOI22X1 U22783 ( .A(reg_A[71]), .B(n25124), .C(reg_A[68]), .D(n25222), .Y(
        n28149) );
  AOI22X1 U22784 ( .A(reg_A[69]), .B(n25637), .C(reg_A[65]), .D(n25234), .Y(
        n28148) );
  NAND3X1 U22785 ( .A(n28152), .B(n28153), .C(n28154), .Y(n28146) );
  NOR2X1 U22786 ( .A(n28155), .B(n28156), .Y(n28154) );
  OAI22X1 U22787 ( .A(n25033), .B(n26439), .C(n25133), .D(n26286), .Y(n28156)
         );
  OAI22X1 U22788 ( .A(n25041), .B(n25863), .C(n25042), .D(n25865), .Y(n28155)
         );
  AOI22X1 U22789 ( .A(reg_A[72]), .B(n25628), .C(reg_A[75]), .D(n25066), .Y(
        n28153) );
  AOI22X1 U22790 ( .A(reg_A[74]), .B(n25123), .C(reg_A[70]), .D(n25629), .Y(
        n28152) );
  AOI22X1 U22791 ( .A(n26267), .B(n28157), .C(n26186), .D(n28158), .Y(n28143)
         );
  INVX1 U22792 ( .A(n28159), .Y(n28141) );
  OAI21X1 U22793 ( .A(n28160), .B(n28161), .C(n25918), .Y(n28159) );
  NAND3X1 U22794 ( .A(n28162), .B(n28163), .C(n28164), .Y(n28161) );
  NOR2X1 U22795 ( .A(n28165), .B(n28166), .Y(n28164) );
  OAI22X1 U22796 ( .A(n25736), .B(n25864), .C(n25737), .D(n25884), .Y(n28166)
         );
  OAI22X1 U22797 ( .A(n25738), .B(n25851), .C(n25739), .D(n25853), .Y(n28165)
         );
  AOI22X1 U22798 ( .A(reg_A[71]), .B(n25615), .C(reg_A[68]), .D(n25616), .Y(
        n28163) );
  AOI22X1 U22799 ( .A(reg_A[69]), .B(n25607), .C(reg_A[65]), .D(n25608), .Y(
        n28162) );
  NAND3X1 U22800 ( .A(n28167), .B(n28168), .C(n28169), .Y(n28160) );
  NOR2X1 U22801 ( .A(n28170), .B(n28171), .Y(n28169) );
  OAI22X1 U22802 ( .A(n25745), .B(n26439), .C(n25746), .D(n26286), .Y(n28171)
         );
  OAI22X1 U22803 ( .A(n25747), .B(n25863), .C(n25748), .D(n25865), .Y(n28170)
         );
  AOI22X1 U22804 ( .A(reg_A[72]), .B(n25613), .C(reg_A[75]), .D(n25749), .Y(
        n28168) );
  AOI22X1 U22805 ( .A(reg_A[74]), .B(n25750), .C(reg_A[70]), .D(n25614), .Y(
        n28167) );
  AOI21X1 U22806 ( .A(reg_A[78]), .B(n28172), .C(n28173), .Y(n28124) );
  OAI21X1 U22807 ( .A(n28174), .B(n26438), .C(n28175), .Y(n28173) );
  OAI21X1 U22808 ( .A(n28176), .B(n28177), .C(n25310), .Y(n28175) );
  NAND3X1 U22809 ( .A(n28178), .B(n28179), .C(n28180), .Y(n28177) );
  NOR2X1 U22810 ( .A(n28181), .B(n28182), .Y(n28180) );
  OAI22X1 U22811 ( .A(n25043), .B(n25864), .C(n25039), .D(n25882), .Y(n28182)
         );
  OAI22X1 U22812 ( .A(n25064), .B(n25973), .C(n25482), .D(n25883), .Y(n28181)
         );
  AOI22X1 U22813 ( .A(reg_A[88]), .B(n25629), .C(reg_A[90]), .D(n25222), .Y(
        n28179) );
  AOI22X1 U22814 ( .A(reg_A[89]), .B(n25637), .C(reg_A[93]), .D(n25234), .Y(
        n28178) );
  NAND3X1 U22815 ( .A(n28183), .B(n28184), .C(n28185), .Y(n28176) );
  NOR2X1 U22816 ( .A(n28186), .B(n28187), .Y(n28185) );
  OAI22X1 U22817 ( .A(n25040), .B(n26094), .C(n25254), .D(n25874), .Y(n28187)
         );
  OAI21X1 U22818 ( .A(n25042), .B(n25584), .C(n28188), .Y(n28186) );
  INVX1 U22819 ( .A(n28189), .Y(n28188) );
  OAI21X1 U22820 ( .A(n25873), .B(n25334), .C(n25836), .Y(n28189) );
  NAND2X1 U22821 ( .A(reg_A[87]), .B(n25124), .Y(n25836) );
  AOI22X1 U22822 ( .A(reg_A[85]), .B(n25253), .C(reg_A[86]), .D(n25628), .Y(
        n28184) );
  AOI22X1 U22823 ( .A(reg_A[83]), .B(n25070), .C(reg_A[84]), .D(n25123), .Y(
        n28183) );
  AOI21X1 U22824 ( .A(n28190), .B(n28191), .C(n25947), .Y(n28174) );
  NOR2X1 U22825 ( .A(n25031), .B(n28192), .Y(n28190) );
  OAI21X1 U22826 ( .A(n28107), .B(n28193), .C(n28194), .Y(n28172) );
  NAND3X1 U22827 ( .A(n28195), .B(n28196), .C(n28197), .Y(result[78]) );
  NOR2X1 U22828 ( .A(n28198), .B(n28199), .Y(n28197) );
  NAND2X1 U22829 ( .A(n28200), .B(n28201), .Y(n28199) );
  NOR2X1 U22830 ( .A(n28202), .B(n28203), .Y(n28201) );
  OAI21X1 U22831 ( .A(n28204), .B(n28193), .C(n28205), .Y(n28203) );
  OAI21X1 U22832 ( .A(n28206), .B(n28207), .C(reg_A[75]), .Y(n28205) );
  OAI22X1 U22833 ( .A(n28107), .B(n28208), .C(n28209), .D(n28210), .Y(n28207)
         );
  INVX1 U22834 ( .A(n28211), .Y(n28107) );
  AOI21X1 U22835 ( .A(n26267), .B(n28157), .C(n28212), .Y(n28204) );
  OAI22X1 U22836 ( .A(n28213), .B(n28214), .C(n26286), .D(n28215), .Y(n28212)
         );
  OAI21X1 U22837 ( .A(n28216), .B(n28217), .C(n28218), .Y(n28202) );
  OAI21X1 U22838 ( .A(n28219), .B(n28220), .C(n26480), .Y(n28218) );
  OAI22X1 U22839 ( .A(n26624), .B(n28093), .C(n28221), .D(n26997), .Y(n28220)
         );
  OAI22X1 U22840 ( .A(n28222), .B(n25964), .C(n28223), .D(n25967), .Y(n28219)
         );
  INVX1 U22841 ( .A(n26114), .Y(n28223) );
  AOI21X1 U22842 ( .A(n28224), .B(n26139), .C(n28225), .Y(n28200) );
  OAI21X1 U22843 ( .A(n28226), .B(n28192), .C(n28227), .Y(n28225) );
  OAI21X1 U22844 ( .A(n28228), .B(n28229), .C(n25932), .Y(n28227) );
  OAI21X1 U22845 ( .A(n25950), .B(n28230), .C(n28231), .Y(n28229) );
  AOI22X1 U22846 ( .A(n26276), .B(n28115), .C(n26149), .D(n28232), .Y(n28231)
         );
  OAI21X1 U22847 ( .A(n28233), .B(n26168), .C(n28234), .Y(n28228) );
  AOI21X1 U22848 ( .A(n25984), .B(n28117), .C(n27537), .Y(n28234) );
  OAI21X1 U22849 ( .A(n25964), .B(n26256), .C(n28235), .Y(n28117) );
  AOI22X1 U22850 ( .A(reg_B[93]), .B(n27916), .C(reg_A[78]), .D(n26057), .Y(
        n28235) );
  INVX1 U22851 ( .A(n28118), .Y(n28233) );
  INVX1 U22852 ( .A(n28236), .Y(n28226) );
  NAND2X1 U22853 ( .A(n28237), .B(n28238), .Y(n28198) );
  NOR2X1 U22854 ( .A(n28239), .B(n28240), .Y(n28238) );
  OAI21X1 U22855 ( .A(n28241), .B(n28242), .C(n28243), .Y(n28240) );
  NAND3X1 U22856 ( .A(n26267), .B(n28244), .C(n28245), .Y(n28243) );
  NAND2X1 U22857 ( .A(n28073), .B(n25188), .Y(n28242) );
  OAI21X1 U22858 ( .A(n26151), .B(n28246), .C(n28247), .Y(n28239) );
  NAND2X1 U22859 ( .A(n28133), .B(n28248), .Y(n28246) );
  OAI21X1 U22860 ( .A(n25863), .B(n28209), .C(n28249), .Y(n28133) );
  AOI22X1 U22861 ( .A(n28250), .B(reg_B[77]), .C(n28251), .D(reg_A[78]), .Y(
        n28249) );
  MUX2X1 U22862 ( .B(n26438), .A(n26547), .S(reg_B[78]), .Y(n28250) );
  AOI21X1 U22863 ( .A(n28252), .B(n28253), .C(n28254), .Y(n28237) );
  NAND2X1 U22864 ( .A(n28255), .B(n28256), .Y(n28254) );
  OAI21X1 U22865 ( .A(n28257), .B(n28258), .C(n28211), .Y(n28256) );
  INVX1 U22866 ( .A(n28259), .Y(n28257) );
  OAI21X1 U22867 ( .A(n28260), .B(n28261), .C(n25310), .Y(n28255) );
  NAND3X1 U22868 ( .A(n28262), .B(n28263), .C(n28264), .Y(n28261) );
  NOR2X1 U22869 ( .A(n28265), .B(n28266), .Y(n28264) );
  OAI22X1 U22870 ( .A(n25035), .B(n25882), .C(n25219), .D(n26195), .Y(n28266)
         );
  OAI21X1 U22871 ( .A(n25027), .B(n25929), .C(n28267), .Y(n28265) );
  AOI22X1 U22872 ( .A(reg_A[87]), .B(n25629), .C(reg_A[86]), .D(n25124), .Y(
        n28267) );
  AOI22X1 U22873 ( .A(reg_A[93]), .B(n25235), .C(reg_A[90]), .D(n25635), .Y(
        n28263) );
  AOI22X1 U22874 ( .A(reg_A[91]), .B(n25325), .C(reg_A[78]), .D(n25125), .Y(
        n28262) );
  NAND3X1 U22875 ( .A(n28268), .B(n28269), .C(n28270), .Y(n28260) );
  NOR2X1 U22876 ( .A(n28271), .B(n28272), .Y(n28270) );
  OAI22X1 U22877 ( .A(n25040), .B(n25584), .C(n25041), .D(n26094), .Y(n28272)
         );
  OAI21X1 U22878 ( .A(n25042), .B(n25864), .C(n28273), .Y(n28271) );
  AOI22X1 U22879 ( .A(reg_A[95]), .B(n25246), .C(reg_A[94]), .D(n25247), .Y(
        n28273) );
  AOI22X1 U22880 ( .A(reg_A[84]), .B(n25253), .C(reg_A[85]), .D(n25628), .Y(
        n28269) );
  AOI22X1 U22881 ( .A(reg_A[82]), .B(n25071), .C(reg_A[83]), .D(n25123), .Y(
        n28268) );
  NOR2X1 U22882 ( .A(n28274), .B(n28275), .Y(n28196) );
  OAI21X1 U22883 ( .A(n28276), .B(n25863), .C(n28277), .Y(n28275) );
  AOI22X1 U22884 ( .A(reg_A[74]), .B(n26026), .C(reg_A[78]), .D(n28082), .Y(
        n28277) );
  NAND2X1 U22885 ( .A(n28278), .B(n28279), .Y(n28274) );
  AOI22X1 U22886 ( .A(reg_A[79]), .B(n28280), .C(reg_A[64]), .D(n28281), .Y(
        n28279) );
  AOI22X1 U22887 ( .A(reg_A[72]), .B(n26043), .C(reg_A[73]), .D(n28282), .Y(
        n28278) );
  NOR2X1 U22888 ( .A(n28283), .B(n28284), .Y(n28195) );
  OAI21X1 U22889 ( .A(n28285), .B(n27020), .C(n28286), .Y(n28284) );
  AOI22X1 U22890 ( .A(n26045), .B(n28287), .C(n28288), .D(n28289), .Y(n28286)
         );
  INVX1 U22891 ( .A(n28129), .Y(n28289) );
  MUX2X1 U22892 ( .B(n28290), .A(n28291), .S(reg_B[78]), .Y(n28129) );
  NAND2X1 U22893 ( .A(n28292), .B(n28293), .Y(n28290) );
  AOI22X1 U22894 ( .A(n28294), .B(reg_B[77]), .C(n28073), .D(reg_A[70]), .Y(
        n28293) );
  NOR2X1 U22895 ( .A(n25884), .B(n28295), .Y(n28294) );
  AOI22X1 U22896 ( .A(n28296), .B(reg_A[74]), .C(n28297), .D(reg_A[78]), .Y(
        n28292) );
  NAND3X1 U22897 ( .A(n28298), .B(n28299), .C(n28300), .Y(n28287) );
  NOR2X1 U22898 ( .A(n28301), .B(n28302), .Y(n28300) );
  OAI21X1 U22899 ( .A(n26286), .B(n28303), .C(n28304), .Y(n28302) );
  OAI21X1 U22900 ( .A(n28305), .B(n28306), .C(n25604), .Y(n28304) );
  NAND2X1 U22901 ( .A(n28307), .B(n28308), .Y(n28306) );
  AOI22X1 U22902 ( .A(reg_A[68]), .B(n25607), .C(reg_A[64]), .D(n25608), .Y(
        n28308) );
  AOI22X1 U22903 ( .A(reg_A[66]), .B(n25609), .C(reg_A[65]), .D(n25610), .Y(
        n28307) );
  NAND2X1 U22904 ( .A(n28309), .B(n28310), .Y(n28305) );
  AOI22X1 U22905 ( .A(reg_A[71]), .B(n25613), .C(reg_A[69]), .D(n25614), .Y(
        n28310) );
  AOI22X1 U22906 ( .A(reg_A[70]), .B(n25615), .C(reg_A[67]), .D(n25616), .Y(
        n28309) );
  OAI22X1 U22907 ( .A(n28311), .B(n26547), .C(n25449), .D(n26439), .Y(n28301)
         );
  AOI22X1 U22908 ( .A(reg_A[75]), .B(n25442), .C(reg_A[74]), .D(n27387), .Y(
        n28299) );
  AOI22X1 U22909 ( .A(reg_A[76]), .B(n28312), .C(reg_A[78]), .D(n25434), .Y(
        n28298) );
  INVX1 U22910 ( .A(n28313), .Y(n28285) );
  OR2X1 U22911 ( .A(n28314), .B(n28315), .Y(n28283) );
  OAI22X1 U22912 ( .A(n28135), .B(n26950), .C(n28316), .D(n26919), .Y(n28315)
         );
  AND2X1 U22913 ( .A(n28317), .B(n28318), .Y(n28135) );
  AOI22X1 U22914 ( .A(n26159), .B(n28319), .C(n25838), .D(n27505), .Y(n28318)
         );
  OAI22X1 U22915 ( .A(n26131), .B(n26256), .C(n25894), .D(n25865), .Y(n27505)
         );
  INVX1 U22916 ( .A(n26112), .Y(n26159) );
  NAND2X1 U22917 ( .A(reg_B[93]), .B(reg_B[94]), .Y(n26112) );
  AOI22X1 U22918 ( .A(n26160), .B(n27691), .C(n26059), .D(n27916), .Y(n28317)
         );
  NAND2X1 U22919 ( .A(reg_B[94]), .B(n26197), .Y(n26338) );
  OAI21X1 U22920 ( .A(n28320), .B(n26286), .C(n28321), .Y(n28314) );
  OAI21X1 U22921 ( .A(n28322), .B(n28323), .C(n25119), .Y(n28321) );
  NAND3X1 U22922 ( .A(n28324), .B(n28325), .C(n28326), .Y(n28323) );
  AOI21X1 U22923 ( .A(reg_A[78]), .B(n25125), .C(n28327), .Y(n28326) );
  OAI22X1 U22924 ( .A(n25039), .B(n25855), .C(n25231), .D(n25884), .Y(n28327)
         );
  AOI22X1 U22925 ( .A(reg_A[69]), .B(n25629), .C(reg_A[70]), .D(n25124), .Y(
        n28325) );
  AOI22X1 U22926 ( .A(reg_A[67]), .B(n25222), .C(reg_A[68]), .D(n25637), .Y(
        n28324) );
  NAND3X1 U22927 ( .A(n28328), .B(n28329), .C(n28330), .Y(n28322) );
  AOI21X1 U22928 ( .A(reg_A[73]), .B(n25123), .C(n28331), .Y(n28330) );
  OAI22X1 U22929 ( .A(n26431), .B(n26438), .C(n25129), .D(n26101), .Y(n28331)
         );
  AOI22X1 U22930 ( .A(reg_A[77]), .B(n25135), .C(reg_A[75]), .D(n25136), .Y(
        n28329) );
  AOI22X1 U22931 ( .A(reg_A[76]), .B(n25252), .C(reg_A[72]), .D(n25253), .Y(
        n28328) );
  INVX1 U22932 ( .A(n28332), .Y(n28320) );
  NAND3X1 U22933 ( .A(n28333), .B(n28334), .C(n28335), .Y(result[77]) );
  NOR2X1 U22934 ( .A(n28336), .B(n28337), .Y(n28335) );
  NAND2X1 U22935 ( .A(n28338), .B(n28339), .Y(n28337) );
  AOI21X1 U22936 ( .A(n28083), .B(n28340), .C(n28341), .Y(n28339) );
  OAI22X1 U22937 ( .A(n25994), .B(n28342), .C(n25148), .D(n25865), .Y(n28341)
         );
  AOI21X1 U22938 ( .A(n28343), .B(reg_A[77]), .C(n28344), .Y(n28338) );
  OAI21X1 U22939 ( .A(n28345), .B(n25835), .C(n28346), .Y(n28344) );
  OAI21X1 U22940 ( .A(n28347), .B(n28348), .C(n26045), .Y(n28346) );
  NAND3X1 U22941 ( .A(n28349), .B(n28350), .C(n28351), .Y(n28348) );
  AOI21X1 U22942 ( .A(reg_A[77]), .B(n25434), .C(n28352), .Y(n28351) );
  OAI22X1 U22943 ( .A(n28353), .B(n26103), .C(n25205), .D(n26439), .Y(n28352)
         );
  AOI22X1 U22944 ( .A(n25097), .B(n28354), .C(reg_A[72]), .D(n28355), .Y(
        n28350) );
  AOI22X1 U22945 ( .A(reg_A[76]), .B(n25441), .C(reg_A[74]), .D(n27241), .Y(
        n28349) );
  NAND3X1 U22946 ( .A(n28356), .B(n28357), .C(n28358), .Y(n28347) );
  NOR2X1 U22947 ( .A(n28359), .B(n28360), .Y(n28358) );
  OAI22X1 U22948 ( .A(n28361), .B(n25853), .C(n28311), .D(n26101), .Y(n28360)
         );
  OAI22X1 U22949 ( .A(n28362), .B(n25851), .C(n28363), .D(n25884), .Y(n28359)
         );
  AOI22X1 U22950 ( .A(reg_A[65]), .B(n28364), .C(reg_A[68]), .D(n25500), .Y(
        n28357) );
  AOI22X1 U22951 ( .A(reg_A[69]), .B(n25501), .C(reg_A[70]), .D(n25502), .Y(
        n28356) );
  INVX1 U22952 ( .A(n28354), .Y(n28345) );
  NAND3X1 U22953 ( .A(n28365), .B(n28366), .C(n28367), .Y(n28354) );
  NOR2X1 U22954 ( .A(n28368), .B(n28369), .Y(n28367) );
  OAI21X1 U22955 ( .A(n25043), .B(n26286), .C(n28370), .Y(n28369) );
  AOI22X1 U22956 ( .A(reg_A[67]), .B(n25637), .C(reg_A[65]), .D(n25635), .Y(
        n28370) );
  OAI21X1 U22957 ( .A(n25027), .B(n25884), .C(n28371), .Y(n28368) );
  AOI22X1 U22958 ( .A(reg_A[68]), .B(n25629), .C(reg_A[69]), .D(n25124), .Y(
        n28371) );
  NOR2X1 U22959 ( .A(n28372), .B(n28373), .Y(n28366) );
  OAI22X1 U22960 ( .A(n25033), .B(n26101), .C(n25040), .D(n26103), .Y(n28373)
         );
  OAI22X1 U22961 ( .A(n25041), .B(n26438), .C(n25784), .D(n25863), .Y(n28372)
         );
  AOI21X1 U22962 ( .A(reg_A[72]), .B(n25123), .C(n28374), .Y(n28365) );
  OAI22X1 U22963 ( .A(n26431), .B(n26439), .C(n25030), .D(n26256), .Y(n28374)
         );
  NAND2X1 U22964 ( .A(n28375), .B(n28376), .Y(n28336) );
  AOI21X1 U22965 ( .A(n28069), .B(n28377), .C(n28378), .Y(n28376) );
  OAI21X1 U22966 ( .A(n26438), .B(n28379), .C(n28380), .Y(n28378) );
  OAI21X1 U22967 ( .A(n28381), .B(n28382), .C(n25932), .Y(n28380) );
  OAI21X1 U22968 ( .A(n28383), .B(n26169), .C(n28384), .Y(n28382) );
  MUX2X1 U22969 ( .B(n28114), .A(n28118), .S(n25984), .Y(n28384) );
  OAI21X1 U22970 ( .A(n25856), .B(n25964), .C(n28385), .Y(n28118) );
  AOI22X1 U22971 ( .A(reg_B[93]), .B(n27882), .C(n26057), .D(reg_A[77]), .Y(
        n28385) );
  OAI21X1 U22972 ( .A(n28386), .B(n25914), .C(n28387), .Y(n28381) );
  AOI21X1 U22973 ( .A(n26148), .B(n28115), .C(n27537), .Y(n28387) );
  INVX1 U22974 ( .A(n28232), .Y(n28386) );
  OAI22X1 U22975 ( .A(n25031), .B(n28388), .C(n28389), .D(n28390), .Y(n28069)
         );
  OAI21X1 U22976 ( .A(n28391), .B(n28192), .C(n25188), .Y(n28390) );
  OAI22X1 U22977 ( .A(n28392), .B(n28393), .C(n28394), .D(n28395), .Y(n28389)
         );
  MUX2X1 U22978 ( .B(n26286), .A(n25863), .S(reg_B[79]), .Y(n28395) );
  MUX2X1 U22979 ( .B(n28158), .A(n28396), .S(reg_B[79]), .Y(n28388) );
  MUX2X1 U22980 ( .B(n25863), .A(n26547), .S(reg_B[77]), .Y(n28396) );
  INVX1 U22981 ( .A(n28214), .Y(n28158) );
  AOI21X1 U22982 ( .A(reg_A[79]), .B(n25153), .C(n28397), .Y(n28375) );
  OAI22X1 U22983 ( .A(n26854), .B(n28123), .C(n28398), .D(n28208), .Y(n28397)
         );
  OAI21X1 U22984 ( .A(n28399), .B(n26452), .C(n28400), .Y(n28123) );
  AOI22X1 U22985 ( .A(n26293), .B(n26216), .C(n26295), .D(n26367), .Y(n28400)
         );
  INVX1 U22986 ( .A(n27682), .Y(n26367) );
  MUX2X1 U22987 ( .B(n25863), .A(n26107), .S(reg_B[1]), .Y(n27682) );
  INVX1 U22988 ( .A(n27927), .Y(n26216) );
  MUX2X1 U22989 ( .B(n26286), .A(n25856), .S(reg_B[1]), .Y(n27927) );
  INVX1 U22990 ( .A(n28401), .Y(n28399) );
  NOR2X1 U22991 ( .A(n28402), .B(n28403), .Y(n28334) );
  INVX1 U22992 ( .A(n28404), .Y(n28403) );
  AOI21X1 U22993 ( .A(n28405), .B(n28132), .C(n28406), .Y(n28404) );
  OAI22X1 U22994 ( .A(n28407), .B(n28408), .C(n28121), .D(n26278), .Y(n28406)
         );
  NAND2X1 U22995 ( .A(n28409), .B(n28410), .Y(n28121) );
  AOI22X1 U22996 ( .A(n26292), .B(n26439), .C(n26293), .D(n26286), .Y(n28410)
         );
  AOI22X1 U22997 ( .A(n26294), .B(n26547), .C(n26295), .D(n25863), .Y(n28409)
         );
  NAND3X1 U22998 ( .A(n28411), .B(n28247), .C(n28412), .Y(n28402) );
  NAND2X1 U22999 ( .A(reg_A[75]), .B(n28413), .Y(n28412) );
  OAI21X1 U23000 ( .A(n28144), .B(n28414), .C(n28415), .Y(n28413) );
  NAND3X1 U23001 ( .A(reg_B[77]), .B(reg_B[78]), .C(n28416), .Y(n28247) );
  OAI21X1 U23002 ( .A(n28417), .B(n28418), .C(n25310), .Y(n28411) );
  NAND3X1 U23003 ( .A(n28419), .B(n28420), .C(n28421), .Y(n28418) );
  NOR2X1 U23004 ( .A(n28422), .B(n28423), .Y(n28421) );
  OAI22X1 U23005 ( .A(n25035), .B(n25973), .C(n25219), .D(n25965), .Y(n28423)
         );
  OAI21X1 U23006 ( .A(n25027), .B(n26195), .C(n28424), .Y(n28422) );
  AOI22X1 U23007 ( .A(reg_A[86]), .B(n25629), .C(reg_A[85]), .D(n25124), .Y(
        n28424) );
  AOI22X1 U23008 ( .A(reg_A[92]), .B(n25235), .C(reg_A[89]), .D(n25635), .Y(
        n28420) );
  AOI22X1 U23009 ( .A(reg_A[90]), .B(n25325), .C(reg_A[77]), .D(n25125), .Y(
        n28419) );
  NAND3X1 U23010 ( .A(n28425), .B(n28426), .C(n28427), .Y(n28417) );
  NOR2X1 U23011 ( .A(n28428), .B(n28429), .Y(n28427) );
  OAI22X1 U23012 ( .A(n25041), .B(n25584), .C(n25042), .D(n25865), .Y(n28429)
         );
  OAI21X1 U23013 ( .A(n25051), .B(n25873), .C(n28430), .Y(n28428) );
  AOI22X1 U23014 ( .A(reg_A[94]), .B(n25246), .C(reg_A[93]), .D(n25247), .Y(
        n28430) );
  AOI21X1 U23015 ( .A(reg_A[84]), .B(n25628), .C(n28431), .Y(n28426) );
  OAI22X1 U23016 ( .A(n25033), .B(n25875), .C(n25040), .D(n25864), .Y(n28431)
         );
  AOI22X1 U23017 ( .A(reg_A[81]), .B(n25070), .C(reg_A[82]), .D(n25123), .Y(
        n28425) );
  NOR2X1 U23018 ( .A(n28432), .B(n28433), .Y(n28333) );
  OAI21X1 U23019 ( .A(n26547), .B(n28434), .C(n28435), .Y(n28433) );
  AOI22X1 U23020 ( .A(n26267), .B(n28436), .C(n25170), .D(n28437), .Y(n28435)
         );
  OAI21X1 U23021 ( .A(n28438), .B(n27053), .C(n28439), .Y(n28437) );
  AOI22X1 U23022 ( .A(n28440), .B(n28441), .C(n27787), .D(n28313), .Y(n28439)
         );
  OAI21X1 U23023 ( .A(n28442), .B(n25950), .C(n28443), .Y(n28313) );
  AOI22X1 U23024 ( .A(n25838), .B(n27550), .C(n26059), .D(n27882), .Y(n28443)
         );
  OAI22X1 U23025 ( .A(n25856), .B(n26131), .C(n25894), .D(n26286), .Y(n27550)
         );
  OAI22X1 U23026 ( .A(n26103), .B(n28209), .C(reg_B[78]), .D(n28214), .Y(
        n28441) );
  MUX2X1 U23027 ( .B(reg_A[77]), .A(reg_A[73]), .S(reg_B[77]), .Y(n28214) );
  OAI21X1 U23028 ( .A(n28444), .B(n28144), .C(n28445), .Y(n28436) );
  AOI22X1 U23029 ( .A(n28446), .B(n28157), .C(n28191), .D(n28291), .Y(n28445)
         );
  INVX1 U23030 ( .A(n28447), .Y(n28291) );
  NAND2X1 U23031 ( .A(n28448), .B(n28449), .Y(n28157) );
  AOI22X1 U23032 ( .A(n28450), .B(reg_B[77]), .C(n28073), .D(reg_A[69]), .Y(
        n28449) );
  NOR2X1 U23033 ( .A(n25855), .B(n28295), .Y(n28450) );
  AOI22X1 U23034 ( .A(n28296), .B(reg_A[73]), .C(n28297), .D(reg_A[77]), .Y(
        n28448) );
  OAI21X1 U23035 ( .A(n28451), .B(n26996), .C(n28452), .Y(n28432) );
  AOI22X1 U23036 ( .A(n28453), .B(reg_A[64]), .C(n28454), .D(n28455), .Y(
        n28452) );
  NOR2X1 U23037 ( .A(n28456), .B(n28457), .Y(n28451) );
  OAI22X1 U23038 ( .A(n26807), .B(n28093), .C(n28458), .D(n26997), .Y(n28457)
         );
  OAI22X1 U23039 ( .A(n28459), .B(n25964), .C(n26182), .D(n25967), .Y(n28456)
         );
  INVX1 U23040 ( .A(n28460), .Y(n26182) );
  INVX1 U23041 ( .A(n28461), .Y(n28459) );
  NAND2X1 U23042 ( .A(n28462), .B(n28463), .Y(result[76]) );
  NOR2X1 U23043 ( .A(n28464), .B(n28465), .Y(n28463) );
  NAND3X1 U23044 ( .A(n28466), .B(n28467), .C(n28468), .Y(n28465) );
  NOR2X1 U23045 ( .A(n28469), .B(n28470), .Y(n28468) );
  NAND2X1 U23046 ( .A(n28471), .B(n28472), .Y(n28470) );
  OAI21X1 U23047 ( .A(n28473), .B(n28474), .C(n28211), .Y(n28472) );
  NAND2X1 U23048 ( .A(n28414), .B(n28215), .Y(n28211) );
  OAI22X1 U23049 ( .A(n25863), .B(n28088), .C(n26439), .D(n28208), .Y(n28474)
         );
  OAI21X1 U23050 ( .A(n26438), .B(n28144), .C(n28475), .Y(n28473) );
  OAI21X1 U23051 ( .A(n28476), .B(n28477), .C(n26267), .Y(n28471) );
  OAI22X1 U23052 ( .A(n28478), .B(n28208), .C(n28479), .D(n28144), .Y(n28477)
         );
  INVX1 U23053 ( .A(n28480), .Y(n28479) );
  OAI22X1 U23054 ( .A(n28444), .B(n28193), .C(n28447), .D(n28088), .Y(n28476)
         );
  NOR2X1 U23055 ( .A(n28481), .B(n28482), .Y(n28447) );
  OAI22X1 U23056 ( .A(n26547), .B(n28483), .C(n25863), .D(n28394), .Y(n28482)
         );
  OAI21X1 U23057 ( .A(n26107), .B(n28393), .C(n28484), .Y(n28481) );
  INVX1 U23058 ( .A(n28244), .Y(n28444) );
  OAI21X1 U23059 ( .A(n28485), .B(n27438), .C(n28486), .Y(n28469) );
  OAI21X1 U23060 ( .A(n28487), .B(n28488), .C(n25188), .Y(n28486) );
  OAI21X1 U23061 ( .A(n28393), .B(n28489), .C(n28484), .Y(n28488) );
  NOR2X1 U23062 ( .A(n28483), .B(n28490), .Y(n28487) );
  INVX1 U23063 ( .A(n28491), .Y(n28485) );
  OAI21X1 U23064 ( .A(n25914), .B(n28383), .C(n28492), .Y(n28491) );
  AOI22X1 U23065 ( .A(n28232), .B(n26148), .C(n28115), .D(n25984), .Y(n28492)
         );
  OAI21X1 U23066 ( .A(n26547), .B(n26997), .C(n28493), .Y(n28115) );
  AOI22X1 U23067 ( .A(reg_A[76]), .B(n26057), .C(reg_A[68]), .D(n26307), .Y(
        n28493) );
  AOI22X1 U23068 ( .A(reg_A[64]), .B(n28494), .C(reg_A[73]), .D(n28495), .Y(
        n28467) );
  AOI22X1 U23069 ( .A(reg_A[74]), .B(n28496), .C(n26149), .D(n28497), .Y(
        n28466) );
  NAND3X1 U23070 ( .A(n28498), .B(n28499), .C(n28500), .Y(n28464) );
  NOR2X1 U23071 ( .A(n28501), .B(n28502), .Y(n28500) );
  OAI21X1 U23072 ( .A(n28503), .B(n28217), .C(n28504), .Y(n28502) );
  OAI21X1 U23073 ( .A(n28505), .B(n28506), .C(n26480), .Y(n28504) );
  OAI22X1 U23074 ( .A(n28507), .B(n26997), .C(n28508), .D(n25964), .Y(n28506)
         );
  INVX1 U23075 ( .A(n28509), .Y(n28508) );
  OAI22X1 U23076 ( .A(n28510), .B(n28093), .C(n26329), .D(n25967), .Y(n28505)
         );
  INVX1 U23077 ( .A(n26992), .Y(n26329) );
  OAI22X1 U23078 ( .A(n28511), .B(n28210), .C(n25884), .D(n28512), .Y(n28501)
         );
  AOI21X1 U23079 ( .A(n28513), .B(n28405), .C(n28514), .Y(n28499) );
  OAI21X1 U23080 ( .A(n28515), .B(n28516), .C(n28517), .Y(n28514) );
  OAI21X1 U23081 ( .A(n28518), .B(n28519), .C(n25310), .Y(n28517) );
  NAND3X1 U23082 ( .A(n28520), .B(n28521), .C(n28522), .Y(n28519) );
  NOR2X1 U23083 ( .A(n28523), .B(n28524), .Y(n28522) );
  OAI22X1 U23084 ( .A(n25043), .B(n25863), .C(n25039), .D(n25929), .Y(n28524)
         );
  OAI21X1 U23085 ( .A(n25064), .B(n26195), .C(n28525), .Y(n28523) );
  AOI22X1 U23086 ( .A(reg_A[90]), .B(n25234), .C(reg_A[91]), .D(n25235), .Y(
        n28525) );
  AOI21X1 U23087 ( .A(reg_A[84]), .B(n25124), .C(n28526), .Y(n28521) );
  OAI22X1 U23088 ( .A(n25037), .B(n26215), .C(n25028), .D(n26094), .Y(n28526)
         );
  AOI22X1 U23089 ( .A(reg_A[87]), .B(n25222), .C(reg_A[86]), .D(n25637), .Y(
        n28520) );
  NAND3X1 U23090 ( .A(n28527), .B(n28528), .C(n28529), .Y(n28518) );
  NOR2X1 U23091 ( .A(n28530), .B(n28531), .Y(n28529) );
  OAI22X1 U23092 ( .A(n25042), .B(n26286), .C(n25331), .D(n25883), .Y(n28531)
         );
  OAI21X1 U23093 ( .A(n25038), .B(n25873), .C(n28532), .Y(n28530) );
  AOI22X1 U23094 ( .A(reg_A[93]), .B(n25246), .C(reg_A[92]), .D(n25247), .Y(
        n28532) );
  AOI21X1 U23095 ( .A(reg_A[82]), .B(n25253), .C(n28533), .Y(n28528) );
  OAI22X1 U23096 ( .A(n25040), .B(n25865), .C(n25041), .D(n25864), .Y(n28533)
         );
  AOI22X1 U23097 ( .A(reg_A[83]), .B(n25628), .C(reg_A[80]), .D(n25067), .Y(
        n28527) );
  AND2X1 U23098 ( .A(n28534), .B(n28535), .Y(n28515) );
  NOR2X1 U23099 ( .A(n28536), .B(n28537), .Y(n28535) );
  OAI21X1 U23100 ( .A(n25043), .B(n25863), .C(n28538), .Y(n28537) );
  AOI22X1 U23101 ( .A(reg_A[75]), .B(n25135), .C(reg_A[74]), .D(n25252), .Y(
        n28538) );
  OAI21X1 U23102 ( .A(n25028), .B(n26101), .C(n28539), .Y(n28536) );
  AOI22X1 U23103 ( .A(reg_A[73]), .B(n25136), .C(reg_A[72]), .D(n25066), .Y(
        n28539) );
  NOR2X1 U23104 ( .A(n28540), .B(n28541), .Y(n28534) );
  OAI21X1 U23105 ( .A(n25034), .B(n26107), .C(n28542), .Y(n28541) );
  AOI22X1 U23106 ( .A(reg_A[70]), .B(n25253), .C(reg_A[69]), .D(n25628), .Y(
        n28542) );
  OAI21X1 U23107 ( .A(n25036), .B(n25884), .C(n28543), .Y(n28540) );
  AOI22X1 U23108 ( .A(reg_A[67]), .B(n25629), .C(reg_A[65]), .D(n25222), .Y(
        n28543) );
  OAI21X1 U23109 ( .A(n26438), .B(n28209), .C(n28544), .Y(n28405) );
  AOI22X1 U23110 ( .A(n28545), .B(reg_B[77]), .C(n28251), .D(reg_A[76]), .Y(
        n28544) );
  NOR2X1 U23111 ( .A(reg_B[78]), .B(n26547), .Y(n28545) );
  INVX1 U23112 ( .A(n28546), .Y(n28209) );
  AOI22X1 U23113 ( .A(n28547), .B(n28548), .C(n28549), .D(reg_A[65]), .Y(
        n28498) );
  NOR2X1 U23114 ( .A(n28550), .B(n28551), .Y(n28462) );
  NAND3X1 U23115 ( .A(n28552), .B(n28553), .C(n28554), .Y(n28551) );
  NOR2X1 U23116 ( .A(n28555), .B(n28556), .Y(n28554) );
  OAI21X1 U23117 ( .A(n28438), .B(n26950), .C(n28557), .Y(n28556) );
  INVX1 U23118 ( .A(n28558), .Y(n28438) );
  OAI21X1 U23119 ( .A(n28559), .B(n25950), .C(n28560), .Y(n28558) );
  AOI22X1 U23120 ( .A(n25838), .B(n27691), .C(n26059), .D(n28319), .Y(n28560)
         );
  INVX1 U23121 ( .A(n25898), .Y(n26059) );
  NAND2X1 U23122 ( .A(reg_B[93]), .B(n25950), .Y(n25898) );
  OAI22X1 U23123 ( .A(n26131), .B(n26107), .C(n25894), .D(n25863), .Y(n27691)
         );
  NAND2X1 U23124 ( .A(n26197), .B(n25950), .Y(n26337) );
  OAI22X1 U23125 ( .A(n28561), .B(n26919), .C(n25856), .D(n28562), .Y(n28555)
         );
  AOI22X1 U23126 ( .A(reg_A[77]), .B(n28280), .C(reg_A[75]), .D(n26358), .Y(
        n28553) );
  AOI22X1 U23127 ( .A(reg_A[76]), .B(n28563), .C(reg_A[72]), .D(n26348), .Y(
        n28552) );
  NAND3X1 U23128 ( .A(n28564), .B(n28565), .C(n28566), .Y(n28550) );
  NOR2X1 U23129 ( .A(n28567), .B(n28568), .Y(n28566) );
  OAI22X1 U23130 ( .A(n28569), .B(n25865), .C(n28570), .D(n25864), .Y(n28568)
         );
  OAI22X1 U23131 ( .A(n28571), .B(n26101), .C(n25178), .D(n26107), .Y(n28567)
         );
  AOI22X1 U23132 ( .A(n28572), .B(reg_A[67]), .C(n28573), .D(n26139), .Y(
        n28565) );
  AOI22X1 U23133 ( .A(n28574), .B(n28575), .C(n28576), .D(reg_A[70]), .Y(
        n28564) );
  NAND2X1 U23134 ( .A(n28577), .B(n28578), .Y(result[75]) );
  NOR2X1 U23135 ( .A(n28579), .B(n28580), .Y(n28578) );
  NAND3X1 U23136 ( .A(n28581), .B(n28582), .C(n28583), .Y(n28580) );
  NOR2X1 U23137 ( .A(n28584), .B(n28585), .Y(n28583) );
  OAI22X1 U23138 ( .A(n28586), .B(n26439), .C(n28587), .D(n25914), .Y(n28585)
         );
  OAI22X1 U23139 ( .A(n28588), .B(n26169), .C(n28398), .D(n28193), .Y(n28584)
         );
  AOI22X1 U23140 ( .A(n28480), .B(n26267), .C(reg_A[74]), .D(n28589), .Y(
        n28398) );
  AOI21X1 U23141 ( .A(reg_A[64]), .B(n28590), .C(n28591), .Y(n28582) );
  OAI21X1 U23142 ( .A(n25864), .B(n28592), .C(n28593), .Y(n28591) );
  OAI21X1 U23143 ( .A(n28594), .B(n28595), .C(n26480), .Y(n28593) );
  OAI22X1 U23144 ( .A(n28596), .B(n26997), .C(n28094), .D(n28093), .Y(n28595)
         );
  INVX1 U23145 ( .A(n28597), .Y(n28094) );
  OAI22X1 U23146 ( .A(n28095), .B(n25964), .C(n27027), .D(n26479), .Y(n28594)
         );
  AOI22X1 U23147 ( .A(n25932), .B(n28598), .C(n26267), .D(n28599), .Y(n28581)
         );
  OAI21X1 U23148 ( .A(n28600), .B(n28208), .C(n28601), .Y(n28599) );
  AOI22X1 U23149 ( .A(n28446), .B(n28244), .C(n28602), .D(n28603), .Y(n28601)
         );
  OAI21X1 U23150 ( .A(n26103), .B(n28394), .C(n28604), .Y(n28244) );
  AOI22X1 U23151 ( .A(n28073), .B(reg_A[67]), .C(n28296), .D(reg_A[71]), .Y(
        n28604) );
  OAI21X1 U23152 ( .A(n28605), .B(n26169), .C(n28606), .Y(n28598) );
  AOI22X1 U23153 ( .A(n25984), .B(n28232), .C(n26148), .D(n28607), .Y(n28606)
         );
  OAI21X1 U23154 ( .A(n25964), .B(n25851), .C(n28608), .Y(n28232) );
  AOI21X1 U23155 ( .A(reg_A[75]), .B(n26057), .C(n28609), .Y(n28608) );
  NAND3X1 U23156 ( .A(n28610), .B(n28611), .C(n28612), .Y(n28579) );
  NOR2X1 U23157 ( .A(n28613), .B(n28614), .Y(n28612) );
  OAI21X1 U23158 ( .A(n28407), .B(n28615), .C(n28616), .Y(n28614) );
  OAI21X1 U23159 ( .A(n28617), .B(n28618), .C(n25310), .Y(n28616) );
  NAND3X1 U23160 ( .A(n28619), .B(n28620), .C(n28621), .Y(n28618) );
  NOR2X1 U23161 ( .A(n28622), .B(n28623), .Y(n28621) );
  OAI22X1 U23162 ( .A(n25043), .B(n26103), .C(n25039), .D(n26195), .Y(n28623)
         );
  OAI21X1 U23163 ( .A(n25064), .B(n25965), .C(n28624), .Y(n28622) );
  AOI22X1 U23164 ( .A(reg_A[89]), .B(n25234), .C(reg_A[90]), .D(n25235), .Y(
        n28624) );
  AOI21X1 U23165 ( .A(reg_A[83]), .B(n25124), .C(n28625), .Y(n28620) );
  OAI22X1 U23166 ( .A(n25037), .B(n26230), .C(n25028), .D(n25584), .Y(n28625)
         );
  AOI22X1 U23167 ( .A(reg_A[86]), .B(n25222), .C(reg_A[85]), .D(n25637), .Y(
        n28619) );
  NAND3X1 U23168 ( .A(n28626), .B(n28627), .C(n28628), .Y(n28617) );
  NOR2X1 U23169 ( .A(n28629), .B(n28630), .Y(n28628) );
  OAI21X1 U23170 ( .A(n25042), .B(n25863), .C(n28631), .Y(n28630) );
  AOI22X1 U23171 ( .A(reg_A[93]), .B(n25241), .C(reg_A[95]), .D(n25339), .Y(
        n28631) );
  OAI21X1 U23172 ( .A(n25038), .B(n25883), .C(n28632), .Y(n28629) );
  AOI22X1 U23173 ( .A(reg_A[92]), .B(n25246), .C(reg_A[91]), .D(n25247), .Y(
        n28632) );
  AOI21X1 U23174 ( .A(reg_A[81]), .B(n25253), .C(n28633), .Y(n28627) );
  OAI22X1 U23175 ( .A(n25040), .B(n26286), .C(n25254), .D(n25865), .Y(n28633)
         );
  AOI22X1 U23176 ( .A(reg_A[82]), .B(n25628), .C(reg_A[79]), .D(n25067), .Y(
        n28626) );
  OAI21X1 U23177 ( .A(n28511), .B(n28634), .C(n28635), .Y(n28613) );
  AOI22X1 U23178 ( .A(n28636), .B(n28637), .C(n28638), .D(n25382), .Y(n28635)
         );
  NOR2X1 U23179 ( .A(n28102), .B(n28639), .Y(n28638) );
  INVX1 U23180 ( .A(n28408), .Y(n28637) );
  OAI21X1 U23181 ( .A(n28072), .B(n28483), .C(n28640), .Y(n28408) );
  AOI21X1 U23182 ( .A(n28641), .B(n28192), .C(n28642), .Y(n28640) );
  INVX1 U23183 ( .A(n28071), .Y(n28641) );
  MUX2X1 U23184 ( .B(n28643), .A(n28644), .S(reg_B[79]), .Y(n28071) );
  INVX1 U23185 ( .A(n28645), .Y(n28644) );
  MUX2X1 U23186 ( .B(reg_A[75]), .A(reg_A[67]), .S(reg_B[76]), .Y(n28643) );
  NOR2X1 U23187 ( .A(reg_B[78]), .B(n25032), .Y(n28636) );
  AOI21X1 U23188 ( .A(n26504), .B(n28248), .C(n28513), .Y(n28634) );
  INVX1 U23189 ( .A(n28646), .Y(n28513) );
  AOI22X1 U23190 ( .A(reg_A[73]), .B(n28546), .C(reg_A[75]), .D(n28251), .Y(
        n28511) );
  AOI22X1 U23191 ( .A(n28647), .B(n28548), .C(n28547), .D(n28648), .Y(n28611)
         );
  INVX1 U23192 ( .A(n28559), .Y(n28648) );
  INVX1 U23193 ( .A(n28442), .Y(n28548) );
  AOI21X1 U23194 ( .A(n27761), .B(n26197), .C(n28609), .Y(n28442) );
  OAI22X1 U23195 ( .A(n26131), .B(n25851), .C(n25894), .D(n26103), .Y(n27761)
         );
  AOI22X1 U23196 ( .A(n28649), .B(reg_A[65]), .C(n28132), .D(n28650), .Y(
        n28610) );
  INVX1 U23197 ( .A(n28651), .Y(n28650) );
  INVX1 U23198 ( .A(n28210), .Y(n28132) );
  NAND2X1 U23199 ( .A(reg_B[79]), .B(n26186), .Y(n28210) );
  NOR2X1 U23200 ( .A(n28652), .B(n28653), .Y(n28577) );
  NAND3X1 U23201 ( .A(n28654), .B(n28655), .C(n28656), .Y(n28653) );
  NOR2X1 U23202 ( .A(n28657), .B(n28658), .Y(n28656) );
  OAI21X1 U23203 ( .A(n28659), .B(n28208), .C(n28557), .Y(n28658) );
  OAI22X1 U23204 ( .A(n28660), .B(n26919), .C(n26107), .D(n28562), .Y(n28657)
         );
  AOI21X1 U23205 ( .A(reg_A[75]), .B(n28661), .C(n28662), .Y(n28655) );
  OAI22X1 U23206 ( .A(n25994), .B(n28663), .C(n28664), .D(n26547), .Y(n28662)
         );
  AOI22X1 U23207 ( .A(reg_A[74]), .B(n26626), .C(n28665), .D(n25119), .Y(
        n28654) );
  NAND3X1 U23208 ( .A(n28666), .B(n28667), .C(n28668), .Y(n28665) );
  NOR2X1 U23209 ( .A(n28669), .B(n28670), .Y(n28668) );
  OAI21X1 U23210 ( .A(n25056), .B(n26101), .C(n28671), .Y(n28670) );
  AOI22X1 U23211 ( .A(reg_A[69]), .B(n25253), .C(reg_A[68]), .D(n25628), .Y(
        n28671) );
  OAI21X1 U23212 ( .A(n25040), .B(n26439), .C(n28672), .Y(n28669) );
  AOI22X1 U23213 ( .A(reg_A[74]), .B(n25135), .C(reg_A[72]), .D(n25136), .Y(
        n28672) );
  AOI21X1 U23214 ( .A(reg_A[67]), .B(n25124), .C(n28673), .Y(n28667) );
  OAI22X1 U23215 ( .A(n25037), .B(n25884), .C(n25028), .D(n26256), .Y(n28673)
         );
  AOI22X1 U23216 ( .A(reg_A[65]), .B(n25637), .C(reg_A[75]), .D(n25125), .Y(
        n28666) );
  NAND3X1 U23217 ( .A(n28674), .B(n28675), .C(n28676), .Y(n28652) );
  NOR2X1 U23218 ( .A(n28677), .B(n28678), .Y(n28676) );
  OAI22X1 U23219 ( .A(n28571), .B(n26256), .C(n25178), .D(n25851), .Y(n28678)
         );
  OAI21X1 U23220 ( .A(n28679), .B(n26101), .C(n28680), .Y(n28677) );
  AOI22X1 U23221 ( .A(n28572), .B(reg_A[66]), .C(n28576), .D(reg_A[69]), .Y(
        n28680) );
  AOI22X1 U23222 ( .A(n28681), .B(n25150), .C(reg_A[78]), .D(n25152), .Y(
        n28675) );
  INVX1 U23223 ( .A(n28342), .Y(n28681) );
  OAI21X1 U23224 ( .A(reg_B[2]), .B(n28137), .C(n28682), .Y(n28342) );
  AOI22X1 U23225 ( .A(n26455), .B(n25853), .C(n26456), .D(n28683), .Y(n28682)
         );
  INVX1 U23226 ( .A(n28684), .Y(n28137) );
  OAI21X1 U23227 ( .A(reg_B[4]), .B(n27823), .C(n28685), .Y(n28684) );
  AOI22X1 U23228 ( .A(n26462), .B(n26438), .C(n26463), .D(n25884), .Y(n28685)
         );
  MUX2X1 U23229 ( .B(n26103), .A(n25851), .S(reg_B[1]), .Y(n27823) );
  AOI22X1 U23230 ( .A(reg_A[77]), .B(n25153), .C(reg_A[76]), .D(n28280), .Y(
        n28674) );
  NAND3X1 U23231 ( .A(n28686), .B(n28687), .C(n28688), .Y(result[74]) );
  NOR2X1 U23232 ( .A(n28689), .B(n28690), .Y(n28688) );
  NAND3X1 U23233 ( .A(n28691), .B(n28692), .C(n28693), .Y(n28690) );
  NOR2X1 U23234 ( .A(n28694), .B(n28695), .Y(n28693) );
  OAI21X1 U23235 ( .A(n28377), .B(n28659), .C(n28557), .Y(n28695) );
  OAI22X1 U23236 ( .A(n28696), .B(n26919), .C(n25851), .D(n28562), .Y(n28694)
         );
  INVX1 U23237 ( .A(n28697), .Y(n28692) );
  OAI21X1 U23238 ( .A(n26438), .B(n28698), .C(n28699), .Y(n28697) );
  AOI22X1 U23239 ( .A(n28700), .B(reg_A[64]), .C(n28280), .D(reg_A[75]), .Y(
        n28699) );
  AOI22X1 U23240 ( .A(reg_A[73]), .B(n26626), .C(n28701), .D(n25119), .Y(
        n28691) );
  NAND3X1 U23241 ( .A(n28702), .B(n28703), .C(n28704), .Y(n28701) );
  NOR2X1 U23242 ( .A(n28705), .B(n28706), .Y(n28704) );
  OAI22X1 U23243 ( .A(n25043), .B(n26438), .C(n25467), .D(n25884), .Y(n28706)
         );
  OAI21X1 U23244 ( .A(n25037), .B(n25855), .C(n28707), .Y(n28705) );
  AOI22X1 U23245 ( .A(reg_A[70]), .B(n25070), .C(reg_A[69]), .D(n25123), .Y(
        n28707) );
  AOI21X1 U23246 ( .A(reg_A[72]), .B(n25252), .C(n28708), .Y(n28703) );
  OAI22X1 U23247 ( .A(n25041), .B(n26101), .C(n25042), .D(n26439), .Y(n28708)
         );
  AOI22X1 U23248 ( .A(reg_A[68]), .B(n25253), .C(reg_A[67]), .D(n25628), .Y(
        n28702) );
  NAND3X1 U23249 ( .A(n28709), .B(n28710), .C(n28711), .Y(n28689) );
  NOR2X1 U23250 ( .A(n28712), .B(n28713), .Y(n28711) );
  OAI22X1 U23251 ( .A(n28679), .B(n26256), .C(n26107), .D(n28714), .Y(n28713)
         );
  OAI21X1 U23252 ( .A(n28715), .B(n26101), .C(n28716), .Y(n28712) );
  AOI22X1 U23253 ( .A(n28572), .B(reg_A[65]), .C(n28224), .D(n28575), .Y(
        n28716) );
  AOI22X1 U23254 ( .A(reg_A[66]), .B(n28717), .C(reg_A[69]), .D(n25149), .Y(
        n28710) );
  AOI22X1 U23255 ( .A(reg_A[77]), .B(n25152), .C(reg_A[76]), .D(n25153), .Y(
        n28709) );
  NOR2X1 U23256 ( .A(n28718), .B(n28719), .Y(n28687) );
  OR2X1 U23257 ( .A(n28720), .B(n28721), .Y(n28719) );
  OAI22X1 U23258 ( .A(n28559), .B(n28722), .C(n28651), .D(n28646), .Y(n28721)
         );
  NAND2X1 U23259 ( .A(n28440), .B(n25170), .Y(n28646) );
  NOR2X1 U23260 ( .A(n26999), .B(reg_B[79]), .Y(n28440) );
  AOI22X1 U23261 ( .A(reg_A[72]), .B(n28546), .C(reg_A[74]), .D(n28251), .Y(
        n28651) );
  NOR2X1 U23262 ( .A(reg_B[77]), .B(reg_B[78]), .Y(n28251) );
  NOR2X1 U23263 ( .A(n28377), .B(reg_B[77]), .Y(n28546) );
  AOI21X1 U23264 ( .A(n27916), .B(n26197), .C(n28723), .Y(n28559) );
  OAI22X1 U23265 ( .A(n25894), .B(n26438), .C(n26131), .D(n25884), .Y(n27916)
         );
  OAI21X1 U23266 ( .A(n28383), .B(n28724), .C(n28725), .Y(n28720) );
  AOI22X1 U23267 ( .A(n28726), .B(reg_A[79]), .C(n28727), .D(n26974), .Y(
        n28725) );
  INVX1 U23268 ( .A(n28728), .Y(n28727) );
  INVX1 U23269 ( .A(n28607), .Y(n28383) );
  OAI21X1 U23270 ( .A(n25964), .B(n25884), .C(n28729), .Y(n28607) );
  AOI21X1 U23271 ( .A(reg_A[74]), .B(n26057), .C(n28723), .Y(n28729) );
  INVX1 U23272 ( .A(n28730), .Y(n28723) );
  NAND3X1 U23273 ( .A(n28731), .B(n28732), .C(n28733), .Y(n28718) );
  AOI22X1 U23274 ( .A(n25188), .B(n28734), .C(n28252), .D(n28735), .Y(n28733)
         );
  NOR2X1 U23275 ( .A(n28736), .B(n28737), .Y(n28252) );
  OAI22X1 U23276 ( .A(n28738), .B(n27454), .C(n27855), .D(n26599), .Y(n28737)
         );
  MUX2X1 U23277 ( .B(n26438), .A(n25884), .S(reg_B[1]), .Y(n27855) );
  OAI21X1 U23278 ( .A(reg_A[64]), .B(n28739), .C(n28740), .Y(n28736) );
  AOI22X1 U23279 ( .A(n28741), .B(n26101), .C(n28742), .D(n26547), .Y(n28740)
         );
  OAI21X1 U23280 ( .A(n28483), .B(n28241), .C(n28484), .Y(n28734) );
  NAND2X1 U23281 ( .A(n28743), .B(reg_B[77]), .Y(n28484) );
  NAND2X1 U23282 ( .A(n28744), .B(n28745), .Y(n28241) );
  AOI22X1 U23283 ( .A(n28602), .B(n26107), .C(n28191), .D(n25856), .Y(n28745)
         );
  AOI22X1 U23284 ( .A(n28245), .B(n25851), .C(n28446), .D(n26256), .Y(n28744)
         );
  OAI21X1 U23285 ( .A(n28746), .B(n28747), .C(n25310), .Y(n28732) );
  NAND3X1 U23286 ( .A(n28748), .B(n28749), .C(n28750), .Y(n28747) );
  NOR2X1 U23287 ( .A(n28751), .B(n28752), .Y(n28750) );
  OAI21X1 U23288 ( .A(n25036), .B(n26230), .C(n28753), .Y(n28752) );
  AOI22X1 U23289 ( .A(reg_A[82]), .B(n25124), .C(reg_A[85]), .D(n25222), .Y(
        n28753) );
  OAI21X1 U23290 ( .A(n25037), .B(n25875), .C(n28754), .Y(n28751) );
  AOI22X1 U23291 ( .A(reg_A[78]), .B(n25071), .C(reg_A[79]), .D(n25123), .Y(
        n28754) );
  AOI21X1 U23292 ( .A(reg_A[86]), .B(n25635), .C(n28755), .Y(n28749) );
  OAI22X1 U23293 ( .A(n25065), .B(n25929), .C(n25475), .D(n26195), .Y(n28755)
         );
  AOI22X1 U23294 ( .A(reg_A[87]), .B(n25325), .C(reg_A[74]), .D(n25125), .Y(
        n28748) );
  NAND3X1 U23295 ( .A(n28756), .B(n28757), .C(n28758), .Y(n28746) );
  NOR2X1 U23296 ( .A(n28759), .B(n28760), .Y(n28758) );
  OAI21X1 U23297 ( .A(n26719), .B(n25873), .C(n28761), .Y(n28760) );
  AOI22X1 U23298 ( .A(reg_A[92]), .B(n25241), .C(reg_A[94]), .D(n25339), .Y(
        n28761) );
  OAI21X1 U23299 ( .A(n25038), .B(n25881), .C(n28762), .Y(n28759) );
  AOI22X1 U23300 ( .A(reg_A[91]), .B(n25246), .C(reg_A[90]), .D(n25247), .Y(
        n28762) );
  AOI21X1 U23301 ( .A(reg_A[76]), .B(n25252), .C(n28763), .Y(n28757) );
  OAI22X1 U23302 ( .A(n25041), .B(n26286), .C(n25042), .D(n26103), .Y(n28763)
         );
  AOI22X1 U23303 ( .A(reg_A[80]), .B(n25253), .C(reg_A[81]), .D(n25628), .Y(
        n28756) );
  AOI22X1 U23304 ( .A(n28764), .B(n28765), .C(n28766), .D(n26149), .Y(n28731)
         );
  NOR2X1 U23305 ( .A(n28767), .B(n25198), .Y(n28766) );
  NOR2X1 U23306 ( .A(n28216), .B(n25087), .Y(n28764) );
  NOR2X1 U23307 ( .A(n28768), .B(n28769), .Y(n28686) );
  NAND2X1 U23308 ( .A(n28770), .B(n28771), .Y(n28769) );
  AOI22X1 U23309 ( .A(reg_A[72]), .B(n28772), .C(n28191), .D(n28773), .Y(
        n28771) );
  AOI22X1 U23310 ( .A(n26276), .B(n28774), .C(n26148), .D(n28497), .Y(n28770)
         );
  INVX1 U23311 ( .A(n28587), .Y(n28497) );
  AOI22X1 U23312 ( .A(n28775), .B(n25699), .C(n28776), .D(n25932), .Y(n28587)
         );
  NAND3X1 U23313 ( .A(n28777), .B(n28778), .C(n28779), .Y(n28768) );
  AOI22X1 U23314 ( .A(n26267), .B(n28780), .C(n28236), .D(n28192), .Y(n28779)
         );
  OAI22X1 U23315 ( .A(n28781), .B(n28782), .C(n25342), .D(n28783), .Y(n28236)
         );
  OAI21X1 U23316 ( .A(n28784), .B(n28193), .C(n25188), .Y(n28782) );
  OAI21X1 U23317 ( .A(n28645), .B(n28088), .C(n28785), .Y(n28781) );
  AOI22X1 U23318 ( .A(n28786), .B(n28295), .C(n28787), .D(reg_B[78]), .Y(
        n28785) );
  INVX1 U23319 ( .A(n28788), .Y(n28787) );
  OAI22X1 U23320 ( .A(reg_A[71]), .B(n28208), .C(reg_A[72]), .D(n28144), .Y(
        n28786) );
  MUX2X1 U23321 ( .B(n26438), .A(n25884), .S(reg_B[76]), .Y(n28645) );
  OAI21X1 U23322 ( .A(n28789), .B(n28208), .C(n28790), .Y(n28780) );
  AOI22X1 U23323 ( .A(n28446), .B(n28480), .C(n28602), .D(n28791), .Y(n28790)
         );
  OAI21X1 U23324 ( .A(n26438), .B(n28394), .C(n28792), .Y(n28480) );
  AOI22X1 U23325 ( .A(n28073), .B(reg_A[66]), .C(n28296), .D(reg_A[70]), .Y(
        n28792) );
  OAI21X1 U23326 ( .A(n28793), .B(n28794), .C(n26480), .Y(n28778) );
  OAI22X1 U23327 ( .A(n28316), .B(n26997), .C(n28221), .D(n25964), .Y(n28794)
         );
  INVX1 U23328 ( .A(n28795), .Y(n28221) );
  INVX1 U23329 ( .A(n28796), .Y(n28316) );
  OAI21X1 U23330 ( .A(n28222), .B(n28093), .C(n28797), .Y(n28793) );
  AOI22X1 U23331 ( .A(n28798), .B(n26114), .C(n26056), .D(n28799), .Y(n28797)
         );
  INVX1 U23332 ( .A(n28800), .Y(n28222) );
  AOI22X1 U23333 ( .A(n28454), .B(n28801), .C(n28802), .D(reg_A[78]), .Y(
        n28777) );
  INVX1 U23334 ( .A(n28217), .Y(n28454) );
  NAND2X1 U23335 ( .A(n28108), .B(n25382), .Y(n28217) );
  NAND3X1 U23336 ( .A(n28803), .B(n28804), .C(n28805), .Y(result[73]) );
  NOR2X1 U23337 ( .A(n28806), .B(n28807), .Y(n28805) );
  NAND3X1 U23338 ( .A(n28808), .B(n28809), .C(n28810), .Y(n28807) );
  NOR2X1 U23339 ( .A(n28811), .B(n28812), .Y(n28810) );
  OAI21X1 U23340 ( .A(n28813), .B(n25087), .C(n28557), .Y(n28812) );
  INVX1 U23341 ( .A(n28814), .Y(n28557) );
  OAI21X1 U23342 ( .A(n28192), .B(n28659), .C(n28815), .Y(n28814) );
  OAI21X1 U23343 ( .A(n28816), .B(n28114), .C(n25932), .Y(n28815) );
  INVX1 U23344 ( .A(n28230), .Y(n28114) );
  OAI21X1 U23345 ( .A(reg_B[93]), .B(reg_B[91]), .C(n26974), .Y(n28230) );
  NOR2X1 U23346 ( .A(n27027), .B(n25853), .Y(n28816) );
  NAND2X1 U23347 ( .A(reg_B[91]), .B(n26063), .Y(n27027) );
  AOI21X1 U23348 ( .A(n28108), .B(n28817), .C(n28818), .Y(n28813) );
  OAI21X1 U23349 ( .A(n28819), .B(n28820), .C(n28821), .Y(n28818) );
  OAI21X1 U23350 ( .A(n28822), .B(n28823), .C(n25044), .Y(n28821) );
  OAI21X1 U23351 ( .A(n28458), .B(n25964), .C(n28824), .Y(n28823) );
  AOI22X1 U23352 ( .A(n26057), .B(n28825), .C(n28826), .D(n28461), .Y(n28824)
         );
  INVX1 U23353 ( .A(n28827), .Y(n28458) );
  OAI21X1 U23354 ( .A(n28828), .B(n26997), .C(n28829), .Y(n28822) );
  AOI22X1 U23355 ( .A(n28798), .B(n28460), .C(n26056), .D(n28830), .Y(n28829)
         );
  INVX1 U23356 ( .A(n28340), .Y(n28828) );
  INVX1 U23357 ( .A(n28831), .Y(n28811) );
  MUX2X1 U23358 ( .B(n28416), .A(n28773), .S(n28446), .Y(n28831) );
  OAI21X1 U23359 ( .A(n28478), .B(n26147), .C(n28832), .Y(n28773) );
  OAI21X1 U23360 ( .A(n28833), .B(n28589), .C(reg_A[73]), .Y(n28832) );
  INVX1 U23361 ( .A(n28414), .Y(n28589) );
  NAND2X1 U23362 ( .A(n26504), .B(n28192), .Y(n28414) );
  NOR2X1 U23363 ( .A(reg_B[77]), .B(n26151), .Y(n28833) );
  INVX1 U23364 ( .A(n28603), .Y(n28478) );
  OAI21X1 U23365 ( .A(n26439), .B(n28394), .C(n28834), .Y(n28603) );
  AOI22X1 U23366 ( .A(n28073), .B(reg_A[65]), .C(n28296), .D(reg_A[69]), .Y(
        n28834) );
  INVX1 U23367 ( .A(n28659), .Y(n28416) );
  NAND2X1 U23368 ( .A(reg_A[72]), .B(n26504), .Y(n28659) );
  AOI22X1 U23369 ( .A(reg_A[73]), .B(n28835), .C(reg_A[64]), .D(n25137), .Y(
        n28809) );
  AOI22X1 U23370 ( .A(reg_A[71]), .B(n25138), .C(n28836), .D(n25119), .Y(
        n28808) );
  NAND3X1 U23371 ( .A(n28837), .B(n28838), .C(n28839), .Y(n28836) );
  NOR2X1 U23372 ( .A(n28840), .B(n28841), .Y(n28839) );
  OAI22X1 U23373 ( .A(n25030), .B(n25884), .C(n25131), .D(n25851), .Y(n28841)
         );
  OAI21X1 U23374 ( .A(n25040), .B(n26101), .C(n28842), .Y(n28840) );
  AOI22X1 U23375 ( .A(reg_A[72]), .B(n25135), .C(reg_A[70]), .D(n25136), .Y(
        n28842) );
  AOI22X1 U23376 ( .A(reg_A[69]), .B(n25071), .C(reg_A[68]), .D(n25123), .Y(
        n28838) );
  AOI22X1 U23377 ( .A(reg_A[65]), .B(n25124), .C(reg_A[73]), .D(n25125), .Y(
        n28837) );
  NAND3X1 U23378 ( .A(n28843), .B(n28844), .C(n28845), .Y(n28806) );
  AOI21X1 U23379 ( .A(reg_A[74]), .B(n28280), .C(n28846), .Y(n28845) );
  OAI22X1 U23380 ( .A(n28569), .B(n26103), .C(n28570), .D(n25863), .Y(n28846)
         );
  AOI22X1 U23381 ( .A(reg_A[69]), .B(n25181), .C(reg_A[65]), .D(n28717), .Y(
        n28844) );
  AOI22X1 U23382 ( .A(reg_A[68]), .B(n25149), .C(n28847), .D(n25150), .Y(
        n28843) );
  INVX1 U23383 ( .A(n28663), .Y(n28847) );
  NAND2X1 U23384 ( .A(n28848), .B(n28849), .Y(n28663) );
  AOI22X1 U23385 ( .A(n26859), .B(n26107), .C(n26860), .D(n25856), .Y(n28849)
         );
  AOI22X1 U23386 ( .A(n26455), .B(n25853), .C(n28401), .D(n26452), .Y(n28848)
         );
  OAI21X1 U23387 ( .A(reg_A[64]), .B(n26861), .C(n28850), .Y(n28401) );
  AOI22X1 U23388 ( .A(n28851), .B(n26863), .C(n26462), .D(n26547), .Y(n28850)
         );
  INVX1 U23389 ( .A(n28738), .Y(n28851) );
  MUX2X1 U23390 ( .B(n26439), .A(n25855), .S(reg_B[1]), .Y(n28738) );
  NOR2X1 U23391 ( .A(n28852), .B(n28853), .Y(n28804) );
  OAI21X1 U23392 ( .A(n26881), .B(n28683), .C(n28854), .Y(n28853) );
  AOI22X1 U23393 ( .A(n28855), .B(n28776), .C(n28647), .D(n28775), .Y(n28854)
         );
  INVX1 U23394 ( .A(n28856), .Y(n28775) );
  AOI21X1 U23395 ( .A(n27882), .B(n26197), .C(n28857), .Y(n28856) );
  OAI22X1 U23396 ( .A(n26439), .B(n25894), .C(n25855), .D(n26131), .Y(n27882)
         );
  OAI21X1 U23397 ( .A(n25855), .B(n25964), .C(n28858), .Y(n28776) );
  AOI21X1 U23398 ( .A(n26057), .B(reg_A[73]), .C(n28857), .Y(n28858) );
  NOR2X1 U23399 ( .A(n26997), .B(n25856), .Y(n28857) );
  INVX1 U23400 ( .A(n28134), .Y(n28683) );
  NAND3X1 U23401 ( .A(n28859), .B(n28860), .C(n28861), .Y(n28852) );
  AOI22X1 U23402 ( .A(n28862), .B(n26756), .C(n26267), .D(n28863), .Y(n28861)
         );
  OAI22X1 U23403 ( .A(n28864), .B(n28208), .C(n28789), .D(n28144), .Y(n28863)
         );
  OAI22X1 U23404 ( .A(n28865), .B(n26169), .C(n28767), .D(n25914), .Y(n28862)
         );
  NAND3X1 U23405 ( .A(n25170), .B(n28866), .C(n28191), .Y(n28860) );
  NAND3X1 U23406 ( .A(n25932), .B(n25972), .C(n26974), .Y(n28859) );
  NOR2X1 U23407 ( .A(n28867), .B(n28868), .Y(n28803) );
  OAI21X1 U23408 ( .A(n28715), .B(n26256), .C(n28869), .Y(n28868) );
  AOI22X1 U23409 ( .A(n26148), .B(n28774), .C(reg_A[72]), .D(n25174), .Y(
        n28869) );
  INVX1 U23410 ( .A(n28870), .Y(n25174) );
  INVX1 U23411 ( .A(n28588), .Y(n28774) );
  AOI22X1 U23412 ( .A(n28871), .B(n25699), .C(n28872), .D(n25932), .Y(n28588)
         );
  OR2X1 U23413 ( .A(n28873), .B(n28874), .Y(n28867) );
  OAI21X1 U23414 ( .A(n25184), .B(n25884), .C(n28875), .Y(n28874) );
  OAI21X1 U23415 ( .A(n28876), .B(n28877), .C(n25188), .Y(n28875) );
  OAI21X1 U23416 ( .A(n28878), .B(n28879), .C(n28880), .Y(n28877) );
  INVX1 U23417 ( .A(n28881), .Y(n28880) );
  MUX2X1 U23418 ( .B(n28615), .A(n28882), .S(reg_B[78]), .Y(n28881) );
  OAI21X1 U23419 ( .A(reg_B[77]), .B(n28391), .C(n28883), .Y(n28615) );
  AOI21X1 U23420 ( .A(n28296), .B(n28884), .C(n28642), .Y(n28883) );
  NOR2X1 U23421 ( .A(n28788), .B(n28192), .Y(n28642) );
  INVX1 U23422 ( .A(n28392), .Y(n28884) );
  MUX2X1 U23423 ( .B(n25856), .A(n26107), .S(reg_B[79]), .Y(n28392) );
  MUX2X1 U23424 ( .B(n28885), .A(n28886), .S(reg_B[79]), .Y(n28391) );
  OAI21X1 U23425 ( .A(reg_B[76]), .B(reg_A[72]), .C(n28788), .Y(n28886) );
  NAND2X1 U23426 ( .A(reg_B[76]), .B(n25853), .Y(n28788) );
  INVX1 U23427 ( .A(n28784), .Y(n28885) );
  MUX2X1 U23428 ( .B(n26439), .A(n25855), .S(reg_B[76]), .Y(n28784) );
  INVX1 U23429 ( .A(n28072), .Y(n28878) );
  MUX2X1 U23430 ( .B(n26101), .A(n26256), .S(reg_B[79]), .Y(n28072) );
  OAI21X1 U23431 ( .A(n28208), .B(n28887), .C(n28888), .Y(n28876) );
  NAND3X1 U23432 ( .A(n28296), .B(reg_A[67]), .C(n28602), .Y(n28888) );
  OAI21X1 U23433 ( .A(n25162), .B(n25851), .C(n28889), .Y(n28873) );
  OAI21X1 U23434 ( .A(n28890), .B(n28891), .C(n25203), .Y(n28889) );
  OAI22X1 U23435 ( .A(n25204), .B(n26439), .C(n25205), .D(n26286), .Y(n28891)
         );
  OAI21X1 U23436 ( .A(n25207), .B(n25865), .C(n28892), .Y(n28890) );
  AOI22X1 U23437 ( .A(n25097), .B(n28893), .C(reg_A[79]), .D(n25211), .Y(
        n28892) );
  NAND3X1 U23438 ( .A(n28894), .B(n28895), .C(n28896), .Y(n28893) );
  AND2X1 U23439 ( .A(n28897), .B(n28898), .Y(n28896) );
  NOR2X1 U23440 ( .A(n28899), .B(n28900), .Y(n28898) );
  OAI21X1 U23441 ( .A(n25036), .B(n25875), .C(n28901), .Y(n28900) );
  AOI22X1 U23442 ( .A(reg_A[81]), .B(n25124), .C(reg_A[84]), .D(n25222), .Y(
        n28901) );
  OAI21X1 U23443 ( .A(n25037), .B(n25874), .C(n28902), .Y(n28899) );
  AOI22X1 U23444 ( .A(reg_A[77]), .B(n25072), .C(reg_A[78]), .D(n25123), .Y(
        n28902) );
  NOR2X1 U23445 ( .A(n28903), .B(n28904), .Y(n28897) );
  OAI22X1 U23446 ( .A(n25043), .B(n26439), .C(n25039), .D(n26039), .Y(n28904)
         );
  OAI21X1 U23447 ( .A(n25064), .B(n26215), .C(n28905), .Y(n28903) );
  AOI22X1 U23448 ( .A(reg_A[87]), .B(n25234), .C(reg_A[88]), .D(n25235), .Y(
        n28905) );
  NOR2X1 U23449 ( .A(n28906), .B(n28907), .Y(n28895) );
  OAI21X1 U23450 ( .A(n25238), .B(n25881), .C(n28908), .Y(n28907) );
  AOI22X1 U23451 ( .A(reg_A[91]), .B(n25241), .C(reg_A[95]), .D(n25242), .Y(
        n28908) );
  OAI21X1 U23452 ( .A(n25038), .B(n25882), .C(n28909), .Y(n28906) );
  AOI22X1 U23453 ( .A(reg_A[90]), .B(n25246), .C(reg_A[89]), .D(n25247), .Y(
        n28909) );
  NOR2X1 U23454 ( .A(n28910), .B(n28911), .Y(n28894) );
  OAI21X1 U23455 ( .A(n25030), .B(n25584), .C(n28912), .Y(n28911) );
  AOI22X1 U23456 ( .A(reg_A[75]), .B(n25252), .C(reg_A[79]), .D(n25253), .Y(
        n28912) );
  OAI21X1 U23457 ( .A(n25041), .B(n25863), .C(n28913), .Y(n28910) );
  AOI22X1 U23458 ( .A(reg_A[94]), .B(n25257), .C(reg_A[74]), .D(n25135), .Y(
        n28913) );
  NAND3X1 U23459 ( .A(n28914), .B(n28915), .C(n28916), .Y(result[72]) );
  NOR2X1 U23460 ( .A(n28917), .B(n28918), .Y(n28916) );
  OR2X1 U23461 ( .A(n28919), .B(n28920), .Y(n28918) );
  OAI21X1 U23462 ( .A(n28921), .B(n25087), .C(n28922), .Y(n28920) );
  AOI22X1 U23463 ( .A(reg_A[72]), .B(n26690), .C(reg_A[73]), .D(n28923), .Y(
        n28922) );
  AOI21X1 U23464 ( .A(n28108), .B(n28924), .C(n28925), .Y(n28921) );
  OAI21X1 U23465 ( .A(n28503), .B(n28820), .C(n28926), .Y(n28925) );
  OAI21X1 U23466 ( .A(n28927), .B(n28928), .C(n25044), .Y(n28926) );
  OAI21X1 U23467 ( .A(n28507), .B(n25964), .C(n28929), .Y(n28928) );
  AOI22X1 U23468 ( .A(n28826), .B(n28509), .C(n28930), .D(n28931), .Y(n28929)
         );
  OAI21X1 U23469 ( .A(n28932), .B(n25966), .C(n28933), .Y(n28927) );
  AOI22X1 U23470 ( .A(n28798), .B(n26992), .C(n26056), .D(n26915), .Y(n28933)
         );
  INVX1 U23471 ( .A(n25967), .Y(n26056) );
  NAND2X1 U23472 ( .A(reg_B[91]), .B(n26275), .Y(n25967) );
  NOR2X1 U23473 ( .A(n26069), .B(n25895), .Y(n28798) );
  INVX1 U23474 ( .A(n28765), .Y(n28820) );
  NOR2X1 U23475 ( .A(n28192), .B(n28102), .Y(n28765) );
  INVX1 U23476 ( .A(n28934), .Y(n28503) );
  NOR2X1 U23477 ( .A(reg_B[77]), .B(n28102), .Y(n28108) );
  AOI21X1 U23478 ( .A(n28295), .B(n25604), .C(n25589), .Y(n28102) );
  OAI21X1 U23479 ( .A(n28935), .B(n26438), .C(n28936), .Y(n28919) );
  AOI22X1 U23480 ( .A(n28573), .B(n28575), .C(reg_A[75]), .D(n26739), .Y(
        n28936) );
  INVX1 U23481 ( .A(n26783), .Y(n28935) );
  NAND3X1 U23482 ( .A(n28937), .B(n28938), .C(n28939), .Y(n28917) );
  AOI21X1 U23483 ( .A(reg_A[71]), .B(n26749), .C(n28940), .Y(n28939) );
  INVX1 U23484 ( .A(n28941), .Y(n28940) );
  AOI22X1 U23485 ( .A(n26748), .B(reg_A[79]), .C(n26747), .D(reg_A[78]), .Y(
        n28941) );
  AOI22X1 U23486 ( .A(reg_A[70]), .B(n28942), .C(reg_A[76]), .D(n28943), .Y(
        n28938) );
  AOI22X1 U23487 ( .A(reg_A[65]), .B(n26673), .C(reg_A[77]), .D(n26746), .Y(
        n28937) );
  NOR2X1 U23488 ( .A(n28944), .B(n28945), .Y(n28915) );
  OAI21X1 U23489 ( .A(n25198), .B(n28946), .C(n28947), .Y(n28945) );
  AOI22X1 U23490 ( .A(n28647), .B(n28871), .C(n28574), .D(n27008), .Y(n28947)
         );
  AND2X1 U23491 ( .A(n28948), .B(n28949), .Y(n28574) );
  AOI22X1 U23492 ( .A(n26601), .B(n26256), .C(n26602), .D(n25856), .Y(n28949)
         );
  AOI22X1 U23493 ( .A(n27012), .B(n26547), .C(n26597), .D(n26101), .Y(n28948)
         );
  OAI21X1 U23494 ( .A(n28950), .B(reg_B[93]), .C(n28951), .Y(n28871) );
  INVX1 U23495 ( .A(n28319), .Y(n28950) );
  OAI22X1 U23496 ( .A(n26131), .B(n25853), .C(n25894), .D(n26547), .Y(n28319)
         );
  INVX1 U23497 ( .A(n28722), .Y(n28647) );
  AOI21X1 U23498 ( .A(n26149), .B(n28952), .C(n28953), .Y(n28946) );
  OAI22X1 U23499 ( .A(n28865), .B(n25914), .C(n28767), .D(n26168), .Y(n28953)
         );
  NAND3X1 U23500 ( .A(n28954), .B(n28955), .C(n28956), .Y(n28944) );
  AOI22X1 U23501 ( .A(reg_A[64]), .B(n28957), .C(n28855), .D(n28872), .Y(
        n28956) );
  OAI21X1 U23502 ( .A(n25966), .B(n26547), .C(n28951), .Y(n28872) );
  NAND2X1 U23503 ( .A(n28930), .B(reg_A[68]), .Y(n28951) );
  INVX1 U23504 ( .A(n28724), .Y(n28855) );
  OAI21X1 U23505 ( .A(n26134), .B(n27438), .C(n26743), .Y(n28957) );
  INVX1 U23506 ( .A(n28958), .Y(n26743) );
  INVX1 U23507 ( .A(n25894), .Y(n26134) );
  NAND2X1 U23508 ( .A(n25895), .B(n26063), .Y(n25894) );
  OAI21X1 U23509 ( .A(n28959), .B(n28960), .C(n25310), .Y(n28955) );
  NAND2X1 U23510 ( .A(n28961), .B(n28962), .Y(n28960) );
  NOR2X1 U23511 ( .A(n28963), .B(n28964), .Y(n28962) );
  OAI21X1 U23512 ( .A(n25043), .B(n26547), .C(n28965), .Y(n28964) );
  AOI22X1 U23513 ( .A(reg_A[73]), .B(n25135), .C(reg_A[74]), .D(n25252), .Y(
        n28965) );
  OAI21X1 U23514 ( .A(n25028), .B(n26286), .C(n28966), .Y(n28963) );
  AOI22X1 U23515 ( .A(reg_A[75]), .B(n25136), .C(reg_A[76]), .D(n25068), .Y(
        n28966) );
  NOR2X1 U23516 ( .A(n28967), .B(n28968), .Y(n28961) );
  OAI21X1 U23517 ( .A(n25034), .B(n25584), .C(n28969), .Y(n28968) );
  AOI22X1 U23518 ( .A(reg_A[78]), .B(n25253), .C(reg_A[79]), .D(n25628), .Y(
        n28969) );
  OAI21X1 U23519 ( .A(n25036), .B(n25874), .C(n28970), .Y(n28967) );
  AOI22X1 U23520 ( .A(reg_A[81]), .B(n25629), .C(reg_A[83]), .D(n25222), .Y(
        n28970) );
  NAND2X1 U23521 ( .A(n28971), .B(n28972), .Y(n28959) );
  NOR2X1 U23522 ( .A(n28973), .B(n28974), .Y(n28972) );
  OAI21X1 U23523 ( .A(n25039), .B(n26215), .C(n28975), .Y(n28974) );
  AOI22X1 U23524 ( .A(reg_A[86]), .B(n25234), .C(reg_A[84]), .D(n25635), .Y(
        n28975) );
  OAI21X1 U23525 ( .A(n25065), .B(n25965), .C(n28976), .Y(n28973) );
  AOI22X1 U23526 ( .A(reg_A[89]), .B(n25246), .C(reg_A[88]), .D(n25247), .Y(
        n28976) );
  NOR2X1 U23527 ( .A(n28977), .B(n28978), .Y(n28971) );
  OAI21X1 U23528 ( .A(n25238), .B(n25882), .C(n28979), .Y(n28978) );
  AOI22X1 U23529 ( .A(reg_A[91]), .B(n25487), .C(reg_A[90]), .D(n25241), .Y(
        n28979) );
  OAI21X1 U23530 ( .A(n26719), .B(n25881), .C(n28980), .Y(n28977) );
  AOI22X1 U23531 ( .A(reg_A[94]), .B(n25242), .C(reg_A[95]), .D(n25338), .Y(
        n28980) );
  NAND3X1 U23532 ( .A(n25170), .B(n28866), .C(n28446), .Y(n28954) );
  OAI21X1 U23533 ( .A(n28600), .B(n25415), .C(n28981), .Y(n28866) );
  NAND3X1 U23534 ( .A(n25589), .B(n28192), .C(reg_A[72]), .Y(n28981) );
  INVX1 U23535 ( .A(n28791), .Y(n28600) );
  OAI21X1 U23536 ( .A(n26547), .B(n28394), .C(n28982), .Y(n28791) );
  AOI22X1 U23537 ( .A(n28743), .B(n28192), .C(n28296), .D(reg_A[68]), .Y(
        n28982) );
  INVX1 U23538 ( .A(n28882), .Y(n28743) );
  NOR2X1 U23539 ( .A(n28983), .B(n28984), .Y(n28914) );
  OAI21X1 U23540 ( .A(n28985), .B(n25856), .C(n28986), .Y(n28984) );
  AOI22X1 U23541 ( .A(reg_A[67]), .B(n26679), .C(reg_A[68]), .D(n26680), .Y(
        n28986) );
  INVX1 U23542 ( .A(n26681), .Y(n28985) );
  OAI21X1 U23543 ( .A(n28987), .B(n25884), .C(n28988), .Y(n28983) );
  AOI22X1 U23544 ( .A(n26267), .B(n28989), .C(n25188), .D(n28990), .Y(n28988)
         );
  OAI21X1 U23545 ( .A(n28394), .B(n28490), .C(n28991), .Y(n28990) );
  INVX1 U23546 ( .A(n28992), .Y(n28991) );
  OAI21X1 U23547 ( .A(n28489), .B(n28483), .C(n28882), .Y(n28992) );
  NAND2X1 U23548 ( .A(n28993), .B(n28994), .Y(n28489) );
  AOI22X1 U23549 ( .A(n28602), .B(n25884), .C(n28191), .D(n25851), .Y(n28994)
         );
  AOI22X1 U23550 ( .A(n28245), .B(n25855), .C(n28446), .D(n26107), .Y(n28993)
         );
  NAND2X1 U23551 ( .A(n28995), .B(n28996), .Y(n28490) );
  AOI22X1 U23552 ( .A(n28602), .B(n26256), .C(n28191), .D(n26101), .Y(n28996)
         );
  AOI22X1 U23553 ( .A(n28245), .B(n25856), .C(n28446), .D(n26547), .Y(n28995)
         );
  OAI21X1 U23554 ( .A(n28997), .B(n28208), .C(n28998), .Y(n28989) );
  AOI22X1 U23555 ( .A(n28191), .B(n28999), .C(n28602), .D(n29000), .Y(n28998)
         );
  INVX1 U23556 ( .A(n26678), .Y(n28987) );
  NAND3X1 U23557 ( .A(n29001), .B(n29002), .C(n29003), .Y(result[71]) );
  NOR2X1 U23558 ( .A(n29004), .B(n29005), .Y(n29003) );
  NAND3X1 U23559 ( .A(n29006), .B(n29007), .C(n29008), .Y(n29005) );
  NOR2X1 U23560 ( .A(n29009), .B(n29010), .Y(n29008) );
  OAI21X1 U23561 ( .A(n27354), .B(n29011), .C(n29012), .Y(n29010) );
  OAI21X1 U23562 ( .A(n29013), .B(n29014), .C(n25170), .Y(n29012) );
  OAI21X1 U23563 ( .A(n26101), .B(n29015), .C(n29016), .Y(n29014) );
  OAI21X1 U23564 ( .A(n29017), .B(n29018), .C(n25044), .Y(n29016) );
  AND2X1 U23565 ( .A(n29019), .B(n26149), .Y(n29017) );
  OAI21X1 U23566 ( .A(n29020), .B(n29021), .C(n29022), .Y(n29013) );
  NAND3X1 U23567 ( .A(n25604), .B(n29023), .C(n28245), .Y(n29022) );
  MUX2X1 U23568 ( .B(n29024), .A(n29025), .S(reg_B[70]), .Y(n29021) );
  NOR2X1 U23569 ( .A(n25851), .B(n29026), .Y(n29024) );
  AOI21X1 U23570 ( .A(n28602), .B(n29027), .C(n29028), .Y(n29011) );
  OAI22X1 U23571 ( .A(n28864), .B(n28193), .C(n28789), .D(n28088), .Y(n29028)
         );
  INVX1 U23572 ( .A(n28999), .Y(n28789) );
  OAI22X1 U23573 ( .A(n26101), .B(n28394), .C(n25851), .D(n28483), .Y(n28999)
         );
  AOI22X1 U23574 ( .A(reg_A[75]), .B(n29029), .C(reg_A[76]), .D(n29030), .Y(
        n29007) );
  AOI22X1 U23575 ( .A(reg_A[77]), .B(n29031), .C(reg_A[78]), .D(n25293), .Y(
        n29006) );
  NAND2X1 U23576 ( .A(n29032), .B(n29033), .Y(n29004) );
  NOR2X1 U23577 ( .A(n29034), .B(n29035), .Y(n29033) );
  OAI21X1 U23578 ( .A(n29036), .B(n26547), .C(n29037), .Y(n29035) );
  OAI21X1 U23579 ( .A(n29038), .B(n29039), .C(n25310), .Y(n29037) );
  NAND3X1 U23580 ( .A(n29040), .B(n29041), .C(n29042), .Y(n29039) );
  NOR2X1 U23581 ( .A(n29043), .B(n29044), .Y(n29042) );
  OAI22X1 U23582 ( .A(n25036), .B(n26094), .C(n25473), .D(n25874), .Y(n29044)
         );
  OAI22X1 U23583 ( .A(n25037), .B(n25584), .C(n25320), .D(n25873), .Y(n29043)
         );
  AOI22X1 U23584 ( .A(reg_A[85]), .B(n25234), .C(reg_A[86]), .D(n25235), .Y(
        n29041) );
  AOI22X1 U23585 ( .A(reg_A[83]), .B(n25635), .C(reg_A[84]), .D(n25325), .Y(
        n29040) );
  NAND3X1 U23586 ( .A(n29045), .B(n29046), .C(n29047), .Y(n29038) );
  NOR2X1 U23587 ( .A(n29048), .B(n29049), .Y(n29047) );
  OAI22X1 U23588 ( .A(n25331), .B(n25929), .C(n25243), .D(n26068), .Y(n29049)
         );
  OAI22X1 U23589 ( .A(n25334), .B(n25965), .C(n25336), .D(n26195), .Y(n29048)
         );
  AOI22X1 U23590 ( .A(reg_A[93]), .B(n25242), .C(reg_A[94]), .D(n25338), .Y(
        n29046) );
  AOI22X1 U23591 ( .A(reg_A[91]), .B(n25339), .C(reg_A[92]), .D(n25257), .Y(
        n29045) );
  OAI22X1 U23592 ( .A(n25945), .B(n29050), .C(n27964), .D(n26101), .Y(n29034)
         );
  AOI21X1 U23593 ( .A(reg_A[74]), .B(n29051), .C(n29052), .Y(n29032) );
  OAI22X1 U23594 ( .A(n27938), .B(n26439), .C(n27512), .D(n25864), .Y(n29052)
         );
  NOR2X1 U23595 ( .A(n29053), .B(n29054), .Y(n29002) );
  OAI21X1 U23596 ( .A(n28208), .B(n29055), .C(n29056), .Y(n29054) );
  AOI22X1 U23597 ( .A(n29057), .B(n29058), .C(n28134), .D(n27110), .Y(n29056)
         );
  MUX2X1 U23598 ( .B(n26101), .A(n26256), .S(reg_B[4]), .Y(n28134) );
  NAND3X1 U23599 ( .A(n29059), .B(n29060), .C(n29061), .Y(n29053) );
  AND2X1 U23600 ( .A(n29062), .B(n29063), .Y(n29061) );
  OAI21X1 U23601 ( .A(n29064), .B(n29018), .C(n25932), .Y(n29063) );
  OAI22X1 U23602 ( .A(n29065), .B(n25914), .C(n28865), .D(n26168), .Y(n29018)
         );
  INVX1 U23603 ( .A(n29066), .Y(n28865) );
  AOI21X1 U23604 ( .A(n29067), .B(n29068), .C(n26169), .Y(n29064) );
  OAI21X1 U23605 ( .A(n29069), .B(n28004), .C(reg_A[68]), .Y(n29062) );
  OAI21X1 U23606 ( .A(n29070), .B(n29071), .C(n27067), .Y(n29060) );
  OAI21X1 U23607 ( .A(n25060), .B(n26101), .C(n29072), .Y(n29071) );
  AOI22X1 U23608 ( .A(reg_A[67]), .B(n25749), .C(reg_A[66]), .D(n25750), .Y(
        n29072) );
  NAND2X1 U23609 ( .A(n29073), .B(n29074), .Y(n29070) );
  AOI22X1 U23610 ( .A(reg_A[70]), .B(n26803), .C(reg_A[68]), .D(n26804), .Y(
        n29074) );
  AOI22X1 U23611 ( .A(reg_A[69]), .B(n26927), .C(reg_A[65]), .D(n26878), .Y(
        n29073) );
  OAI21X1 U23612 ( .A(n29075), .B(n29076), .C(n25119), .Y(n29059) );
  OAI21X1 U23613 ( .A(n25043), .B(n26101), .C(n29077), .Y(n29076) );
  AOI22X1 U23614 ( .A(reg_A[67]), .B(n25071), .C(reg_A[66]), .D(n25123), .Y(
        n29077) );
  NAND2X1 U23615 ( .A(n29078), .B(n29079), .Y(n29075) );
  AOI22X1 U23616 ( .A(reg_A[70]), .B(n25135), .C(reg_A[68]), .D(n25136), .Y(
        n29079) );
  AOI22X1 U23617 ( .A(reg_A[69]), .B(n25252), .C(reg_A[65]), .D(n25253), .Y(
        n29078) );
  NOR2X1 U23618 ( .A(n29080), .B(n29081), .Y(n29001) );
  OAI21X1 U23619 ( .A(n29082), .B(n25853), .C(n29083), .Y(n29081) );
  AOI22X1 U23620 ( .A(n29084), .B(n29085), .C(n27132), .D(reg_A[67]), .Y(
        n29083) );
  INVX1 U23621 ( .A(n28767), .Y(n29085) );
  AOI21X1 U23622 ( .A(reg_A[67]), .B(n28930), .C(n29086), .Y(n28767) );
  NAND3X1 U23623 ( .A(n29087), .B(n29088), .C(n29089), .Y(n29080) );
  AOI22X1 U23624 ( .A(n28050), .B(reg_A[66]), .C(n25999), .D(n29090), .Y(
        n29089) );
  OAI21X1 U23625 ( .A(n25754), .B(n25855), .C(n29091), .Y(n29090) );
  AOI22X1 U23626 ( .A(reg_A[70]), .B(n26007), .C(reg_A[69]), .D(n26009), .Y(
        n29091) );
  OAI21X1 U23627 ( .A(n29092), .B(n29093), .C(n26504), .Y(n29088) );
  OAI22X1 U23628 ( .A(n29094), .B(n29095), .C(n29096), .D(n29097), .Y(n29093)
         );
  MUX2X1 U23629 ( .B(reg_A[71]), .A(reg_A[67]), .S(reg_B[69]), .Y(n29097) );
  AND2X1 U23630 ( .A(reg_B[70]), .B(n29098), .Y(n29092) );
  OAI21X1 U23631 ( .A(n29099), .B(n29100), .C(n25382), .Y(n29087) );
  OAI21X1 U23632 ( .A(n29101), .B(n29102), .C(n29103), .Y(n29100) );
  AOI22X1 U23633 ( .A(n29104), .B(reg_A[71]), .C(n29086), .D(n25963), .Y(
        n29103) );
  INVX1 U23634 ( .A(n29015), .Y(n29104) );
  INVX1 U23635 ( .A(n29105), .Y(n29101) );
  OAI21X1 U23636 ( .A(n29106), .B(n29107), .C(n29108), .Y(n29099) );
  AND2X1 U23637 ( .A(n29109), .B(n29110), .Y(n29108) );
  NAND3X1 U23638 ( .A(n28103), .B(reg_A[79]), .C(n28446), .Y(n29110) );
  OAI21X1 U23639 ( .A(n29111), .B(n29112), .C(n25044), .Y(n29109) );
  OAI22X1 U23640 ( .A(n28660), .B(n26997), .C(n28596), .D(n25964), .Y(n29112)
         );
  INVX1 U23641 ( .A(n28084), .Y(n28596) );
  OAI21X1 U23642 ( .A(n28095), .B(n28093), .C(n29113), .Y(n29111) );
  AOI22X1 U23643 ( .A(n26057), .B(n29114), .C(reg_B[91]), .D(n27150), .Y(
        n29113) );
  OAI21X1 U23644 ( .A(n28092), .B(n26069), .C(n29115), .Y(n27150) );
  AOI22X1 U23645 ( .A(n25902), .B(n25988), .C(n26275), .D(n28597), .Y(n29115)
         );
  INVX1 U23646 ( .A(n29116), .Y(n28092) );
  INVX1 U23647 ( .A(n29117), .Y(n28095) );
  INVX1 U23648 ( .A(n29118), .Y(n29106) );
  NAND3X1 U23649 ( .A(n29119), .B(n29120), .C(n29121), .Y(result[70]) );
  NOR2X1 U23650 ( .A(n29122), .B(n29123), .Y(n29121) );
  NAND3X1 U23651 ( .A(n29124), .B(n29125), .C(n29126), .Y(n29123) );
  AOI21X1 U23652 ( .A(reg_A[64]), .B(n29127), .C(n29128), .Y(n29126) );
  OAI22X1 U23653 ( .A(n29129), .B(n25884), .C(n26781), .D(n26101), .Y(n29128)
         );
  AOI21X1 U23654 ( .A(reg_A[65]), .B(n29130), .C(n29131), .Y(n29124) );
  AOI21X1 U23655 ( .A(n29132), .B(n29133), .C(n25087), .Y(n29131) );
  AOI21X1 U23656 ( .A(n29134), .B(n28801), .C(n29135), .Y(n29133) );
  OAI21X1 U23657 ( .A(n29136), .B(n29137), .C(n29138), .Y(n29135) );
  OAI21X1 U23658 ( .A(n29139), .B(n29140), .C(n25044), .Y(n29138) );
  OAI21X1 U23659 ( .A(n28696), .B(n26997), .C(n29141), .Y(n29140) );
  AOI22X1 U23660 ( .A(n28826), .B(n28795), .C(n26307), .D(n28796), .Y(n29141)
         );
  OAI21X1 U23661 ( .A(n29142), .B(n25895), .C(n29143), .Y(n29139) );
  AOI22X1 U23662 ( .A(n26057), .B(n29144), .C(n29086), .D(n26148), .Y(n29143)
         );
  NOR2X1 U23663 ( .A(n26101), .B(n25966), .Y(n29086) );
  INVX1 U23664 ( .A(n27270), .Y(n29142) );
  OAI21X1 U23665 ( .A(n26624), .B(n26069), .C(n29145), .Y(n27270) );
  AOI22X1 U23666 ( .A(n26275), .B(n28800), .C(n25988), .D(n26114), .Y(n29145)
         );
  INVX1 U23667 ( .A(n28799), .Y(n26624) );
  AOI21X1 U23668 ( .A(n29146), .B(n29147), .C(n29148), .Y(n29132) );
  OAI22X1 U23669 ( .A(n28216), .B(n29149), .C(n29150), .D(n29151), .Y(n29148)
         );
  NAND3X1 U23670 ( .A(n29152), .B(n29153), .C(n29154), .Y(n29122) );
  AOI21X1 U23671 ( .A(reg_A[67]), .B(n29155), .C(n29156), .Y(n29154) );
  OAI21X1 U23672 ( .A(n29157), .B(n25856), .C(n29158), .Y(n29156) );
  OAI21X1 U23673 ( .A(n29159), .B(n29160), .C(n25310), .Y(n29158) );
  NAND3X1 U23674 ( .A(n29161), .B(n29162), .C(n29163), .Y(n29160) );
  NOR2X1 U23675 ( .A(n29164), .B(n29165), .Y(n29163) );
  OAI21X1 U23676 ( .A(n25043), .B(n26256), .C(n29166), .Y(n29165) );
  AOI22X1 U23677 ( .A(reg_A[82]), .B(n25635), .C(reg_A[83]), .D(n25325), .Y(
        n29166) );
  OAI21X1 U23678 ( .A(n25065), .B(n26215), .C(n29167), .Y(n29164) );
  AOI22X1 U23679 ( .A(reg_A[80]), .B(n25637), .C(reg_A[84]), .D(n25234), .Y(
        n29167) );
  NOR2X1 U23680 ( .A(n29168), .B(n29169), .Y(n29162) );
  OAI22X1 U23681 ( .A(n25028), .B(n26103), .C(n26431), .D(n26438), .Y(n29169)
         );
  OAI22X1 U23682 ( .A(n25030), .B(n26286), .C(n25131), .D(n25863), .Y(n29168)
         );
  AOI21X1 U23683 ( .A(reg_A[81]), .B(n25222), .C(n29170), .Y(n29161) );
  OAI22X1 U23684 ( .A(n25034), .B(n25865), .C(n25223), .D(n25864), .Y(n29170)
         );
  NAND3X1 U23685 ( .A(n29171), .B(n29172), .C(n29173), .Y(n29159) );
  NOR2X1 U23686 ( .A(n29174), .B(n29175), .Y(n29173) );
  OAI21X1 U23687 ( .A(n25040), .B(n26547), .C(n29176), .Y(n29175) );
  AOI22X1 U23688 ( .A(reg_A[71]), .B(n25135), .C(reg_A[73]), .D(n25136), .Y(
        n29176) );
  OAI21X1 U23689 ( .A(n25057), .B(n25883), .C(n29177), .Y(n29174) );
  AOI22X1 U23690 ( .A(reg_A[91]), .B(n25257), .C(reg_A[95]), .D(n25857), .Y(
        n29177) );
  NOR2X1 U23691 ( .A(n29178), .B(n29179), .Y(n29172) );
  OAI22X1 U23692 ( .A(n25331), .B(n26195), .C(n25243), .D(n25929), .Y(n29179)
         );
  OAI22X1 U23693 ( .A(n25334), .B(n26039), .C(n25336), .D(n25965), .Y(n29178)
         );
  AOI21X1 U23694 ( .A(reg_A[90]), .B(n25339), .C(n29180), .Y(n29171) );
  OAI22X1 U23695 ( .A(n25491), .B(n25881), .C(n25492), .D(n25882), .Y(n29180)
         );
  OAI21X1 U23696 ( .A(n29181), .B(n29182), .C(n25730), .Y(n29153) );
  NAND2X1 U23697 ( .A(n29183), .B(n29184), .Y(n29182) );
  AOI22X1 U23698 ( .A(reg_A[74]), .B(n25749), .C(reg_A[75]), .D(n25750), .Y(
        n29184) );
  AOI22X1 U23699 ( .A(reg_A[79]), .B(n25614), .C(reg_A[78]), .D(n25615), .Y(
        n29183) );
  NAND2X1 U23700 ( .A(n29185), .B(n29186), .Y(n29181) );
  AOI22X1 U23701 ( .A(reg_A[73]), .B(n26804), .C(reg_A[72]), .D(n26927), .Y(
        n29186) );
  AOI22X1 U23702 ( .A(reg_A[76]), .B(n26878), .C(reg_A[77]), .D(n25613), .Y(
        n29185) );
  AOI22X1 U23703 ( .A(n29084), .B(n29066), .C(n28602), .D(n29187), .Y(n29152)
         );
  OAI21X1 U23704 ( .A(n25884), .B(n26997), .C(n29137), .Y(n29066) );
  NAND2X1 U23705 ( .A(n28722), .B(n28724), .Y(n29084) );
  NAND2X1 U23706 ( .A(n25984), .B(n25932), .Y(n28724) );
  NAND2X1 U23707 ( .A(n25963), .B(n25170), .Y(n28722) );
  NOR2X1 U23708 ( .A(n29188), .B(n29189), .Y(n29120) );
  OAI21X1 U23709 ( .A(n29190), .B(n25914), .C(n29191), .Y(n29189) );
  AOI22X1 U23710 ( .A(n29192), .B(n27155), .C(n29193), .D(n29194), .Y(n29191)
         );
  NAND2X1 U23711 ( .A(n26298), .B(n26583), .Y(n29193) );
  NAND2X1 U23712 ( .A(n25980), .B(n25170), .Y(n26583) );
  NAND2X1 U23713 ( .A(reg_B[95]), .B(n25932), .Y(n26298) );
  OAI22X1 U23714 ( .A(n29195), .B(n28248), .C(n28864), .D(n28088), .Y(n29192)
         );
  INVX1 U23715 ( .A(n29000), .Y(n28864) );
  OAI21X1 U23716 ( .A(n26256), .B(n28394), .C(n28887), .Y(n29000) );
  NAND2X1 U23717 ( .A(n28296), .B(reg_A[66]), .Y(n28887) );
  INVX1 U23718 ( .A(n29196), .Y(n29195) );
  AOI22X1 U23719 ( .A(n25699), .B(n29019), .C(n29197), .D(n25932), .Y(n29190)
         );
  OAI21X1 U23720 ( .A(n29020), .B(n29198), .C(n29199), .Y(n29188) );
  AOI22X1 U23721 ( .A(n29200), .B(n29201), .C(n29202), .D(reg_B[71]), .Y(
        n29199) );
  NOR2X1 U23722 ( .A(n28213), .B(n29203), .Y(n29202) );
  NOR2X1 U23723 ( .A(n29094), .B(n25031), .Y(n29200) );
  NAND2X1 U23724 ( .A(n25170), .B(n29058), .Y(n29198) );
  MUX2X1 U23725 ( .B(n29094), .A(n29204), .S(reg_B[70]), .Y(n29058) );
  MUX2X1 U23726 ( .B(reg_A[70]), .A(reg_A[66]), .S(reg_B[69]), .Y(n29094) );
  NOR2X1 U23727 ( .A(n29205), .B(n29206), .Y(n29119) );
  OAI21X1 U23728 ( .A(n29207), .B(n26256), .C(n29208), .Y(n29206) );
  AOI22X1 U23729 ( .A(n28224), .B(n29209), .C(n29210), .D(reg_B[78]), .Y(
        n29208) );
  AND2X1 U23730 ( .A(n29211), .B(n29212), .Y(n28224) );
  AOI22X1 U23731 ( .A(n26601), .B(n26107), .C(n26602), .D(n25851), .Y(n29212)
         );
  AOI22X1 U23732 ( .A(n27012), .B(n26256), .C(n26597), .D(n25856), .Y(n29211)
         );
  OAI21X1 U23733 ( .A(n29067), .B(n28728), .C(n29213), .Y(n29205) );
  AOI22X1 U23734 ( .A(reg_A[68]), .B(n29214), .C(n29215), .D(n29216), .Y(
        n29213) );
  OAI21X1 U23735 ( .A(n29217), .B(n29218), .C(n29219), .Y(n29214) );
  INVX1 U23736 ( .A(n29220), .Y(n29219) );
  NAND2X1 U23737 ( .A(n29026), .B(n29221), .Y(n29218) );
  OR2X1 U23738 ( .A(n29222), .B(n29223), .Y(result[6]) );
  NAND3X1 U23739 ( .A(n29224), .B(n29225), .C(n29226), .Y(n29223) );
  NOR2X1 U23740 ( .A(n29227), .B(n29228), .Y(n29226) );
  OAI21X1 U23741 ( .A(n29229), .B(n25087), .C(n26754), .Y(n29228) );
  AND2X1 U23742 ( .A(n29230), .B(n29231), .Y(n29229) );
  AOI21X1 U23743 ( .A(n28023), .B(n29232), .C(n29233), .Y(n29231) );
  OAI21X1 U23744 ( .A(n29234), .B(n29235), .C(n29236), .Y(n29233) );
  OAI21X1 U23745 ( .A(n29237), .B(n29238), .C(n25044), .Y(n29236) );
  OAI22X1 U23746 ( .A(n29239), .B(n25106), .C(n29240), .D(n25099), .Y(n29238)
         );
  OAI21X1 U23747 ( .A(n29241), .B(n28033), .C(n29242), .Y(n29237) );
  AOI22X1 U23748 ( .A(n25110), .B(n29243), .C(reg_B[27]), .D(n29244), .Y(
        n29242) );
  AOI22X1 U23749 ( .A(n29245), .B(n29246), .C(n28038), .D(n29247), .Y(n29230)
         );
  OAI21X1 U23750 ( .A(n29248), .B(n25177), .C(n29249), .Y(n29227) );
  AOI22X1 U23751 ( .A(reg_A[7]), .B(n28923), .C(reg_A[2]), .D(n29250), .Y(
        n29249) );
  AOI21X1 U23752 ( .A(n25730), .B(n29251), .C(n29252), .Y(n29225) );
  OAI21X1 U23753 ( .A(n27994), .B(n25189), .C(n29253), .Y(n29252) );
  OAI21X1 U23754 ( .A(n29127), .B(n29254), .C(reg_A[0]), .Y(n29253) );
  OAI22X1 U23755 ( .A(n27438), .B(n29255), .C(n29256), .D(n28057), .Y(n29254)
         );
  AOI22X1 U23756 ( .A(n29257), .B(n26267), .C(reg_A[4]), .D(n29258), .Y(n27994) );
  INVX1 U23757 ( .A(n26727), .Y(n29258) );
  NAND3X1 U23758 ( .A(n29259), .B(n29260), .C(n29261), .Y(n29251) );
  NOR2X1 U23759 ( .A(n29262), .B(n29263), .Y(n29261) );
  OAI22X1 U23760 ( .A(n26936), .B(n25206), .C(n25745), .D(n25255), .Y(n29263)
         );
  OAI22X1 U23761 ( .A(n26701), .B(n25746), .C(n25146), .D(n25747), .Y(n29262)
         );
  AOI22X1 U23762 ( .A(reg_A[10]), .B(n25749), .C(reg_A[11]), .D(n25750), .Y(
        n29260) );
  AOI22X1 U23763 ( .A(n25614), .B(reg_A[15]), .C(n25615), .D(reg_A[14]), .Y(
        n29259) );
  AOI21X1 U23764 ( .A(reg_A[3]), .B(n29155), .C(n29264), .Y(n29224) );
  OAI21X1 U23765 ( .A(n29157), .B(n29265), .C(n29266), .Y(n29264) );
  OAI21X1 U23766 ( .A(n29267), .B(n29268), .C(n25310), .Y(n29266) );
  NAND3X1 U23767 ( .A(n29269), .B(n29270), .C(n29271), .Y(n29268) );
  NOR2X1 U23768 ( .A(n29272), .B(n29273), .Y(n29271) );
  OAI21X1 U23769 ( .A(n26677), .B(n25043), .C(n29274), .Y(n29273) );
  AOI22X1 U23770 ( .A(n25635), .B(reg_A[18]), .C(n25325), .D(reg_A[19]), .Y(
        n29274) );
  OAI21X1 U23771 ( .A(n25065), .B(n25232), .C(n29275), .Y(n29272) );
  AOI22X1 U23772 ( .A(n25637), .B(reg_A[16]), .C(n25234), .D(reg_A[20]), .Y(
        n29275) );
  NOR2X1 U23773 ( .A(n29276), .B(n29277), .Y(n29270) );
  OAI22X1 U23774 ( .A(n27967), .B(n26703), .C(n25147), .D(n26431), .Y(n29277)
         );
  OAI22X1 U23775 ( .A(n25030), .B(n25206), .C(n25255), .D(n25131), .Y(n29276)
         );
  AOI21X1 U23776 ( .A(n25222), .B(reg_A[17]), .C(n29278), .Y(n29269) );
  OAI22X1 U23777 ( .A(n25208), .B(n25467), .C(n29279), .D(n25223), .Y(n29278)
         );
  NAND3X1 U23778 ( .A(n29280), .B(n29281), .C(n29282), .Y(n29267) );
  NOR2X1 U23779 ( .A(n29283), .B(n29284), .Y(n29282) );
  OAI21X1 U23780 ( .A(n26701), .B(n25133), .C(n29285), .Y(n29284) );
  AOI22X1 U23781 ( .A(n25135), .B(reg_A[7]), .C(n25136), .D(reg_A[9]), .Y(
        n29285) );
  OAI21X1 U23782 ( .A(n29286), .B(n25320), .C(n29287), .Y(n29283) );
  AOI22X1 U23783 ( .A(n25257), .B(reg_A[27]), .C(n25857), .D(reg_A[31]), .Y(
        n29287) );
  NOR2X1 U23784 ( .A(n29288), .B(n29289), .Y(n29281) );
  OAI22X1 U23785 ( .A(n25331), .B(n27962), .C(n27960), .D(n25243), .Y(n29289)
         );
  OAI22X1 U23786 ( .A(n25334), .B(n25230), .C(n25336), .D(n26714), .Y(n29288)
         );
  AOI21X1 U23787 ( .A(n25339), .B(reg_A[26]), .C(n29290), .Y(n29280) );
  OAI22X1 U23788 ( .A(n25239), .B(n25491), .C(n25244), .D(n25492), .Y(n29290)
         );
  INVX1 U23789 ( .A(n29291), .Y(n29157) );
  NAND3X1 U23790 ( .A(n29292), .B(n29293), .C(n29294), .Y(n29222) );
  NOR2X1 U23791 ( .A(n29295), .B(n29296), .Y(n29294) );
  OAI21X1 U23792 ( .A(n25198), .B(n29297), .C(n29298), .Y(n29296) );
  AOI22X1 U23793 ( .A(n29299), .B(n25699), .C(n29300), .D(n27155), .Y(n29298)
         );
  OAI22X1 U23794 ( .A(n29301), .B(n29302), .C(n29303), .D(n26692), .Y(n29300)
         );
  INVX1 U23795 ( .A(n25160), .Y(n29303) );
  OAI21X1 U23796 ( .A(n29304), .B(n26677), .C(n25195), .Y(n25160) );
  NAND2X1 U23797 ( .A(reg_A[2]), .B(n26691), .Y(n25195) );
  NOR2X1 U23798 ( .A(n27979), .B(n29305), .Y(n29299) );
  AOI22X1 U23799 ( .A(n25156), .B(n26760), .C(n29306), .D(reg_B[31]), .Y(
        n29297) );
  INVX1 U23800 ( .A(n25263), .Y(n26760) );
  AOI21X1 U23801 ( .A(reg_A[2]), .B(n25101), .C(n29307), .Y(n25263) );
  OAI21X1 U23802 ( .A(n28041), .B(n29308), .C(n29309), .Y(n29295) );
  AOI21X1 U23803 ( .A(n29310), .B(n27986), .C(n29311), .Y(n29309) );
  INVX1 U23804 ( .A(n29312), .Y(n29311) );
  NOR2X1 U23805 ( .A(n29313), .B(n25031), .Y(n29310) );
  NAND2X1 U23806 ( .A(n29314), .B(n29315), .Y(n29308) );
  AOI21X1 U23807 ( .A(n29316), .B(n29317), .C(n29318), .Y(n29293) );
  OAI21X1 U23808 ( .A(n28049), .B(n29319), .C(n29320), .Y(n29318) );
  OAI21X1 U23809 ( .A(n29321), .B(n29220), .C(reg_A[4]), .Y(n29320) );
  INVX1 U23810 ( .A(n29322), .Y(n29321) );
  MUX2X1 U23811 ( .B(n28010), .A(n29323), .S(reg_B[6]), .Y(n28049) );
  INVX1 U23812 ( .A(n29313), .Y(n28010) );
  MUX2X1 U23813 ( .B(reg_A[6]), .A(reg_A[2]), .S(reg_B[5]), .Y(n29313) );
  AOI22X1 U23814 ( .A(n29324), .B(n29209), .C(reg_A[6]), .D(n29325), .Y(n29292) );
  NAND3X1 U23815 ( .A(n29326), .B(n29327), .C(n29328), .Y(result[69]) );
  NOR2X1 U23816 ( .A(n29329), .B(n29330), .Y(n29328) );
  NAND3X1 U23817 ( .A(n29331), .B(n29125), .C(n29332), .Y(n29330) );
  AOI21X1 U23818 ( .A(n25730), .B(n29333), .C(n29334), .Y(n29332) );
  OAI21X1 U23819 ( .A(n29335), .B(n26919), .C(n29336), .Y(n29334) );
  OAI21X1 U23820 ( .A(n29337), .B(n29338), .C(n27358), .Y(n29336) );
  OAI21X1 U23821 ( .A(n29339), .B(n25856), .C(n29340), .Y(n29338) );
  AOI22X1 U23822 ( .A(reg_A[65]), .B(n25650), .C(reg_A[68]), .D(n29341), .Y(
        n29340) );
  NAND2X1 U23823 ( .A(n29342), .B(n29343), .Y(n29337) );
  AOI22X1 U23824 ( .A(n29344), .B(n29345), .C(reg_A[66]), .D(n29346), .Y(
        n29343) );
  INVX1 U23825 ( .A(n29050), .Y(n29344) );
  NAND2X1 U23826 ( .A(n29347), .B(n29348), .Y(n29050) );
  AOI22X1 U23827 ( .A(n26292), .B(n25855), .C(n26293), .D(n25856), .Y(n29348)
         );
  AOI22X1 U23828 ( .A(n26294), .B(n25853), .C(n26295), .D(n26107), .Y(n29347)
         );
  AOI22X1 U23829 ( .A(reg_A[67]), .B(n29349), .C(reg_A[64]), .D(n29350), .Y(
        n29342) );
  INVX1 U23830 ( .A(n29351), .Y(n29335) );
  NAND3X1 U23831 ( .A(n29352), .B(n29353), .C(n29354), .Y(n29333) );
  NOR2X1 U23832 ( .A(n29355), .B(n29356), .Y(n29354) );
  OAI21X1 U23833 ( .A(n26801), .B(n26439), .C(n29357), .Y(n29356) );
  AOI22X1 U23834 ( .A(reg_A[75]), .B(n26878), .C(reg_A[76]), .D(n25613), .Y(
        n29357) );
  OAI21X1 U23835 ( .A(n25062), .B(n26101), .C(n29358), .Y(n29355) );
  AOI22X1 U23836 ( .A(reg_A[70]), .B(n26803), .C(reg_A[72]), .D(n26804), .Y(
        n29358) );
  AOI21X1 U23837 ( .A(reg_A[77]), .B(n25615), .C(n29359), .Y(n29353) );
  OAI22X1 U23838 ( .A(n27253), .B(n25865), .C(n26800), .D(n26438), .Y(n29359)
         );
  AOI22X1 U23839 ( .A(reg_A[79]), .B(n25607), .C(reg_A[69]), .D(n26924), .Y(
        n29352) );
  INVX1 U23840 ( .A(n29009), .Y(n29125) );
  OAI21X1 U23841 ( .A(n25032), .B(n28882), .C(n29360), .Y(n29009) );
  OAI21X1 U23842 ( .A(n27537), .B(n26974), .C(n25932), .Y(n29360) );
  INVX1 U23843 ( .A(n28605), .Y(n26974) );
  NAND2X1 U23844 ( .A(reg_A[64]), .B(reg_B[92]), .Y(n28605) );
  INVX1 U23845 ( .A(n27664), .Y(n27537) );
  NAND2X1 U23846 ( .A(reg_A[64]), .B(reg_B[91]), .Y(n27664) );
  NAND2X1 U23847 ( .A(reg_B[76]), .B(reg_A[64]), .Y(n28882) );
  AOI22X1 U23848 ( .A(reg_A[70]), .B(n27402), .C(reg_A[71]), .D(n29361), .Y(
        n29331) );
  NAND3X1 U23849 ( .A(n29362), .B(n29363), .C(n29364), .Y(n29329) );
  INVX1 U23850 ( .A(n29365), .Y(n29364) );
  OAI21X1 U23851 ( .A(n29366), .B(n26107), .C(n29367), .Y(n29365) );
  AOI22X1 U23852 ( .A(n29187), .B(n28191), .C(reg_A[64]), .D(n29368), .Y(
        n29367) );
  OAI22X1 U23853 ( .A(n29369), .B(n26147), .C(n26107), .D(n28215), .Y(n29187)
         );
  OAI21X1 U23854 ( .A(n29370), .B(n29371), .C(n25310), .Y(n29363) );
  NAND3X1 U23855 ( .A(n29372), .B(n29373), .C(n29374), .Y(n29371) );
  NOR2X1 U23856 ( .A(n29375), .B(n29376), .Y(n29374) );
  OAI21X1 U23857 ( .A(n25043), .B(n25856), .C(n29377), .Y(n29376) );
  AOI22X1 U23858 ( .A(reg_A[81]), .B(n25635), .C(reg_A[82]), .D(n25325), .Y(
        n29377) );
  OAI21X1 U23859 ( .A(n25065), .B(n26230), .C(n29378), .Y(n29375) );
  AOI22X1 U23860 ( .A(reg_A[79]), .B(n25637), .C(reg_A[83]), .D(n25234), .Y(
        n29378) );
  NOR2X1 U23861 ( .A(n29379), .B(n29380), .Y(n29373) );
  OAI22X1 U23862 ( .A(n25028), .B(n26438), .C(n26431), .D(n26439), .Y(n29380)
         );
  OAI22X1 U23863 ( .A(n25030), .B(n25863), .C(n25131), .D(n26103), .Y(n29379)
         );
  AOI21X1 U23864 ( .A(reg_A[80]), .B(n25222), .C(n29381), .Y(n29372) );
  OAI22X1 U23865 ( .A(n25034), .B(n26286), .C(n25223), .D(n25865), .Y(n29381)
         );
  NAND3X1 U23866 ( .A(n29382), .B(n29383), .C(n29384), .Y(n29370) );
  NOR2X1 U23867 ( .A(n29385), .B(n29386), .Y(n29384) );
  OAI21X1 U23868 ( .A(n25238), .B(n25929), .C(n29387), .Y(n29386) );
  AOI22X1 U23869 ( .A(reg_A[91]), .B(n25242), .C(reg_A[92]), .D(n25338), .Y(
        n29387) );
  NAND2X1 U23870 ( .A(n29388), .B(n29389), .Y(n29385) );
  AOI22X1 U23871 ( .A(reg_A[86]), .B(n25246), .C(reg_A[85]), .D(n25247), .Y(
        n29389) );
  AOI22X1 U23872 ( .A(reg_A[88]), .B(n25487), .C(reg_A[87]), .D(n25241), .Y(
        n29388) );
  NOR2X1 U23873 ( .A(n29390), .B(n29391), .Y(n29383) );
  OAI22X1 U23874 ( .A(n25316), .B(n25873), .C(n25320), .D(n25881), .Y(n29391)
         );
  OAI22X1 U23875 ( .A(n25322), .B(n25883), .C(n26719), .D(n26068), .Y(n29390)
         );
  AOI21X1 U23876 ( .A(reg_A[71]), .B(n25252), .C(n29392), .Y(n29382) );
  OAI22X1 U23877 ( .A(n25041), .B(n26547), .C(n25042), .D(n26256), .Y(n29392)
         );
  AOI22X1 U23878 ( .A(reg_A[69]), .B(n29393), .C(n29394), .D(reg_A[67]), .Y(
        n29362) );
  NOR2X1 U23879 ( .A(n29395), .B(n29396), .Y(n29327) );
  OAI21X1 U23880 ( .A(n25855), .B(n29397), .C(n29398), .Y(n29396) );
  AOI22X1 U23881 ( .A(n29399), .B(n29400), .C(n29057), .D(n29401), .Y(n29398)
         );
  INVX1 U23882 ( .A(n29203), .Y(n29400) );
  MUX2X1 U23883 ( .B(n29025), .A(n29402), .S(reg_B[70]), .Y(n29203) );
  NOR2X1 U23884 ( .A(reg_B[69]), .B(n25851), .Y(n29402) );
  INVX1 U23885 ( .A(n29403), .Y(n29025) );
  NAND3X1 U23886 ( .A(n29404), .B(n29405), .C(n29406), .Y(n29395) );
  AOI22X1 U23887 ( .A(n29407), .B(n29098), .C(n29408), .D(n29196), .Y(n29406)
         );
  OAI22X1 U23888 ( .A(n25851), .B(n28879), .C(reg_B[78]), .D(n28997), .Y(
        n29196) );
  INVX1 U23889 ( .A(n29027), .Y(n28997) );
  OAI22X1 U23890 ( .A(n25856), .B(n28394), .C(n25855), .D(n28483), .Y(n29027)
         );
  OAI21X1 U23891 ( .A(reg_B[79]), .B(n25794), .C(n29409), .Y(n29408) );
  MUX2X1 U23892 ( .B(n29403), .A(n29410), .S(reg_B[71]), .Y(n29098) );
  MUX2X1 U23893 ( .B(reg_A[68]), .A(reg_A[64]), .S(reg_B[69]), .Y(n29410) );
  MUX2X1 U23894 ( .B(reg_A[69]), .A(reg_A[65]), .S(reg_B[69]), .Y(n29403) );
  NOR2X1 U23895 ( .A(reg_B[70]), .B(n25031), .Y(n29407) );
  OAI21X1 U23896 ( .A(n26125), .B(n26050), .C(n29194), .Y(n29405) );
  OAI22X1 U23897 ( .A(n29065), .B(reg_B[94]), .C(n25851), .D(n29411), .Y(
        n29194) );
  INVX1 U23898 ( .A(n29412), .Y(n29411) );
  INVX1 U23899 ( .A(n28952), .Y(n29065) );
  OAI21X1 U23900 ( .A(n25855), .B(n26997), .C(n29413), .Y(n28952) );
  INVX1 U23901 ( .A(n26950), .Y(n26050) );
  INVX1 U23902 ( .A(n25886), .Y(n26125) );
  NAND2X1 U23903 ( .A(n25932), .B(n25976), .Y(n25886) );
  OAI21X1 U23904 ( .A(n29215), .B(n29414), .C(n29216), .Y(n29404) );
  INVX1 U23905 ( .A(n29217), .Y(n29216) );
  MUX2X1 U23906 ( .B(n29415), .A(n29416), .S(reg_B[71]), .Y(n29414) );
  NAND2X1 U23907 ( .A(reg_A[67]), .B(n29026), .Y(n29415) );
  NOR2X1 U23908 ( .A(n29417), .B(n29418), .Y(n29326) );
  NAND3X1 U23909 ( .A(n29419), .B(n29420), .C(n29421), .Y(n29418) );
  OAI21X1 U23910 ( .A(n29422), .B(n29423), .C(n25932), .Y(n29421) );
  OAI22X1 U23911 ( .A(n26168), .B(n29068), .C(n25984), .D(n29067), .Y(n29423)
         );
  NAND2X1 U23912 ( .A(reg_A[64]), .B(reg_B[93]), .Y(n29067) );
  NOR2X1 U23913 ( .A(n26169), .B(n29424), .Y(n29422) );
  INVX1 U23914 ( .A(n29425), .Y(n29420) );
  AOI21X1 U23915 ( .A(n29426), .B(n29427), .C(n26996), .Y(n29425) );
  AOI22X1 U23916 ( .A(n28827), .B(n28826), .C(n28825), .D(n28930), .Y(n29427)
         );
  AOI22X1 U23917 ( .A(n28340), .B(n26307), .C(n27401), .D(reg_B[91]), .Y(
        n29426) );
  OAI21X1 U23918 ( .A(n26807), .B(n26069), .C(n29428), .Y(n27401) );
  AOI22X1 U23919 ( .A(n26275), .B(n28461), .C(n25988), .D(n28460), .Y(n29428)
         );
  INVX1 U23920 ( .A(n28830), .Y(n26807) );
  OAI21X1 U23921 ( .A(n29429), .B(n29430), .C(n25382), .Y(n29419) );
  OAI22X1 U23922 ( .A(n29431), .B(n29102), .C(n28819), .D(n29149), .Y(n29430)
         );
  INVX1 U23923 ( .A(n29432), .Y(n29429) );
  AOI22X1 U23924 ( .A(n29433), .B(n29434), .C(n28817), .D(n29134), .Y(n29432)
         );
  OAI21X1 U23925 ( .A(n29435), .B(n27020), .C(n29436), .Y(n29417) );
  AOI22X1 U23926 ( .A(n29210), .B(n28088), .C(reg_A[66]), .D(n29437), .Y(
        n29436) );
  OAI21X1 U23927 ( .A(n28130), .B(n28879), .C(n29438), .Y(n29437) );
  NOR2X1 U23928 ( .A(n29439), .B(n29069), .Y(n29438) );
  NOR2X1 U23929 ( .A(n28215), .B(n28208), .Y(n29069) );
  NAND2X1 U23930 ( .A(n28297), .B(n25188), .Y(n28215) );
  INVX1 U23931 ( .A(n29055), .Y(n29210) );
  NAND3X1 U23932 ( .A(reg_A[64]), .B(n25188), .C(reg_B[77]), .Y(n29055) );
  NAND3X1 U23933 ( .A(n29440), .B(n29441), .C(n29442), .Y(result[68]) );
  NOR2X1 U23934 ( .A(n29443), .B(n29444), .Y(n29442) );
  NAND3X1 U23935 ( .A(n29445), .B(n29446), .C(n29447), .Y(n29444) );
  AOI22X1 U23936 ( .A(n25372), .B(n29448), .C(n26116), .D(n29449), .Y(n29447)
         );
  INVX1 U23937 ( .A(n27020), .Y(n26116) );
  NAND3X1 U23938 ( .A(n29450), .B(n29451), .C(n29452), .Y(n29448) );
  NOR2X1 U23939 ( .A(n29453), .B(n29454), .Y(n29452) );
  OAI21X1 U23940 ( .A(n29424), .B(n29455), .C(n29456), .Y(n29454) );
  NAND3X1 U23941 ( .A(reg_B[71]), .B(n25589), .C(n29457), .Y(n29456) );
  NAND2X1 U23942 ( .A(n26276), .B(n25044), .Y(n29455) );
  OAI21X1 U23943 ( .A(n28248), .B(n29458), .C(n29459), .Y(n29453) );
  NAND2X1 U23944 ( .A(n25604), .B(n29460), .Y(n29458) );
  AOI22X1 U23945 ( .A(n25980), .B(n29449), .C(n29197), .D(n25963), .Y(n29451)
         );
  INVX1 U23946 ( .A(n27053), .Y(n25980) );
  NAND2X1 U23947 ( .A(reg_B[95]), .B(n25044), .Y(n27053) );
  AOI22X1 U23948 ( .A(reg_A[66]), .B(n29461), .C(reg_A[68]), .D(n29462), .Y(
        n29450) );
  OAI21X1 U23949 ( .A(n29463), .B(n29464), .C(n27358), .Y(n29446) );
  OAI21X1 U23950 ( .A(n25598), .B(n25884), .C(n29465), .Y(n29464) );
  AOI22X1 U23951 ( .A(reg_A[65]), .B(n27740), .C(reg_A[68]), .D(n29466), .Y(
        n29465) );
  OAI21X1 U23952 ( .A(n29467), .B(n25851), .C(n29468), .Y(n29463) );
  AOI22X1 U23953 ( .A(reg_A[64]), .B(n29469), .C(n28573), .D(n29470), .Y(
        n29468) );
  INVX1 U23954 ( .A(n27449), .Y(n29470) );
  AND2X1 U23955 ( .A(n29471), .B(n29472), .Y(n28573) );
  AOI22X1 U23956 ( .A(n26601), .B(n25884), .C(n26602), .D(n25855), .Y(n29472)
         );
  AOI22X1 U23957 ( .A(n27012), .B(n26107), .C(n26597), .D(n25851), .Y(n29471)
         );
  NAND2X1 U23958 ( .A(n29473), .B(n27448), .Y(n29469) );
  AOI22X1 U23959 ( .A(reg_A[69]), .B(n28923), .C(n28083), .D(n29474), .Y(
        n29445) );
  INVX1 U23960 ( .A(n26919), .Y(n28083) );
  NAND2X1 U23961 ( .A(n26480), .B(n26057), .Y(n26919) );
  NAND3X1 U23962 ( .A(n29475), .B(n29476), .C(n29477), .Y(n29443) );
  AOI22X1 U23963 ( .A(reg_A[71]), .B(n26739), .C(reg_A[70]), .D(n26783), .Y(
        n29477) );
  OAI21X1 U23964 ( .A(n29478), .B(n29479), .C(n25310), .Y(n29476) );
  NAND3X1 U23965 ( .A(n29480), .B(n29481), .C(n29482), .Y(n29479) );
  NOR2X1 U23966 ( .A(n29483), .B(n29484), .Y(n29482) );
  OAI21X1 U23967 ( .A(n25034), .B(n25863), .C(n29485), .Y(n29484) );
  AOI22X1 U23968 ( .A(reg_A[73]), .B(n25123), .C(reg_A[77]), .D(n25629), .Y(
        n29485) );
  NAND2X1 U23969 ( .A(n29486), .B(n29487), .Y(n29483) );
  AOI22X1 U23970 ( .A(reg_A[70]), .B(n25252), .C(reg_A[74]), .D(n25253), .Y(
        n29487) );
  AOI22X1 U23971 ( .A(reg_A[75]), .B(n25628), .C(reg_A[72]), .D(n25068), .Y(
        n29486) );
  NOR2X1 U23972 ( .A(n29488), .B(n29489), .Y(n29481) );
  OAI22X1 U23973 ( .A(n25065), .B(n25875), .C(n25035), .D(n25874), .Y(n29489)
         );
  OAI22X1 U23974 ( .A(n25036), .B(n25865), .C(n25473), .D(n25864), .Y(n29488)
         );
  AOI21X1 U23975 ( .A(reg_A[68]), .B(n25125), .C(n29490), .Y(n29480) );
  OAI22X1 U23976 ( .A(n25039), .B(n26094), .C(n25231), .D(n25584), .Y(n29490)
         );
  NAND3X1 U23977 ( .A(n29491), .B(n29492), .C(n29493), .Y(n29478) );
  NOR2X1 U23978 ( .A(n29494), .B(n29495), .Y(n29493) );
  OAI21X1 U23979 ( .A(n25238), .B(n26195), .C(n29496), .Y(n29495) );
  AOI22X1 U23980 ( .A(reg_A[90]), .B(n25242), .C(reg_A[91]), .D(n25338), .Y(
        n29496) );
  NAND2X1 U23981 ( .A(n29497), .B(n29498), .Y(n29494) );
  AOI22X1 U23982 ( .A(reg_A[85]), .B(n25246), .C(reg_A[84]), .D(n25247), .Y(
        n29498) );
  AOI22X1 U23983 ( .A(reg_A[87]), .B(n25487), .C(reg_A[86]), .D(n25241), .Y(
        n29497) );
  NOR2X1 U23984 ( .A(n29499), .B(n29500), .Y(n29492) );
  OAI22X1 U23985 ( .A(n25318), .B(n25873), .C(n25320), .D(n25882), .Y(n29500)
         );
  OAI22X1 U23986 ( .A(n25322), .B(n25881), .C(n26719), .D(n25929), .Y(n29499)
         );
  AOI21X1 U23987 ( .A(reg_A[71]), .B(n25136), .C(n29501), .Y(n29491) );
  OAI22X1 U23988 ( .A(n25042), .B(n25856), .C(n25316), .D(n25883), .Y(n29501)
         );
  AOI22X1 U23989 ( .A(n29502), .B(reg_A[67]), .C(n29439), .D(reg_A[65]), .Y(
        n29475) );
  NOR2X1 U23990 ( .A(n29503), .B(n29504), .Y(n29441) );
  OAI21X1 U23991 ( .A(n29505), .B(n28130), .C(n29506), .Y(n29504) );
  AOI22X1 U23992 ( .A(n29457), .B(n29057), .C(n29507), .D(reg_A[64]), .Y(
        n29506) );
  OAI21X1 U23993 ( .A(n29508), .B(n29509), .C(n29510), .Y(n29503) );
  AOI22X1 U23994 ( .A(n29511), .B(n28288), .C(reg_A[66]), .D(n29512), .Y(
        n29510) );
  OAI21X1 U23995 ( .A(n29409), .B(n28879), .C(n29513), .Y(n29512) );
  NOR2X1 U23996 ( .A(reg_B[78]), .B(n29369), .Y(n29511) );
  INVX1 U23997 ( .A(n29023), .Y(n29369) );
  OAI22X1 U23998 ( .A(n26107), .B(n28394), .C(n25853), .D(n28483), .Y(n29023)
         );
  INVX1 U23999 ( .A(n29401), .Y(n29508) );
  MUX2X1 U24000 ( .B(n29204), .A(n29416), .S(reg_B[70]), .Y(n29401) );
  AOI21X1 U24001 ( .A(n29026), .B(reg_A[68]), .C(n29215), .Y(n29204) );
  NOR2X1 U24002 ( .A(n29026), .B(n25853), .Y(n29215) );
  NOR2X1 U24003 ( .A(n29514), .B(n29515), .Y(n29440) );
  OAI21X1 U24004 ( .A(n29435), .B(n26950), .C(n29516), .Y(n29515) );
  OAI21X1 U24005 ( .A(n29517), .B(n29518), .C(n25730), .Y(n29516) );
  NAND2X1 U24006 ( .A(n29519), .B(n29520), .Y(n29518) );
  AOI22X1 U24007 ( .A(reg_A[77]), .B(n25614), .C(reg_A[76]), .D(n25615), .Y(
        n29520) );
  AOI22X1 U24008 ( .A(reg_A[79]), .B(n25616), .C(reg_A[78]), .D(n25607), .Y(
        n29519) );
  NAND2X1 U24009 ( .A(n29521), .B(n29522), .Y(n29517) );
  AOI22X1 U24010 ( .A(reg_A[74]), .B(n26878), .C(reg_A[75]), .D(n25613), .Y(
        n29522) );
  AOI22X1 U24011 ( .A(reg_A[72]), .B(n25749), .C(reg_A[73]), .D(n25750), .Y(
        n29521) );
  MUX2X1 U24012 ( .B(n29019), .A(n29523), .S(reg_B[94]), .Y(n29435) );
  OAI21X1 U24013 ( .A(n25853), .B(n26997), .C(n29068), .Y(n29019) );
  NAND3X1 U24014 ( .A(n29524), .B(n29525), .C(n29526), .Y(n29514) );
  INVX1 U24015 ( .A(n29527), .Y(n29526) );
  AOI21X1 U24016 ( .A(n29528), .B(n29529), .C(n25087), .Y(n29527) );
  AOI22X1 U24017 ( .A(n29530), .B(n29146), .C(n29531), .D(n29434), .Y(n29529)
         );
  INVX1 U24018 ( .A(n29102), .Y(n29146) );
  AOI22X1 U24019 ( .A(n28924), .B(n29134), .C(n28934), .D(n28103), .Y(n29528)
         );
  OR2X1 U24020 ( .A(n26107), .B(n29532), .Y(n29525) );
  OAI21X1 U24021 ( .A(n29533), .B(n29534), .C(n26480), .Y(n29524) );
  OAI22X1 U24022 ( .A(n28932), .B(n26997), .C(n28561), .D(n25964), .Y(n29534)
         );
  INVX1 U24023 ( .A(n29535), .Y(n28932) );
  OAI22X1 U24024 ( .A(n28507), .B(n28093), .C(n29536), .D(n25895), .Y(n29533)
         );
  INVX1 U24025 ( .A(n27499), .Y(n29536) );
  OAI21X1 U24026 ( .A(n28510), .B(n26069), .C(n29537), .Y(n27499) );
  AOI22X1 U24027 ( .A(n26275), .B(n28509), .C(n25988), .D(n26992), .Y(n29537)
         );
  INVX1 U24028 ( .A(n26915), .Y(n28510) );
  INVX1 U24029 ( .A(n29538), .Y(n28507) );
  NAND3X1 U24030 ( .A(n29539), .B(n29540), .C(n29541), .Y(result[67]) );
  NOR2X1 U24031 ( .A(n29542), .B(n29543), .Y(n29541) );
  NAND2X1 U24032 ( .A(n29544), .B(n29545), .Y(n29543) );
  AOI22X1 U24033 ( .A(n29546), .B(reg_A[67]), .C(reg_A[68]), .D(n27402), .Y(
        n29545) );
  AOI22X1 U24034 ( .A(reg_A[70]), .B(n29547), .C(reg_A[69]), .D(n29361), .Y(
        n29544) );
  NAND2X1 U24035 ( .A(n29548), .B(n29549), .Y(n29542) );
  AOI21X1 U24036 ( .A(n28288), .B(n29460), .C(n29550), .Y(n29549) );
  OAI21X1 U24037 ( .A(n29551), .B(n26950), .C(n29552), .Y(n29550) );
  OAI21X1 U24038 ( .A(n29553), .B(n29554), .C(n25730), .Y(n29552) );
  OR2X1 U24039 ( .A(n29555), .B(n29556), .Y(n29554) );
  OAI21X1 U24040 ( .A(n25060), .B(n25851), .C(n29557), .Y(n29556) );
  AOI22X1 U24041 ( .A(reg_A[77]), .B(n25607), .C(reg_A[79]), .D(n25609), .Y(
        n29557) );
  OAI21X1 U24042 ( .A(n29558), .B(n25865), .C(n29559), .Y(n29555) );
  AOI22X1 U24043 ( .A(reg_A[76]), .B(n25614), .C(reg_A[75]), .D(n25615), .Y(
        n29559) );
  NAND3X1 U24044 ( .A(n29560), .B(n29561), .C(n29562), .Y(n29553) );
  AOI21X1 U24045 ( .A(reg_A[72]), .B(n25750), .C(n29563), .Y(n29562) );
  OAI22X1 U24046 ( .A(n26801), .B(n26101), .C(n26936), .D(n26438), .Y(n29563)
         );
  AOI22X1 U24047 ( .A(reg_A[68]), .B(n26803), .C(reg_A[70]), .D(n26804), .Y(
        n29561) );
  AOI22X1 U24048 ( .A(reg_A[69]), .B(n26927), .C(reg_A[73]), .D(n26878), .Y(
        n29560) );
  INVX1 U24049 ( .A(n29409), .Y(n28288) );
  AOI22X1 U24050 ( .A(n29564), .B(n29565), .C(reg_A[71]), .D(n25722), .Y(
        n29548) );
  OAI21X1 U24051 ( .A(n29566), .B(n25851), .C(n29567), .Y(n29564) );
  AOI22X1 U24052 ( .A(reg_A[66]), .B(n29568), .C(reg_A[65]), .D(n29569), .Y(
        n29567) );
  NOR2X1 U24053 ( .A(n29570), .B(n29571), .Y(n29540) );
  OAI21X1 U24054 ( .A(n29572), .B(n27020), .C(n29573), .Y(n29571) );
  OAI21X1 U24055 ( .A(n29574), .B(n29575), .C(n25382), .Y(n29573) );
  NAND2X1 U24056 ( .A(n29576), .B(n29577), .Y(n29575) );
  AOI22X1 U24057 ( .A(n29134), .B(n29105), .C(reg_A[68]), .D(n29578), .Y(
        n29577) );
  NAND2X1 U24058 ( .A(n29579), .B(n29580), .Y(n29105) );
  AOI22X1 U24059 ( .A(n28602), .B(reg_A[73]), .C(n28191), .D(reg_A[72]), .Y(
        n29580) );
  AOI22X1 U24060 ( .A(n28245), .B(reg_A[74]), .C(n28446), .D(reg_A[71]), .Y(
        n29579) );
  AOI22X1 U24061 ( .A(reg_A[69]), .B(n29461), .C(reg_A[70]), .D(n29581), .Y(
        n29576) );
  NAND3X1 U24062 ( .A(n29582), .B(n29583), .C(n29584), .Y(n29574) );
  AOI22X1 U24063 ( .A(reg_A[67]), .B(n29585), .C(n28609), .D(n25963), .Y(
        n29584) );
  OAI21X1 U24064 ( .A(n29586), .B(n29587), .C(n25044), .Y(n29583) );
  OAI21X1 U24065 ( .A(n28660), .B(n25964), .C(n29588), .Y(n29587) );
  AOI22X1 U24066 ( .A(reg_B[91]), .B(n27594), .C(n28826), .D(n28084), .Y(
        n29588) );
  NAND2X1 U24067 ( .A(n29589), .B(n29590), .Y(n28084) );
  AOI22X1 U24068 ( .A(n26276), .B(reg_A[81]), .C(n26149), .D(reg_A[82]), .Y(
        n29590) );
  AOI22X1 U24069 ( .A(n26148), .B(reg_A[80]), .C(reg_A[79]), .D(n25984), .Y(
        n29589) );
  OAI21X1 U24070 ( .A(n26063), .B(n26479), .C(n29591), .Y(n27594) );
  AOI22X1 U24071 ( .A(n26275), .B(n29117), .C(n26274), .D(n28597), .Y(n29591)
         );
  NAND2X1 U24072 ( .A(n29592), .B(n29593), .Y(n28597) );
  AOI22X1 U24073 ( .A(n26276), .B(reg_A[89]), .C(n26149), .D(reg_A[90]), .Y(
        n29593) );
  AOI22X1 U24074 ( .A(n26148), .B(reg_A[88]), .C(reg_A[87]), .D(n25984), .Y(
        n29592) );
  NAND2X1 U24075 ( .A(n29594), .B(n29595), .Y(n29117) );
  AOI22X1 U24076 ( .A(n26276), .B(reg_A[85]), .C(n26149), .D(reg_A[86]), .Y(
        n29595) );
  AOI22X1 U24077 ( .A(n26148), .B(reg_A[84]), .C(reg_A[83]), .D(n25984), .Y(
        n29594) );
  MUX2X1 U24078 ( .B(n25902), .A(n29116), .S(n26197), .Y(n26479) );
  NAND2X1 U24079 ( .A(n29596), .B(n29597), .Y(n29116) );
  AOI22X1 U24080 ( .A(n26276), .B(reg_A[93]), .C(n26149), .D(reg_A[94]), .Y(
        n29597) );
  AOI22X1 U24081 ( .A(n26148), .B(reg_A[92]), .C(reg_A[91]), .D(n25984), .Y(
        n29596) );
  NOR2X1 U24082 ( .A(n25873), .B(n25972), .Y(n25902) );
  AND2X1 U24083 ( .A(n29598), .B(n29599), .Y(n28660) );
  AOI22X1 U24084 ( .A(n26276), .B(reg_A[77]), .C(n26148), .D(reg_A[76]), .Y(
        n29599) );
  AOI22X1 U24085 ( .A(reg_A[75]), .B(n25984), .C(n26149), .D(reg_A[78]), .Y(
        n29598) );
  OAI21X1 U24086 ( .A(n26169), .B(n29137), .C(n29600), .Y(n29586) );
  AOI22X1 U24087 ( .A(n29601), .B(n26276), .C(n28930), .D(n29114), .Y(n29600)
         );
  OAI21X1 U24088 ( .A(n26547), .B(n26168), .C(n29602), .Y(n29114) );
  AOI22X1 U24089 ( .A(n26276), .B(reg_A[73]), .C(n26149), .D(reg_A[74]), .Y(
        n29602) );
  INVX1 U24090 ( .A(n29413), .Y(n29601) );
  NAND2X1 U24091 ( .A(reg_A[70]), .B(n26057), .Y(n29137) );
  AOI22X1 U24092 ( .A(n29603), .B(reg_B[76]), .C(n29604), .D(n29605), .Y(
        n29582) );
  NOR2X1 U24093 ( .A(n26101), .B(n29096), .Y(n29604) );
  NOR2X1 U24094 ( .A(n28639), .B(n25415), .Y(n29603) );
  MUX2X1 U24095 ( .B(n29118), .A(n29606), .S(reg_B[77]), .Y(n28639) );
  NOR2X1 U24096 ( .A(n25864), .B(n28088), .Y(n29606) );
  NAND2X1 U24097 ( .A(n29607), .B(n29608), .Y(n29118) );
  AOI22X1 U24098 ( .A(n28602), .B(reg_A[77]), .C(n28191), .D(reg_A[76]), .Y(
        n29608) );
  AOI22X1 U24099 ( .A(n28245), .B(reg_A[78]), .C(n28446), .D(reg_A[75]), .Y(
        n29607) );
  NAND2X1 U24100 ( .A(reg_B[95]), .B(n25699), .Y(n27020) );
  OAI21X1 U24101 ( .A(n29609), .B(n28130), .C(n29610), .Y(n29570) );
  AOI22X1 U24102 ( .A(n29457), .B(n29399), .C(n29057), .D(n29611), .Y(n29610)
         );
  NOR2X1 U24103 ( .A(n29221), .B(n26151), .Y(n29057) );
  INVX1 U24104 ( .A(n29509), .Y(n29399) );
  NAND2X1 U24105 ( .A(reg_B[79]), .B(n26267), .Y(n28130) );
  NOR2X1 U24106 ( .A(n29612), .B(n29613), .Y(n29539) );
  OAI21X1 U24107 ( .A(n29614), .B(n26990), .C(n29615), .Y(n29613) );
  OAI21X1 U24108 ( .A(n29616), .B(n29617), .C(n25372), .Y(n29615) );
  OAI21X1 U24109 ( .A(n29618), .B(n25884), .C(n29619), .Y(n29617) );
  AOI22X1 U24110 ( .A(n29457), .B(n29620), .C(n27787), .D(n29449), .Y(n29619)
         );
  INVX1 U24111 ( .A(n29551), .Y(n29449) );
  AOI22X1 U24112 ( .A(reg_A[65]), .B(n29412), .C(n25950), .D(n29621), .Y(
        n29551) );
  INVX1 U24113 ( .A(n26896), .Y(n27787) );
  NAND2X1 U24114 ( .A(n25044), .B(n25976), .Y(n26896) );
  INVX1 U24115 ( .A(n29020), .Y(n29620) );
  NAND2X1 U24116 ( .A(n25029), .B(n29221), .Y(n29020) );
  AND2X1 U24117 ( .A(n29622), .B(n29026), .Y(n29457) );
  MUX2X1 U24118 ( .B(n25851), .A(n25855), .S(reg_B[70]), .Y(n29622) );
  OAI21X1 U24119 ( .A(n29623), .B(n25853), .C(n29624), .Y(n29616) );
  AOI21X1 U24120 ( .A(n29625), .B(n25604), .C(n29626), .Y(n29624) );
  INVX1 U24121 ( .A(n29459), .Y(n29626) );
  NOR2X1 U24122 ( .A(reg_B[79]), .B(n29505), .Y(n29625) );
  INVX1 U24123 ( .A(n29460), .Y(n29505) );
  OAI21X1 U24124 ( .A(n25855), .B(n28879), .C(n29627), .Y(n29460) );
  NAND3X1 U24125 ( .A(reg_A[67]), .B(n28377), .C(n28297), .Y(n29627) );
  AOI21X1 U24126 ( .A(n26149), .B(n25097), .C(n29628), .Y(n29623) );
  OAI22X1 U24127 ( .A(n25415), .B(n28208), .C(n26999), .D(n29629), .Y(n29628)
         );
  NOR2X1 U24128 ( .A(n29630), .B(n29631), .Y(n29614) );
  NAND3X1 U24129 ( .A(n29632), .B(n29633), .C(n29634), .Y(n29631) );
  NOR2X1 U24130 ( .A(n29635), .B(n29636), .Y(n29634) );
  OAI21X1 U24131 ( .A(n25034), .B(n26103), .C(n29637), .Y(n29636) );
  AOI22X1 U24132 ( .A(reg_A[72]), .B(n25123), .C(reg_A[76]), .D(n25629), .Y(
        n29637) );
  NAND2X1 U24133 ( .A(n29638), .B(n29639), .Y(n29635) );
  AOI22X1 U24134 ( .A(reg_A[69]), .B(n25252), .C(reg_A[73]), .D(n25253), .Y(
        n29639) );
  AOI22X1 U24135 ( .A(reg_A[74]), .B(n25628), .C(reg_A[71]), .D(n25069), .Y(
        n29638) );
  NOR2X1 U24136 ( .A(n29640), .B(n29641), .Y(n29633) );
  OAI22X1 U24137 ( .A(n25065), .B(n25874), .C(n25035), .D(n26094), .Y(n29641)
         );
  OAI22X1 U24138 ( .A(n25036), .B(n26286), .C(n25473), .D(n25865), .Y(n29640)
         );
  AOI21X1 U24139 ( .A(reg_A[67]), .B(n25125), .C(n29642), .Y(n29632) );
  OAI22X1 U24140 ( .A(n25039), .B(n25584), .C(n25231), .D(n25864), .Y(n29642)
         );
  NAND3X1 U24141 ( .A(n29643), .B(n29644), .C(n29645), .Y(n29630) );
  NOR2X1 U24142 ( .A(n29646), .B(n29647), .Y(n29645) );
  OAI21X1 U24143 ( .A(n25041), .B(n26256), .C(n29648), .Y(n29647) );
  AOI22X1 U24144 ( .A(reg_A[95]), .B(n25324), .C(reg_A[68]), .D(n25135), .Y(
        n29648) );
  NAND2X1 U24145 ( .A(n29649), .B(n29650), .Y(n29646) );
  AOI22X1 U24146 ( .A(reg_A[92]), .B(n25857), .C(reg_A[91]), .D(n25647), .Y(
        n29650) );
  AOI22X1 U24147 ( .A(reg_A[94]), .B(n25648), .C(reg_A[93]), .D(n26432), .Y(
        n29649) );
  NOR2X1 U24148 ( .A(n29651), .B(n29652), .Y(n29644) );
  OAI22X1 U24149 ( .A(n25331), .B(n26215), .C(n25243), .D(n26039), .Y(n29652)
         );
  INVX1 U24150 ( .A(reg_A[86]), .Y(n26039) );
  INVX1 U24151 ( .A(reg_A[85]), .Y(n26215) );
  OAI22X1 U24152 ( .A(n25334), .B(n25875), .C(n25336), .D(n26230), .Y(n29651)
         );
  NOR2X1 U24153 ( .A(n29653), .B(n29654), .Y(n29643) );
  OAI22X1 U24154 ( .A(n26719), .B(n26195), .C(n25238), .D(n25965), .Y(n29654)
         );
  OAI22X1 U24155 ( .A(n25491), .B(n26068), .C(n25492), .D(n25929), .Y(n29653)
         );
  OAI22X1 U24156 ( .A(n25583), .B(n29655), .C(n29656), .D(n25853), .Y(n29612)
         );
  OR2X1 U24157 ( .A(n29657), .B(n29658), .Y(result[66]) );
  NAND3X1 U24158 ( .A(n29659), .B(n29660), .C(n29661), .Y(n29658) );
  NOR2X1 U24159 ( .A(n29662), .B(n29663), .Y(n29661) );
  OAI21X1 U24160 ( .A(n29609), .B(n29409), .C(n29664), .Y(n29663) );
  OAI21X1 U24161 ( .A(n29665), .B(n29666), .C(n25203), .Y(n29664) );
  NAND3X1 U24162 ( .A(n29667), .B(n29668), .C(n29669), .Y(n29666) );
  AOI21X1 U24163 ( .A(reg_A[66]), .B(n25434), .C(n29670), .Y(n29669) );
  OAI22X1 U24164 ( .A(n25437), .B(n26107), .C(n25438), .D(n26256), .Y(n29670)
         );
  AOI22X1 U24165 ( .A(reg_A[76]), .B(n25439), .C(reg_A[72]), .D(n25440), .Y(
        n29668) );
  AOI22X1 U24166 ( .A(reg_A[67]), .B(n25441), .C(reg_A[69]), .D(n25442), .Y(
        n29667) );
  NAND3X1 U24167 ( .A(n29671), .B(n29672), .C(n29673), .Y(n29665) );
  NOR2X1 U24168 ( .A(n29674), .B(n29675), .Y(n29673) );
  OAI22X1 U24169 ( .A(n25449), .B(n26101), .C(n25451), .D(n25865), .Y(n29675)
         );
  OAI21X1 U24170 ( .A(n25453), .B(n25864), .C(n29676), .Y(n29674) );
  OAI21X1 U24171 ( .A(n29677), .B(n29678), .C(n25044), .Y(n29676) );
  NAND3X1 U24172 ( .A(n29679), .B(n29680), .C(n29681), .Y(n29678) );
  NOR2X1 U24173 ( .A(n29682), .B(n29683), .Y(n29681) );
  OAI21X1 U24174 ( .A(n25043), .B(n25884), .C(n29684), .Y(n29683) );
  AOI22X1 U24175 ( .A(reg_A[67]), .B(n25135), .C(reg_A[68]), .D(n25252), .Y(
        n29684) );
  NAND2X1 U24176 ( .A(n29685), .B(n29686), .Y(n29682) );
  AOI22X1 U24177 ( .A(reg_A[69]), .B(n25136), .C(reg_A[72]), .D(n25253), .Y(
        n29686) );
  AOI22X1 U24178 ( .A(reg_A[70]), .B(n25071), .C(reg_A[71]), .D(n25123), .Y(
        n29685) );
  NOR2X1 U24179 ( .A(n29687), .B(n29688), .Y(n29680) );
  OAI22X1 U24180 ( .A(n25034), .B(n26438), .C(n25129), .D(n26439), .Y(n29688)
         );
  OAI22X1 U24181 ( .A(n25036), .B(n25863), .C(n25223), .D(n26103), .Y(n29687)
         );
  INVX1 U24182 ( .A(reg_A[75]), .Y(n26103) );
  NOR2X1 U24183 ( .A(n29689), .B(n29690), .Y(n29679) );
  OAI22X1 U24184 ( .A(n25064), .B(n25865), .C(n25473), .D(n26286), .Y(n29690)
         );
  OAI22X1 U24185 ( .A(n25039), .B(n25864), .C(n25035), .D(n25584), .Y(n29689)
         );
  NAND3X1 U24186 ( .A(n29691), .B(n29692), .C(n29693), .Y(n29677) );
  NOR2X1 U24187 ( .A(n29694), .B(n29695), .Y(n29693) );
  OAI21X1 U24188 ( .A(n25065), .B(n26094), .C(n29696), .Y(n29695) );
  AOI22X1 U24189 ( .A(reg_A[83]), .B(n25246), .C(reg_A[82]), .D(n25247), .Y(
        n29696) );
  NAND2X1 U24190 ( .A(n29697), .B(n29698), .Y(n29694) );
  AOI22X1 U24191 ( .A(reg_A[85]), .B(n25487), .C(reg_A[84]), .D(n25241), .Y(
        n29698) );
  AOI22X1 U24192 ( .A(reg_A[86]), .B(n25339), .C(reg_A[87]), .D(n25257), .Y(
        n29697) );
  NOR2X1 U24193 ( .A(n29699), .B(n29700), .Y(n29692) );
  OAI22X1 U24194 ( .A(n25491), .B(n25929), .C(n25492), .D(n26195), .Y(n29700)
         );
  OAI22X1 U24195 ( .A(n25320), .B(n26068), .C(n25322), .D(n25973), .Y(n29699)
         );
  NOR2X1 U24196 ( .A(n29701), .B(n29702), .Y(n29691) );
  OAI22X1 U24197 ( .A(n25316), .B(n25882), .C(n25318), .D(n25881), .Y(n29702)
         );
  INVX1 U24198 ( .A(reg_A[92]), .Y(n25882) );
  OAI22X1 U24199 ( .A(n25498), .B(n25873), .C(n25499), .D(n25883), .Y(n29701)
         );
  AOI22X1 U24200 ( .A(reg_A[75]), .B(n25500), .C(reg_A[74]), .D(n25501), .Y(
        n29672) );
  AOI22X1 U24201 ( .A(reg_A[73]), .B(n25502), .C(reg_A[77]), .D(n25503), .Y(
        n29671) );
  NAND2X1 U24202 ( .A(n26267), .B(n28248), .Y(n29409) );
  INVX1 U24203 ( .A(n29703), .Y(n29609) );
  OAI21X1 U24204 ( .A(n25853), .B(n28879), .C(n29704), .Y(n29703) );
  NAND3X1 U24205 ( .A(reg_A[66]), .B(n28377), .C(n28297), .Y(n29704) );
  NAND2X1 U24206 ( .A(n28297), .B(reg_B[78]), .Y(n28879) );
  AOI22X1 U24207 ( .A(reg_A[68]), .B(n25506), .C(reg_A[69]), .D(n25507), .Y(
        n29660) );
  AOI22X1 U24208 ( .A(reg_A[70]), .B(n25508), .C(reg_A[71]), .D(n25509), .Y(
        n29659) );
  NAND3X1 U24209 ( .A(n29705), .B(n29706), .C(n29707), .Y(n29657) );
  NOR2X1 U24210 ( .A(n29708), .B(n29709), .Y(n29707) );
  OAI21X1 U24211 ( .A(n29710), .B(n25517), .C(n29711), .Y(n29709) );
  OAI21X1 U24212 ( .A(n29712), .B(n29713), .C(reg_A[65]), .Y(n29711) );
  OAI21X1 U24213 ( .A(n29618), .B(n25517), .C(n25566), .Y(n29713) );
  INVX1 U24214 ( .A(n29578), .Y(n29618) );
  OAI21X1 U24215 ( .A(n26168), .B(n29714), .C(n29715), .Y(n29578) );
  NAND2X1 U24216 ( .A(n26057), .B(n25044), .Y(n29714) );
  INVX1 U24217 ( .A(n29716), .Y(n29712) );
  OAI21X1 U24218 ( .A(n29717), .B(n29509), .C(n29718), .Y(n29708) );
  OAI21X1 U24219 ( .A(n29719), .B(n29720), .C(reg_A[64]), .Y(n29718) );
  NAND2X1 U24220 ( .A(n25528), .B(n29217), .Y(n29720) );
  NAND2X1 U24221 ( .A(reg_B[70]), .B(n26504), .Y(n29217) );
  NAND2X1 U24222 ( .A(n28407), .B(n28728), .Y(n29719) );
  NAND2X1 U24223 ( .A(reg_B[94]), .B(n25932), .Y(n28728) );
  NAND2X1 U24224 ( .A(reg_B[78]), .B(n25188), .Y(n28407) );
  NAND2X1 U24225 ( .A(n26186), .B(n29221), .Y(n29509) );
  INVX1 U24226 ( .A(n29611), .Y(n29717) );
  MUX2X1 U24227 ( .B(n29416), .A(n29721), .S(reg_B[70]), .Y(n29611) );
  NAND2X1 U24228 ( .A(n29026), .B(reg_A[64]), .Y(n29721) );
  NAND2X1 U24229 ( .A(reg_A[66]), .B(n29026), .Y(n29416) );
  OAI21X1 U24230 ( .A(n29722), .B(n29723), .C(n25382), .Y(n29706) );
  OR2X1 U24231 ( .A(n29724), .B(n29725), .Y(n29723) );
  OAI21X1 U24232 ( .A(n29726), .B(n25856), .C(n29710), .Y(n29725) );
  AOI22X1 U24233 ( .A(n29462), .B(reg_A[66]), .C(n25963), .D(n29523), .Y(
        n29710) );
  INVX1 U24234 ( .A(n29136), .Y(n25963) );
  OAI21X1 U24235 ( .A(n29715), .B(n25851), .C(n29727), .Y(n29724) );
  AOI22X1 U24236 ( .A(n29134), .B(n29147), .C(reg_A[68]), .D(n29461), .Y(
        n29727) );
  NAND2X1 U24237 ( .A(n29728), .B(n29729), .Y(n29147) );
  AOI22X1 U24238 ( .A(n28602), .B(reg_A[72]), .C(n28191), .D(reg_A[71]), .Y(
        n29729) );
  AOI22X1 U24239 ( .A(n28245), .B(reg_A[73]), .C(n28446), .D(reg_A[70]), .Y(
        n29728) );
  NAND2X1 U24240 ( .A(n29730), .B(n29731), .Y(n29722) );
  AOI21X1 U24241 ( .A(n28103), .B(n28801), .C(n29732), .Y(n29731) );
  OAI21X1 U24242 ( .A(n29136), .B(n28730), .C(n29733), .Y(n29732) );
  OAI21X1 U24243 ( .A(n29734), .B(n29735), .C(n25044), .Y(n29733) );
  OAI21X1 U24244 ( .A(n28696), .B(n25964), .C(n29736), .Y(n29735) );
  AOI22X1 U24245 ( .A(reg_B[91]), .B(n27706), .C(n28826), .D(n28796), .Y(
        n29736) );
  NAND2X1 U24246 ( .A(n29737), .B(n29738), .Y(n28796) );
  AOI22X1 U24247 ( .A(n26276), .B(reg_A[80]), .C(n26149), .D(reg_A[81]), .Y(
        n29738) );
  AOI22X1 U24248 ( .A(n26148), .B(reg_A[79]), .C(reg_A[78]), .D(n25984), .Y(
        n29737) );
  NAND2X1 U24249 ( .A(n29739), .B(n29740), .Y(n27706) );
  AOI22X1 U24250 ( .A(n26274), .B(n28800), .C(n25989), .D(n26114), .Y(n29740)
         );
  OAI21X1 U24251 ( .A(n25873), .B(n26168), .C(n26170), .Y(n26114) );
  NAND2X1 U24252 ( .A(reg_A[94]), .B(n25984), .Y(n26170) );
  INVX1 U24253 ( .A(reg_A[95]), .Y(n25873) );
  NAND2X1 U24254 ( .A(n29741), .B(n29742), .Y(n28800) );
  AOI22X1 U24255 ( .A(reg_A[88]), .B(n26276), .C(n26149), .D(reg_A[89]), .Y(
        n29742) );
  AOI22X1 U24256 ( .A(n26148), .B(reg_A[87]), .C(reg_A[86]), .D(n25984), .Y(
        n29741) );
  AOI22X1 U24257 ( .A(n26275), .B(n28795), .C(n25988), .D(n28799), .Y(n29739)
         );
  NAND2X1 U24258 ( .A(n29743), .B(n29744), .Y(n28799) );
  AOI22X1 U24259 ( .A(reg_A[92]), .B(n26276), .C(n26149), .D(reg_A[93]), .Y(
        n29744) );
  AOI22X1 U24260 ( .A(n26148), .B(reg_A[91]), .C(reg_A[90]), .D(n25984), .Y(
        n29743) );
  NAND2X1 U24261 ( .A(n29745), .B(n29746), .Y(n28795) );
  AOI22X1 U24262 ( .A(reg_A[84]), .B(n26276), .C(n26149), .D(reg_A[85]), .Y(
        n29746) );
  AOI22X1 U24263 ( .A(n26148), .B(reg_A[83]), .C(reg_A[82]), .D(n25984), .Y(
        n29745) );
  AND2X1 U24264 ( .A(n29747), .B(n29748), .Y(n28696) );
  AOI22X1 U24265 ( .A(reg_A[76]), .B(n26276), .C(n26148), .D(reg_A[75]), .Y(
        n29748) );
  AOI22X1 U24266 ( .A(reg_A[74]), .B(n25984), .C(n26149), .D(reg_A[77]), .Y(
        n29747) );
  NAND2X1 U24267 ( .A(n29749), .B(n29750), .Y(n29734) );
  AOI22X1 U24268 ( .A(n26276), .B(n29197), .C(n29144), .D(n28930), .Y(n29750)
         );
  OAI22X1 U24269 ( .A(n26439), .B(n26169), .C(n25914), .D(n26547), .Y(n29144)
         );
  INVX1 U24270 ( .A(n29751), .Y(n29749) );
  OAI21X1 U24271 ( .A(n26169), .B(n29413), .C(n29752), .Y(n29751) );
  OAI21X1 U24272 ( .A(n29621), .B(n28609), .C(n26148), .Y(n29752) );
  NOR2X1 U24273 ( .A(n26997), .B(n26101), .Y(n28609) );
  NAND2X1 U24274 ( .A(n26057), .B(reg_A[69]), .Y(n29413) );
  NAND2X1 U24275 ( .A(n28930), .B(reg_A[70]), .Y(n28730) );
  NAND3X1 U24276 ( .A(n28259), .B(n28783), .C(n29753), .Y(n28801) );
  INVX1 U24277 ( .A(n29754), .Y(n29753) );
  OAI21X1 U24278 ( .A(n28208), .B(n26286), .C(n28475), .Y(n29754) );
  NAND2X1 U24279 ( .A(n28191), .B(reg_A[75]), .Y(n28475) );
  NAND2X1 U24280 ( .A(n28446), .B(reg_A[74]), .Y(n28783) );
  NAND2X1 U24281 ( .A(n28602), .B(reg_A[76]), .Y(n28259) );
  INVX1 U24282 ( .A(n29755), .Y(n29730) );
  OAI22X1 U24283 ( .A(n29756), .B(n29150), .C(n29757), .D(n28216), .Y(n29755)
         );
  AOI21X1 U24284 ( .A(reg_A[79]), .B(n28191), .C(n28258), .Y(n28216) );
  NOR2X1 U24285 ( .A(n28088), .B(n25865), .Y(n28258) );
  AOI22X1 U24286 ( .A(reg_A[70]), .B(n29201), .C(reg_A[71]), .D(n29758), .Y(
        n29150) );
  INVX1 U24287 ( .A(n29759), .Y(n29705) );
  OAI22X1 U24288 ( .A(n25518), .B(n25884), .C(n26950), .D(n29572), .Y(n29759)
         );
  AOI22X1 U24289 ( .A(n25950), .B(n29523), .C(reg_A[64]), .D(n29412), .Y(
        n29572) );
  NOR2X1 U24290 ( .A(n25966), .B(n25950), .Y(n29412) );
  NAND2X1 U24291 ( .A(n25699), .B(n25976), .Y(n26950) );
  NAND3X1 U24292 ( .A(n29760), .B(n29761), .C(n29762), .Y(result[65]) );
  NOR2X1 U24293 ( .A(n29763), .B(n29764), .Y(n29762) );
  OAI22X1 U24294 ( .A(n29765), .B(n26107), .C(n29766), .D(n25851), .Y(n29764)
         );
  NAND3X1 U24295 ( .A(n29767), .B(n29768), .C(n29769), .Y(n29763) );
  OAI21X1 U24296 ( .A(n29770), .B(n29771), .C(reg_A[65]), .Y(n29769) );
  OAI21X1 U24297 ( .A(n29772), .B(n25517), .C(n25706), .Y(n29771) );
  INVX1 U24298 ( .A(n29773), .Y(n25706) );
  INVX1 U24299 ( .A(n29585), .Y(n29772) );
  OAI21X1 U24300 ( .A(n25966), .B(n29136), .C(n29774), .Y(n29585) );
  NAND2X1 U24301 ( .A(n25984), .B(n25044), .Y(n29136) );
  OAI21X1 U24302 ( .A(n29775), .B(n29776), .C(reg_A[64]), .Y(n29768) );
  NAND2X1 U24303 ( .A(n29716), .B(n25693), .Y(n29776) );
  AOI22X1 U24304 ( .A(n29777), .B(n25170), .C(n26057), .D(n28547), .Y(n29716)
         );
  NOR2X1 U24305 ( .A(n26168), .B(n26610), .Y(n28547) );
  OAI21X1 U24306 ( .A(n25984), .B(n27438), .C(n29778), .Y(n29775) );
  AOI22X1 U24307 ( .A(n25188), .B(n28088), .C(n26504), .D(n29096), .Y(n29778)
         );
  NAND2X1 U24308 ( .A(reg_A[71]), .B(n29779), .Y(n29767) );
  AOI21X1 U24309 ( .A(n25203), .B(n29780), .C(n29781), .Y(n29761) );
  OAI22X1 U24310 ( .A(n25652), .B(n26256), .C(n29782), .D(n25856), .Y(n29781)
         );
  NAND3X1 U24311 ( .A(n29783), .B(n29784), .C(n29785), .Y(n29780) );
  NOR2X1 U24312 ( .A(n29786), .B(n29787), .Y(n29785) );
  OAI22X1 U24313 ( .A(n25598), .B(n25851), .C(n25599), .D(n26107), .Y(n29787)
         );
  OAI21X1 U24314 ( .A(n25600), .B(n26256), .C(n29788), .Y(n29786) );
  OAI21X1 U24315 ( .A(n29789), .B(n29790), .C(n25604), .Y(n29788) );
  NAND2X1 U24316 ( .A(n29791), .B(n29792), .Y(n29790) );
  AOI22X1 U24317 ( .A(reg_A[75]), .B(n25607), .C(reg_A[79]), .D(n25608), .Y(
        n29792) );
  AOI22X1 U24318 ( .A(reg_A[77]), .B(n25609), .C(reg_A[78]), .D(n25610), .Y(
        n29791) );
  NAND2X1 U24319 ( .A(n29793), .B(n29794), .Y(n29789) );
  AOI22X1 U24320 ( .A(reg_A[72]), .B(n25613), .C(reg_A[74]), .D(n25614), .Y(
        n29794) );
  AOI22X1 U24321 ( .A(reg_A[73]), .B(n25615), .C(reg_A[76]), .D(n25616), .Y(
        n29793) );
  AOI21X1 U24322 ( .A(reg_A[66]), .B(n25617), .C(n29795), .Y(n29784) );
  OAI21X1 U24323 ( .A(n25619), .B(n25855), .C(n29796), .Y(n29795) );
  OAI21X1 U24324 ( .A(n29797), .B(n29798), .C(n25044), .Y(n29796) );
  NAND2X1 U24325 ( .A(n29799), .B(n29800), .Y(n29798) );
  NOR2X1 U24326 ( .A(n29801), .B(n29802), .Y(n29800) );
  OAI21X1 U24327 ( .A(n25034), .B(n26439), .C(n29803), .Y(n29802) );
  AOI22X1 U24328 ( .A(reg_A[72]), .B(n25628), .C(reg_A[74]), .D(n25629), .Y(
        n29803) );
  OAI21X1 U24329 ( .A(n25498), .B(n25883), .C(n29804), .Y(n29801) );
  AOI22X1 U24330 ( .A(reg_A[95]), .B(n25631), .C(reg_A[93]), .D(n25324), .Y(
        n29804) );
  INVX1 U24331 ( .A(reg_A[94]), .Y(n25883) );
  NOR2X1 U24332 ( .A(n29805), .B(n29806), .Y(n29799) );
  OAI21X1 U24333 ( .A(n25039), .B(n25865), .C(n29807), .Y(n29806) );
  AOI22X1 U24334 ( .A(reg_A[80]), .B(n25235), .C(reg_A[77]), .D(n25635), .Y(
        n29807) );
  INVX1 U24335 ( .A(reg_A[78]), .Y(n25865) );
  OAI21X1 U24336 ( .A(n25035), .B(n25864), .C(n29808), .Y(n29805) );
  AOI22X1 U24337 ( .A(reg_A[76]), .B(n25222), .C(reg_A[75]), .D(n25637), .Y(
        n29808) );
  NAND2X1 U24338 ( .A(n29809), .B(n29810), .Y(n29797) );
  NOR2X1 U24339 ( .A(n29811), .B(n29812), .Y(n29810) );
  OAI21X1 U24340 ( .A(n25050), .B(n26195), .C(n29813), .Y(n29812) );
  AOI22X1 U24341 ( .A(reg_A[83]), .B(n25241), .C(reg_A[87]), .D(n25242), .Y(
        n29813) );
  OAI21X1 U24342 ( .A(n25038), .B(n26230), .C(n29814), .Y(n29811) );
  AOI22X1 U24343 ( .A(reg_A[82]), .B(n25246), .C(reg_A[81]), .D(n25247), .Y(
        n29814) );
  NOR2X1 U24344 ( .A(n29815), .B(n29816), .Y(n29809) );
  OAI21X1 U24345 ( .A(n25059), .B(n25973), .C(n29817), .Y(n29816) );
  AOI22X1 U24346 ( .A(reg_A[89]), .B(n25647), .C(reg_A[92]), .D(n25648), .Y(
        n29817) );
  OAI21X1 U24347 ( .A(n25054), .B(n26068), .C(n29818), .Y(n29815) );
  AOI22X1 U24348 ( .A(reg_A[85]), .B(n25339), .C(reg_A[86]), .D(n25257), .Y(
        n29818) );
  AOI22X1 U24349 ( .A(reg_A[69]), .B(n25650), .C(reg_A[71]), .D(n25651), .Y(
        n29783) );
  AOI21X1 U24350 ( .A(n25382), .B(n29819), .C(n29662), .Y(n29760) );
  OAI22X1 U24351 ( .A(n25517), .B(n29459), .C(n25583), .D(n29655), .Y(n29662)
         );
  OAI21X1 U24352 ( .A(n29820), .B(n29821), .C(reg_A[64]), .Y(n29459) );
  OAI21X1 U24353 ( .A(n26057), .B(n25403), .C(n29756), .Y(n29821) );
  NOR2X1 U24354 ( .A(n28297), .B(n25415), .Y(n29820) );
  NAND3X1 U24355 ( .A(n29822), .B(n29823), .C(n29824), .Y(n29819) );
  NOR2X1 U24356 ( .A(n29825), .B(n29826), .Y(n29824) );
  OAI21X1 U24357 ( .A(n29431), .B(n29107), .C(n29827), .Y(n29826) );
  OAI21X1 U24358 ( .A(n29828), .B(n29829), .C(n25044), .Y(n29827) );
  NAND2X1 U24359 ( .A(n29830), .B(n29831), .Y(n29829) );
  AOI22X1 U24360 ( .A(n28826), .B(n28340), .C(n26307), .D(n28825), .Y(n29831)
         );
  NAND2X1 U24361 ( .A(n29832), .B(n29833), .Y(n28825) );
  AOI22X1 U24362 ( .A(reg_A[75]), .B(n26276), .C(n26149), .D(reg_A[76]), .Y(
        n29833) );
  AOI22X1 U24363 ( .A(n26148), .B(reg_A[74]), .C(reg_A[73]), .D(n25984), .Y(
        n29832) );
  NAND2X1 U24364 ( .A(n29834), .B(n29835), .Y(n28340) );
  AOI22X1 U24365 ( .A(reg_A[79]), .B(n26276), .C(n26149), .D(reg_A[80]), .Y(
        n29835) );
  AOI22X1 U24366 ( .A(n26148), .B(reg_A[78]), .C(reg_A[77]), .D(n25984), .Y(
        n29834) );
  INVX1 U24367 ( .A(n28093), .Y(n28826) );
  AOI22X1 U24368 ( .A(reg_B[91]), .B(n27818), .C(n28930), .D(n29351), .Y(
        n29830) );
  NAND2X1 U24369 ( .A(n29836), .B(n29837), .Y(n29351) );
  AOI22X1 U24370 ( .A(reg_A[71]), .B(n26276), .C(n26149), .D(reg_A[72]), .Y(
        n29837) );
  AOI22X1 U24371 ( .A(n26148), .B(reg_A[70]), .C(reg_A[69]), .D(n25984), .Y(
        n29836) );
  INVX1 U24372 ( .A(n26997), .Y(n28930) );
  NAND2X1 U24373 ( .A(n29838), .B(n29839), .Y(n27818) );
  AOI22X1 U24374 ( .A(n26274), .B(n28461), .C(n25989), .D(n28460), .Y(n29839)
         );
  OAI21X1 U24375 ( .A(n25972), .B(n25881), .C(n29840), .Y(n28460) );
  AOI22X1 U24376 ( .A(reg_A[95]), .B(n26276), .C(n26148), .D(reg_A[94]), .Y(
        n29840) );
  NAND2X1 U24377 ( .A(n29841), .B(n29842), .Y(n28461) );
  AOI22X1 U24378 ( .A(reg_A[87]), .B(n26276), .C(n26149), .D(reg_A[88]), .Y(
        n29842) );
  AOI22X1 U24379 ( .A(n26148), .B(reg_A[86]), .C(reg_A[85]), .D(n25984), .Y(
        n29841) );
  AOI22X1 U24380 ( .A(n26275), .B(n28827), .C(n25988), .D(n28830), .Y(n29838)
         );
  NAND2X1 U24381 ( .A(n29843), .B(n29844), .Y(n28830) );
  AOI22X1 U24382 ( .A(reg_A[91]), .B(n26276), .C(n26149), .D(reg_A[92]), .Y(
        n29844) );
  AOI22X1 U24383 ( .A(n26148), .B(reg_A[90]), .C(reg_A[89]), .D(n25984), .Y(
        n29843) );
  NAND2X1 U24384 ( .A(n29845), .B(n29846), .Y(n28827) );
  AOI22X1 U24385 ( .A(reg_A[83]), .B(n26276), .C(n26149), .D(reg_A[84]), .Y(
        n29846) );
  AOI22X1 U24386 ( .A(n26148), .B(reg_A[82]), .C(reg_A[81]), .D(n25984), .Y(
        n29845) );
  NAND2X1 U24387 ( .A(n29847), .B(n29848), .Y(n29828) );
  AOI22X1 U24388 ( .A(n29849), .B(n26057), .C(n29621), .D(n26276), .Y(n29848)
         );
  NOR2X1 U24389 ( .A(n25851), .B(n25966), .Y(n29621) );
  NOR2X1 U24390 ( .A(n25972), .B(n25855), .Y(n29849) );
  AOI22X1 U24391 ( .A(n29197), .B(n26149), .C(n29523), .D(n26148), .Y(n29847)
         );
  INVX1 U24392 ( .A(n29068), .Y(n29197) );
  NAND2X1 U24393 ( .A(reg_A[68]), .B(n26057), .Y(n29068) );
  AND2X1 U24394 ( .A(n29850), .B(n29851), .Y(n29431) );
  AOI22X1 U24395 ( .A(n28602), .B(reg_A[71]), .C(n28191), .D(reg_A[70]), .Y(
        n29851) );
  AOI22X1 U24396 ( .A(n28245), .B(reg_A[72]), .C(n28446), .D(reg_A[69]), .Y(
        n29850) );
  OAI21X1 U24397 ( .A(n28819), .B(n29757), .C(n29852), .Y(n29825) );
  AOI22X1 U24398 ( .A(n28103), .B(n28817), .C(n29605), .D(n29433), .Y(n29852)
         );
  OAI21X1 U24399 ( .A(n25856), .B(n29096), .C(n29853), .Y(n29433) );
  AOI22X1 U24400 ( .A(n29758), .B(reg_A[70]), .C(n29854), .D(reg_A[71]), .Y(
        n29853) );
  INVX1 U24401 ( .A(n29855), .Y(n29854) );
  NAND2X1 U24402 ( .A(n29856), .B(n29857), .Y(n28817) );
  AOI22X1 U24403 ( .A(n28602), .B(reg_A[75]), .C(n28191), .D(reg_A[74]), .Y(
        n29857) );
  AOI22X1 U24404 ( .A(n28245), .B(reg_A[76]), .C(n28446), .D(reg_A[73]), .Y(
        n29856) );
  INVX1 U24405 ( .A(n28455), .Y(n28819) );
  OAI21X1 U24406 ( .A(n26286), .B(n28088), .C(n29858), .Y(n28455) );
  AOI22X1 U24407 ( .A(n28602), .B(reg_A[79]), .C(n28191), .D(reg_A[78]), .Y(
        n29858) );
  AOI22X1 U24408 ( .A(reg_A[67]), .B(n29461), .C(reg_A[66]), .D(n29777), .Y(
        n29823) );
  AOI22X1 U24409 ( .A(reg_A[68]), .B(n29581), .C(reg_A[65]), .D(n29462), .Y(
        n29822) );
  NAND3X1 U24410 ( .A(n29859), .B(n29860), .C(n29861), .Y(result[64]) );
  NOR2X1 U24411 ( .A(n29862), .B(n29863), .Y(n29861) );
  OAI22X1 U24412 ( .A(n25717), .B(n25884), .C(n25718), .D(n25851), .Y(n29863)
         );
  OAI21X1 U24413 ( .A(n25719), .B(n25855), .C(n29864), .Y(n29862) );
  AOI22X1 U24414 ( .A(reg_A[48]), .B(n25721), .C(reg_A[68]), .D(n25722), .Y(
        n29864) );
  AOI21X1 U24415 ( .A(n26928), .B(n29865), .C(n29866), .Y(n29860) );
  OAI21X1 U24416 ( .A(n29867), .B(n25853), .C(n29868), .Y(n29866) );
  OAI21X1 U24417 ( .A(n29869), .B(n29870), .C(n25730), .Y(n29868) );
  NAND3X1 U24418 ( .A(n29871), .B(n29872), .C(n29873), .Y(n29870) );
  NOR2X1 U24419 ( .A(n29874), .B(n29875), .Y(n29873) );
  OAI22X1 U24420 ( .A(n25736), .B(n25853), .C(n25737), .D(n26286), .Y(n29875)
         );
  OAI22X1 U24421 ( .A(n25738), .B(n25863), .C(n25739), .D(n25864), .Y(n29874)
         );
  AOI22X1 U24422 ( .A(reg_A[72]), .B(n25615), .C(reg_A[75]), .D(n25616), .Y(
        n29872) );
  AOI22X1 U24423 ( .A(reg_A[74]), .B(n25607), .C(reg_A[78]), .D(n25608), .Y(
        n29871) );
  NAND3X1 U24424 ( .A(n29876), .B(n29877), .C(n29878), .Y(n29869) );
  NOR2X1 U24425 ( .A(n29879), .B(n29880), .Y(n29878) );
  OAI22X1 U24426 ( .A(n25061), .B(n26256), .C(n25746), .D(n25884), .Y(n29880)
         );
  OAI22X1 U24427 ( .A(n25747), .B(n25851), .C(n25748), .D(n25855), .Y(n29879)
         );
  AOI22X1 U24428 ( .A(reg_A[71]), .B(n25613), .C(reg_A[68]), .D(n25749), .Y(
        n29877) );
  AOI22X1 U24429 ( .A(reg_A[69]), .B(n25750), .C(reg_A[73]), .D(n25614), .Y(
        n29876) );
  NOR2X1 U24430 ( .A(n29770), .B(n29881), .Y(n29867) );
  OAI21X1 U24431 ( .A(n29774), .B(n25697), .C(n29882), .Y(n29770) );
  NAND3X1 U24432 ( .A(n25984), .B(n25699), .C(n26057), .Y(n29882) );
  OAI21X1 U24433 ( .A(n26944), .B(n25856), .C(n29883), .Y(n29865) );
  AOI22X1 U24434 ( .A(reg_A[70]), .B(n26010), .C(reg_A[71]), .D(n26002), .Y(
        n29883) );
  AOI22X1 U24435 ( .A(n25310), .B(n29884), .C(n25382), .D(n29885), .Y(n29859)
         );
  NAND3X1 U24436 ( .A(n29886), .B(n29887), .C(n29888), .Y(n29885) );
  NOR2X1 U24437 ( .A(n29889), .B(n29890), .Y(n29888) );
  OAI21X1 U24438 ( .A(n29774), .B(n25853), .C(n29891), .Y(n29890) );
  OAI21X1 U24439 ( .A(n29892), .B(n29893), .C(n25044), .Y(n29891) );
  OAI21X1 U24440 ( .A(n29894), .B(n26997), .C(n29895), .Y(n29893) );
  AOI22X1 U24441 ( .A(n26307), .B(n29535), .C(reg_B[91]), .D(n27886), .Y(
        n29895) );
  NAND2X1 U24442 ( .A(n29896), .B(n29897), .Y(n27886) );
  AOI22X1 U24443 ( .A(n26274), .B(n28509), .C(n25989), .D(n26992), .Y(n29897)
         );
  NAND2X1 U24444 ( .A(n29898), .B(n29899), .Y(n26992) );
  AOI22X1 U24445 ( .A(reg_A[94]), .B(n26276), .C(n26149), .D(reg_A[95]), .Y(
        n29899) );
  AOI22X1 U24446 ( .A(n26148), .B(reg_A[93]), .C(reg_A[92]), .D(n25984), .Y(
        n29898) );
  NOR2X1 U24447 ( .A(n26197), .B(n26063), .Y(n25989) );
  NAND2X1 U24448 ( .A(n29900), .B(n29901), .Y(n28509) );
  AOI22X1 U24449 ( .A(reg_A[86]), .B(n26276), .C(n26149), .D(reg_A[87]), .Y(
        n29901) );
  AOI22X1 U24450 ( .A(n26148), .B(reg_A[85]), .C(reg_A[84]), .D(n25984), .Y(
        n29900) );
  AOI22X1 U24451 ( .A(n26275), .B(n29538), .C(n25988), .D(n26915), .Y(n29896)
         );
  NAND2X1 U24452 ( .A(n29902), .B(n29903), .Y(n26915) );
  AOI22X1 U24453 ( .A(reg_A[90]), .B(n26276), .C(n26149), .D(reg_A[91]), .Y(
        n29903) );
  AOI22X1 U24454 ( .A(n26148), .B(reg_A[89]), .C(reg_A[88]), .D(n25984), .Y(
        n29902) );
  NAND2X1 U24455 ( .A(n29904), .B(n29905), .Y(n29538) );
  AOI22X1 U24456 ( .A(reg_A[82]), .B(n26276), .C(n26149), .D(reg_A[83]), .Y(
        n29905) );
  AOI22X1 U24457 ( .A(n26148), .B(reg_A[81]), .C(reg_A[80]), .D(n25984), .Y(
        n29904) );
  NAND2X1 U24458 ( .A(n29906), .B(n29907), .Y(n29535) );
  AOI22X1 U24459 ( .A(reg_A[74]), .B(n26276), .C(n26149), .D(reg_A[75]), .Y(
        n29907) );
  AOI22X1 U24460 ( .A(n26148), .B(reg_A[73]), .C(reg_A[72]), .D(n25984), .Y(
        n29906) );
  INVX1 U24461 ( .A(n25964), .Y(n26307) );
  NAND2X1 U24462 ( .A(n25988), .B(n25895), .Y(n25964) );
  INVX1 U24463 ( .A(n26199), .Y(n25988) );
  NAND2X1 U24464 ( .A(reg_B[92]), .B(n26197), .Y(n26199) );
  NAND2X1 U24465 ( .A(n26274), .B(n25895), .Y(n26997) );
  INVX1 U24466 ( .A(n26069), .Y(n26274) );
  NAND2X1 U24467 ( .A(reg_B[93]), .B(n26063), .Y(n26069) );
  INVX1 U24468 ( .A(n29474), .Y(n29894) );
  NAND2X1 U24469 ( .A(n29908), .B(n29909), .Y(n29474) );
  AOI22X1 U24470 ( .A(reg_A[70]), .B(n26276), .C(n26149), .D(reg_A[71]), .Y(
        n29909) );
  AOI22X1 U24471 ( .A(n26148), .B(reg_A[69]), .C(reg_A[68]), .D(n25984), .Y(
        n29908) );
  OAI21X1 U24472 ( .A(n28561), .B(n28093), .C(n29910), .Y(n29892) );
  AOI22X1 U24473 ( .A(n26057), .B(n29911), .C(n29523), .D(n26276), .Y(n29910)
         );
  INVX1 U24474 ( .A(n29424), .Y(n29523) );
  NAND2X1 U24475 ( .A(reg_A[66]), .B(n26057), .Y(n29424) );
  OAI21X1 U24476 ( .A(n25972), .B(n25853), .C(n29912), .Y(n29911) );
  AOI22X1 U24477 ( .A(n26149), .B(reg_A[67]), .C(n26148), .D(reg_A[65]), .Y(
        n29912) );
  INVX1 U24478 ( .A(n25966), .Y(n26057) );
  NAND2X1 U24479 ( .A(n26275), .B(n25895), .Y(n25966) );
  NAND2X1 U24480 ( .A(reg_B[93]), .B(n25892), .Y(n28093) );
  INVX1 U24481 ( .A(n26131), .Y(n25892) );
  NAND2X1 U24482 ( .A(reg_B[92]), .B(n25895), .Y(n26131) );
  INVX1 U24483 ( .A(reg_B[91]), .Y(n25895) );
  INVX1 U24484 ( .A(n28931), .Y(n28561) );
  NAND2X1 U24485 ( .A(n29913), .B(n29914), .Y(n28931) );
  AOI22X1 U24486 ( .A(reg_A[78]), .B(n26276), .C(n26149), .D(reg_A[79]), .Y(
        n29914) );
  NAND2X1 U24487 ( .A(reg_B[95]), .B(reg_B[94]), .Y(n26169) );
  NAND2X1 U24488 ( .A(reg_B[94]), .B(n25976), .Y(n25914) );
  AOI22X1 U24489 ( .A(n26148), .B(reg_A[77]), .C(reg_A[76]), .D(n25984), .Y(
        n29913) );
  NAND2X1 U24490 ( .A(reg_B[95]), .B(n25950), .Y(n26168) );
  INVX1 U24491 ( .A(n29462), .Y(n29774) );
  OAI21X1 U24492 ( .A(n28088), .B(n29102), .C(n29015), .Y(n29462) );
  NAND2X1 U24493 ( .A(n29434), .B(n29201), .Y(n29015) );
  INVX1 U24494 ( .A(n29151), .Y(n29434) );
  OAI22X1 U24495 ( .A(n29726), .B(n25851), .C(n29715), .D(n25855), .Y(n29889)
         );
  INVX1 U24496 ( .A(n29777), .Y(n29715) );
  OAI22X1 U24497 ( .A(n28193), .B(n29102), .C(n29095), .D(n29151), .Y(n29777)
         );
  INVX1 U24498 ( .A(n29581), .Y(n29726) );
  OAI22X1 U24499 ( .A(n28208), .B(n29102), .C(n29151), .D(n29629), .Y(n29581)
         );
  AOI21X1 U24500 ( .A(n29605), .B(n29531), .C(n29915), .Y(n29887) );
  INVX1 U24501 ( .A(n29916), .Y(n29915) );
  AOI22X1 U24502 ( .A(n29461), .B(reg_A[66]), .C(n28924), .D(n28103), .Y(
        n29916) );
  INVX1 U24503 ( .A(n29149), .Y(n28103) );
  NAND2X1 U24504 ( .A(n28073), .B(n25604), .Y(n29149) );
  INVX1 U24505 ( .A(n28393), .Y(n28073) );
  NAND2X1 U24506 ( .A(reg_B[76]), .B(n28192), .Y(n28393) );
  NAND2X1 U24507 ( .A(n29917), .B(n29918), .Y(n28924) );
  AOI22X1 U24508 ( .A(n28602), .B(reg_A[74]), .C(n28191), .D(reg_A[73]), .Y(
        n29918) );
  AOI22X1 U24509 ( .A(n28245), .B(reg_A[75]), .C(n28446), .D(reg_A[72]), .Y(
        n29917) );
  OAI22X1 U24510 ( .A(n28144), .B(n29102), .C(n29151), .D(n29855), .Y(n29461)
         );
  NAND2X1 U24511 ( .A(n25029), .B(n29026), .Y(n29151) );
  INVX1 U24512 ( .A(reg_B[69]), .Y(n29026) );
  NAND2X1 U24513 ( .A(n28297), .B(n25604), .Y(n29102) );
  INVX1 U24514 ( .A(n28394), .Y(n28297) );
  NAND2X1 U24515 ( .A(n28295), .B(n28192), .Y(n28394) );
  INVX1 U24516 ( .A(reg_B[77]), .Y(n28192) );
  OR2X1 U24517 ( .A(n29919), .B(n29920), .Y(n29531) );
  OAI22X1 U24518 ( .A(n29629), .B(n26101), .C(n29095), .D(n25856), .Y(n29920)
         );
  INVX1 U24519 ( .A(n29758), .Y(n29095) );
  NOR2X1 U24520 ( .A(n29221), .B(reg_B[70]), .Y(n29758) );
  NAND2X1 U24521 ( .A(reg_B[70]), .B(reg_B[71]), .Y(n29629) );
  OAI22X1 U24522 ( .A(n29855), .B(n26256), .C(n29096), .D(n26107), .Y(n29919)
         );
  INVX1 U24523 ( .A(n29201), .Y(n29096) );
  NOR2X1 U24524 ( .A(reg_B[71]), .B(reg_B[70]), .Y(n29201) );
  NAND2X1 U24525 ( .A(reg_B[70]), .B(n29221), .Y(n29855) );
  INVX1 U24526 ( .A(reg_B[71]), .Y(n29221) );
  INVX1 U24527 ( .A(n29756), .Y(n29605) );
  NAND2X1 U24528 ( .A(reg_B[69]), .B(n25029), .Y(n29756) );
  AOI22X1 U24529 ( .A(n28104), .B(n28934), .C(n29134), .D(n29530), .Y(n29886)
         );
  NAND2X1 U24530 ( .A(n29921), .B(n29922), .Y(n29530) );
  AOI22X1 U24531 ( .A(n28602), .B(reg_A[70]), .C(n28191), .D(reg_A[69]), .Y(
        n29922) );
  AOI22X1 U24532 ( .A(n28245), .B(reg_A[71]), .C(n28446), .D(reg_A[68]), .Y(
        n29921) );
  INVX1 U24533 ( .A(n29107), .Y(n29134) );
  NAND2X1 U24534 ( .A(n28296), .B(n25604), .Y(n29107) );
  INVX1 U24535 ( .A(n28483), .Y(n28296) );
  NAND2X1 U24536 ( .A(reg_B[77]), .B(n28295), .Y(n28483) );
  INVX1 U24537 ( .A(reg_B[76]), .Y(n28295) );
  NAND2X1 U24538 ( .A(n29923), .B(n29924), .Y(n28934) );
  AOI22X1 U24539 ( .A(n28602), .B(reg_A[78]), .C(n28191), .D(reg_A[77]), .Y(
        n29924) );
  INVX1 U24540 ( .A(n28193), .Y(n28191) );
  NAND2X1 U24541 ( .A(reg_B[79]), .B(n28377), .Y(n28193) );
  INVX1 U24542 ( .A(n28144), .Y(n28602) );
  NAND2X1 U24543 ( .A(reg_B[78]), .B(n28248), .Y(n28144) );
  AOI22X1 U24544 ( .A(n28245), .B(reg_A[79]), .C(n28446), .D(reg_A[76]), .Y(
        n29923) );
  INVX1 U24545 ( .A(n28088), .Y(n28446) );
  NAND2X1 U24546 ( .A(n28377), .B(n28248), .Y(n28088) );
  INVX1 U24547 ( .A(reg_B[79]), .Y(n28248) );
  INVX1 U24548 ( .A(reg_B[78]), .Y(n28377) );
  INVX1 U24549 ( .A(n28208), .Y(n28245) );
  NAND2X1 U24550 ( .A(reg_B[79]), .B(reg_B[78]), .Y(n28208) );
  INVX1 U24551 ( .A(n29757), .Y(n28104) );
  NAND3X1 U24552 ( .A(reg_B[76]), .B(n25604), .C(reg_B[77]), .Y(n29757) );
  NAND2X1 U24553 ( .A(n29925), .B(n29926), .Y(n29884) );
  NOR2X1 U24554 ( .A(n29927), .B(n29928), .Y(n29926) );
  NAND3X1 U24555 ( .A(n29929), .B(n29930), .C(n29931), .Y(n29928) );
  NOR2X1 U24556 ( .A(n29932), .B(n29933), .Y(n29931) );
  OAI22X1 U24557 ( .A(n25316), .B(n26068), .C(n25318), .D(n25973), .Y(n29933)
         );
  INVX1 U24558 ( .A(reg_A[91]), .Y(n25973) );
  INVX1 U24559 ( .A(reg_A[90]), .Y(n26068) );
  OAI22X1 U24560 ( .A(n25320), .B(n26195), .C(n25322), .D(n25929), .Y(n29932)
         );
  AOI22X1 U24561 ( .A(reg_A[94]), .B(n25631), .C(reg_A[95]), .D(n25764), .Y(
        n29930) );
  AOI22X1 U24562 ( .A(reg_A[92]), .B(n25324), .C(reg_A[93]), .D(n25765), .Y(
        n29929) );
  NAND3X1 U24563 ( .A(n29934), .B(n29935), .C(n29936), .Y(n29927) );
  NOR2X1 U24564 ( .A(n29937), .B(n29938), .Y(n29936) );
  OAI22X1 U24565 ( .A(n25051), .B(n25874), .C(n25038), .D(n25875), .Y(n29938)
         );
  INVX1 U24566 ( .A(reg_A[83]), .Y(n25875) );
  OAI22X1 U24567 ( .A(n25334), .B(n25584), .C(n25336), .D(n26094), .Y(n29937)
         );
  AOI22X1 U24568 ( .A(reg_A[86]), .B(n25242), .C(reg_A[87]), .D(n25338), .Y(
        n29935) );
  AOI22X1 U24569 ( .A(reg_A[84]), .B(n25339), .C(reg_A[85]), .D(n25257), .Y(
        n29934) );
  NOR2X1 U24570 ( .A(n29939), .B(n29940), .Y(n29925) );
  NAND3X1 U24571 ( .A(n29941), .B(n29942), .C(n29943), .Y(n29940) );
  NOR2X1 U24572 ( .A(n29944), .B(n29945), .Y(n29943) );
  OAI22X1 U24573 ( .A(n25043), .B(n25853), .C(n25039), .D(n26286), .Y(n29945)
         );
  OAI22X1 U24574 ( .A(n25064), .B(n25863), .C(n25482), .D(n25864), .Y(n29944)
         );
  AOI22X1 U24575 ( .A(reg_A[72]), .B(n25124), .C(reg_A[75]), .D(n25222), .Y(
        n29942) );
  AOI22X1 U24576 ( .A(reg_A[74]), .B(n25637), .C(reg_A[78]), .D(n25234), .Y(
        n29941) );
  NAND3X1 U24577 ( .A(n29946), .B(n29947), .C(n29948), .Y(n29939) );
  NOR2X1 U24578 ( .A(n29949), .B(n29950), .Y(n29948) );
  OAI22X1 U24579 ( .A(n25033), .B(n26256), .C(n25040), .D(n25884), .Y(n29950)
         );
  OAI22X1 U24580 ( .A(n25041), .B(n25851), .C(n25042), .D(n25855), .Y(n29949)
         );
  AOI22X1 U24581 ( .A(reg_A[71]), .B(n25628), .C(reg_A[68]), .D(n25068), .Y(
        n29947) );
  AOI22X1 U24582 ( .A(reg_A[69]), .B(n25123), .C(reg_A[73]), .D(n25629), .Y(
        n29946) );
  NAND3X1 U24583 ( .A(n29951), .B(n29952), .C(n29953), .Y(result[63]) );
  NOR2X1 U24584 ( .A(n29954), .B(n29955), .Y(n29953) );
  OR2X1 U24585 ( .A(n29956), .B(n29957), .Y(n29955) );
  OAI21X1 U24586 ( .A(n29958), .B(n29959), .C(n29960), .Y(n29957) );
  AOI22X1 U24587 ( .A(n29961), .B(n28138), .C(n29962), .D(n29963), .Y(n29960)
         );
  OAI21X1 U24588 ( .A(n29964), .B(n29965), .C(n29966), .Y(n29956) );
  AOI22X1 U24589 ( .A(reg_A[62]), .B(n29967), .C(reg_A[63]), .D(n29968), .Y(
        n29966) );
  OAI21X1 U24590 ( .A(n29969), .B(n29970), .C(n29971), .Y(n29968) );
  INVX1 U24591 ( .A(n29972), .Y(n29971) );
  AOI21X1 U24592 ( .A(n26504), .B(n29973), .C(n29974), .Y(n29969) );
  OAI22X1 U24593 ( .A(n25794), .B(n29975), .C(n27438), .D(n29976), .Y(n29974)
         );
  OAI21X1 U24594 ( .A(n29977), .B(n29978), .C(n28194), .Y(n29967) );
  NAND2X1 U24595 ( .A(n29979), .B(n29980), .Y(n29954) );
  AOI21X1 U24596 ( .A(n29981), .B(n29982), .C(n29983), .Y(n29980) );
  OAI21X1 U24597 ( .A(n29984), .B(n29985), .C(n29986), .Y(n29983) );
  NAND3X1 U24598 ( .A(n29987), .B(n26186), .C(n29988), .Y(n29986) );
  MUX2X1 U24599 ( .B(n29989), .A(n29990), .S(reg_B[61]), .Y(n29988) );
  NAND2X1 U24600 ( .A(n29991), .B(n29992), .Y(n29985) );
  OAI21X1 U24601 ( .A(n29993), .B(n25697), .C(n25031), .Y(n29992) );
  OAI22X1 U24602 ( .A(n26996), .B(n29994), .C(n28105), .D(n29993), .Y(n29982)
         );
  AOI21X1 U24603 ( .A(n25188), .B(n29995), .C(n29996), .Y(n29979) );
  OAI21X1 U24604 ( .A(n29997), .B(n29998), .C(n29999), .Y(n29996) );
  OAI21X1 U24605 ( .A(n30000), .B(n30001), .C(n25918), .Y(n29999) );
  NAND3X1 U24606 ( .A(n30002), .B(n30003), .C(n30004), .Y(n30001) );
  NOR2X1 U24607 ( .A(n30005), .B(n30006), .Y(n30004) );
  OAI22X1 U24608 ( .A(n25736), .B(n30007), .C(n25737), .D(n30008), .Y(n30006)
         );
  OAI22X1 U24609 ( .A(n25738), .B(n30009), .C(n25739), .D(n29655), .Y(n30005)
         );
  AOI22X1 U24610 ( .A(reg_A[55]), .B(n25615), .C(reg_A[52]), .D(n25616), .Y(
        n30003) );
  AOI22X1 U24611 ( .A(reg_A[53]), .B(n25607), .C(reg_A[49]), .D(n25608), .Y(
        n30002) );
  NAND3X1 U24612 ( .A(n30010), .B(n30011), .C(n30012), .Y(n30000) );
  NOR2X1 U24613 ( .A(n30013), .B(n30014), .Y(n30012) );
  OAI22X1 U24614 ( .A(n25061), .B(n29990), .C(n25746), .D(n29989), .Y(n30014)
         );
  OAI22X1 U24615 ( .A(n25747), .B(n30015), .C(n25748), .D(n30016), .Y(n30013)
         );
  AOI22X1 U24616 ( .A(reg_A[56]), .B(n25613), .C(reg_A[59]), .D(n25749), .Y(
        n30011) );
  AOI22X1 U24617 ( .A(reg_A[58]), .B(n25750), .C(reg_A[54]), .D(n25614), .Y(
        n30010) );
  AOI21X1 U24618 ( .A(n30017), .B(n26601), .C(n30018), .Y(n29997) );
  INVX1 U24619 ( .A(n30019), .Y(n30018) );
  OAI21X1 U24620 ( .A(n30020), .B(n30021), .C(n30022), .Y(n29995) );
  NAND3X1 U24621 ( .A(n30023), .B(n30024), .C(reg_B[60]), .Y(n30022) );
  NOR2X1 U24622 ( .A(n30025), .B(n30026), .Y(n29952) );
  OAI21X1 U24623 ( .A(n30027), .B(n30028), .C(n30029), .Y(n30026) );
  AOI22X1 U24624 ( .A(n25932), .B(n30030), .C(reg_B[62]), .D(n30031), .Y(
        n30029) );
  OAI21X1 U24625 ( .A(n30032), .B(n30033), .C(n30034), .Y(n30030) );
  INVX1 U24626 ( .A(n30035), .Y(n30034) );
  OAI22X1 U24627 ( .A(n29970), .B(n30036), .C(n30037), .D(n30038), .Y(n30035)
         );
  AOI22X1 U24628 ( .A(reg_A[55]), .B(n30039), .C(n30040), .D(n30041), .Y(
        n30036) );
  INVX1 U24629 ( .A(n30042), .Y(n30027) );
  OAI21X1 U24630 ( .A(n30043), .B(n30044), .C(n30045), .Y(n30025) );
  AOI22X1 U24631 ( .A(n30046), .B(n25900), .C(n25840), .D(n30047), .Y(n30045)
         );
  NAND2X1 U24632 ( .A(n30048), .B(n30049), .Y(n30047) );
  NOR2X1 U24633 ( .A(n30050), .B(n30051), .Y(n30049) );
  NAND3X1 U24634 ( .A(n30052), .B(n30053), .C(n30054), .Y(n30051) );
  NOR2X1 U24635 ( .A(n30055), .B(n30056), .Y(n30054) );
  OAI22X1 U24636 ( .A(n25316), .B(n30057), .C(n25318), .D(n30058), .Y(n30056)
         );
  OAI22X1 U24637 ( .A(n25320), .B(n30059), .C(n25322), .D(n30060), .Y(n30055)
         );
  AOI22X1 U24638 ( .A(reg_A[33]), .B(n25631), .C(reg_A[32]), .D(n25764), .Y(
        n30053) );
  AOI22X1 U24639 ( .A(reg_A[35]), .B(n25324), .C(reg_A[34]), .D(n25765), .Y(
        n30052) );
  NAND3X1 U24640 ( .A(n30061), .B(n30062), .C(n30063), .Y(n30050) );
  NOR2X1 U24641 ( .A(n30064), .B(n30065), .Y(n30063) );
  OAI22X1 U24642 ( .A(n25051), .B(n30066), .C(n25038), .D(n30067), .Y(n30065)
         );
  OAI22X1 U24643 ( .A(n25334), .B(n30068), .C(n25336), .D(n30069), .Y(n30064)
         );
  AOI22X1 U24644 ( .A(reg_A[41]), .B(n25242), .C(reg_A[40]), .D(n25338), .Y(
        n30062) );
  AOI22X1 U24645 ( .A(reg_A[43]), .B(n25339), .C(reg_A[42]), .D(n25257), .Y(
        n30061) );
  NOR2X1 U24646 ( .A(n30070), .B(n30071), .Y(n30048) );
  NAND3X1 U24647 ( .A(n30072), .B(n30073), .C(n30074), .Y(n30071) );
  NOR2X1 U24648 ( .A(n30075), .B(n30076), .Y(n30074) );
  OAI22X1 U24649 ( .A(n25043), .B(n30007), .C(n25039), .D(n30008), .Y(n30076)
         );
  OAI22X1 U24650 ( .A(n25064), .B(n30009), .C(n25482), .D(n29655), .Y(n30075)
         );
  AOI22X1 U24651 ( .A(reg_A[55]), .B(n25124), .C(reg_A[52]), .D(n25222), .Y(
        n30073) );
  AOI22X1 U24652 ( .A(reg_A[53]), .B(n25637), .C(reg_A[49]), .D(n25234), .Y(
        n30072) );
  NAND3X1 U24653 ( .A(n30077), .B(n30078), .C(n30079), .Y(n30070) );
  NOR2X1 U24654 ( .A(n30080), .B(n30081), .Y(n30079) );
  OAI22X1 U24655 ( .A(n25033), .B(n29990), .C(n25040), .D(n29989), .Y(n30081)
         );
  OAI22X1 U24656 ( .A(n25041), .B(n30015), .C(n25042), .D(n30016), .Y(n30080)
         );
  AOI22X1 U24657 ( .A(reg_A[56]), .B(n25628), .C(reg_A[59]), .D(n25069), .Y(
        n30078) );
  AOI22X1 U24658 ( .A(reg_A[58]), .B(n25123), .C(reg_A[54]), .D(n25629), .Y(
        n30077) );
  NOR2X1 U24659 ( .A(n30082), .B(n30083), .Y(n29951) );
  OAI21X1 U24660 ( .A(n30084), .B(n25697), .C(n30085), .Y(n30083) );
  OAI21X1 U24661 ( .A(n30086), .B(n30087), .C(n25999), .Y(n30085) );
  OAI21X1 U24662 ( .A(n26943), .B(n30007), .C(n30019), .Y(n30087) );
  NOR2X1 U24663 ( .A(n30088), .B(n30089), .Y(n30019) );
  OAI22X1 U24664 ( .A(n26944), .B(n26107), .C(n26945), .D(n25856), .Y(n30089)
         );
  OAI21X1 U24665 ( .A(n30090), .B(n30015), .C(n30091), .Y(n30088) );
  OAI21X1 U24666 ( .A(n25754), .B(n25851), .C(n30092), .Y(n30086) );
  AOI22X1 U24667 ( .A(reg_A[62]), .B(n26007), .C(reg_A[61]), .D(n26009), .Y(
        n30092) );
  INVX1 U24668 ( .A(n30093), .Y(n30084) );
  OAI21X1 U24669 ( .A(n30094), .B(n30095), .C(n30096), .Y(n30093) );
  AOI22X1 U24670 ( .A(n25097), .B(n30097), .C(n25604), .D(n30098), .Y(n30096)
         );
  OAI21X1 U24671 ( .A(n30099), .B(n30038), .C(n30100), .Y(n30098) );
  AOI22X1 U24672 ( .A(reg_B[60]), .B(n30101), .C(reg_B[63]), .D(n30102), .Y(
        n30100) );
  OAI22X1 U24673 ( .A(n30103), .B(n30043), .C(n30032), .D(n30009), .Y(n30101)
         );
  NAND2X1 U24674 ( .A(n30104), .B(n30105), .Y(n30097) );
  AOI22X1 U24675 ( .A(n29987), .B(n30106), .C(n30107), .D(n30108), .Y(n30105)
         );
  OAI21X1 U24676 ( .A(n30043), .B(n30109), .C(n30110), .Y(n30108) );
  AOI22X1 U24677 ( .A(n30111), .B(reg_A[39]), .C(n30112), .D(reg_A[47]), .Y(
        n30110) );
  INVX1 U24678 ( .A(n30113), .Y(n30106) );
  AOI21X1 U24679 ( .A(n30114), .B(reg_B[61]), .C(n30115), .Y(n30113) );
  AOI22X1 U24680 ( .A(n29991), .B(n30116), .C(n29981), .D(n30117), .Y(n30104)
         );
  OAI21X1 U24681 ( .A(n25994), .B(n30118), .C(n30119), .Y(n30082) );
  AOI22X1 U24682 ( .A(n30120), .B(n30121), .C(n30122), .D(n26260), .Y(n30119)
         );
  INVX1 U24683 ( .A(n30123), .Y(n30122) );
  NAND3X1 U24684 ( .A(n30124), .B(n30125), .C(n30126), .Y(result[62]) );
  NOR2X1 U24685 ( .A(n30127), .B(n30128), .Y(n30126) );
  NAND3X1 U24686 ( .A(n30129), .B(n30130), .C(n30131), .Y(n30128) );
  AOI22X1 U24687 ( .A(reg_A[59]), .B(n26161), .C(n30132), .D(n26139), .Y(
        n30131) );
  OAI21X1 U24688 ( .A(n30133), .B(n30134), .C(n25188), .Y(n30130) );
  OAI22X1 U24689 ( .A(n29973), .B(n30135), .C(n30136), .D(n30137), .Y(n30134)
         );
  OAI21X1 U24690 ( .A(n29989), .B(n30138), .C(n30139), .Y(n30133) );
  NAND3X1 U24691 ( .A(n30140), .B(reg_A[59]), .C(n30141), .Y(n30139) );
  AOI22X1 U24692 ( .A(n26045), .B(n30142), .C(reg_A[61]), .D(n27188), .Y(
        n30129) );
  NAND3X1 U24693 ( .A(n30143), .B(n30144), .C(n30145), .Y(n30142) );
  NOR2X1 U24694 ( .A(n30146), .B(n30147), .Y(n30145) );
  OAI21X1 U24695 ( .A(n25600), .B(n29990), .C(n30148), .Y(n30147) );
  AOI22X1 U24696 ( .A(reg_A[58]), .B(n25650), .C(reg_A[56]), .D(n25651), .Y(
        n30148) );
  OAI21X1 U24697 ( .A(n30149), .B(n29989), .C(n30150), .Y(n30146) );
  AOI22X1 U24698 ( .A(n25097), .B(n30151), .C(reg_A[62]), .D(n27639), .Y(
        n30150) );
  NAND3X1 U24699 ( .A(n30152), .B(n30153), .C(n30154), .Y(n30151) );
  AND2X1 U24700 ( .A(n30155), .B(n30156), .Y(n30154) );
  NOR2X1 U24701 ( .A(n30157), .B(n30158), .Y(n30156) );
  OAI21X1 U24702 ( .A(n25491), .B(n30059), .C(n30159), .Y(n30158) );
  AOI22X1 U24703 ( .A(reg_A[44]), .B(n25241), .C(reg_A[40]), .D(n25242), .Y(
        n30159) );
  OAI21X1 U24704 ( .A(n25038), .B(n30160), .C(n30161), .Y(n30157) );
  AOI22X1 U24705 ( .A(reg_A[45]), .B(n25246), .C(reg_A[46]), .D(n25247), .Y(
        n30161) );
  NOR2X1 U24706 ( .A(n30162), .B(n30163), .Y(n30155) );
  OAI21X1 U24707 ( .A(n25059), .B(n30058), .C(n30164), .Y(n30163) );
  AOI22X1 U24708 ( .A(reg_A[38]), .B(n25647), .C(reg_A[35]), .D(n25648), .Y(
        n30164) );
  OAI21X1 U24709 ( .A(n25054), .B(n30057), .C(n30165), .Y(n30162) );
  AOI22X1 U24710 ( .A(reg_A[42]), .B(n25339), .C(reg_A[41]), .D(n25257), .Y(
        n30165) );
  NOR2X1 U24711 ( .A(n30166), .B(n30167), .Y(n30153) );
  OAI21X1 U24712 ( .A(n25034), .B(n30168), .C(n30169), .Y(n30167) );
  AOI22X1 U24713 ( .A(reg_A[55]), .B(n25628), .C(reg_A[53]), .D(n25629), .Y(
        n30169) );
  OAI21X1 U24714 ( .A(n25498), .B(n30170), .C(n30171), .Y(n30166) );
  AOI22X1 U24715 ( .A(reg_A[32]), .B(n25631), .C(reg_A[34]), .D(n25324), .Y(
        n30171) );
  NOR2X1 U24716 ( .A(n30172), .B(n30173), .Y(n30152) );
  OAI21X1 U24717 ( .A(n25039), .B(n30174), .C(n30175), .Y(n30173) );
  AOI22X1 U24718 ( .A(reg_A[47]), .B(n25235), .C(reg_A[50]), .D(n25635), .Y(
        n30175) );
  OAI21X1 U24719 ( .A(n25035), .B(n29655), .C(n30176), .Y(n30172) );
  AOI22X1 U24720 ( .A(reg_A[51]), .B(n25222), .C(reg_A[52]), .D(n25637), .Y(
        n30176) );
  AOI21X1 U24721 ( .A(reg_A[67]), .B(n30177), .C(n30178), .Y(n30144) );
  OAI21X1 U24722 ( .A(n30179), .B(n25884), .C(n30180), .Y(n30178) );
  OAI21X1 U24723 ( .A(n30181), .B(n30182), .C(n25604), .Y(n30180) );
  NAND2X1 U24724 ( .A(n30183), .B(n30184), .Y(n30182) );
  AOI22X1 U24725 ( .A(reg_A[52]), .B(n25607), .C(reg_A[48]), .D(n25608), .Y(
        n30184) );
  AOI22X1 U24726 ( .A(reg_A[50]), .B(n25609), .C(reg_A[49]), .D(n25610), .Y(
        n30183) );
  NAND2X1 U24727 ( .A(n30185), .B(n30186), .Y(n30181) );
  AOI22X1 U24728 ( .A(reg_A[55]), .B(n25613), .C(reg_A[53]), .D(n25614), .Y(
        n30186) );
  AOI22X1 U24729 ( .A(reg_A[54]), .B(n25615), .C(reg_A[51]), .D(n25616), .Y(
        n30185) );
  AOI22X1 U24730 ( .A(reg_A[59]), .B(n27740), .C(reg_A[60]), .D(n27637), .Y(
        n30143) );
  NAND2X1 U24731 ( .A(n30187), .B(n30188), .Y(n30127) );
  AOI21X1 U24732 ( .A(reg_A[62]), .B(n30189), .C(n30190), .Y(n30188) );
  OAI21X1 U24733 ( .A(n30191), .B(n29998), .C(n30192), .Y(n30190) );
  OAI21X1 U24734 ( .A(n27183), .B(n30193), .C(reg_A[60]), .Y(n30192) );
  AOI22X1 U24735 ( .A(n30194), .B(n26601), .C(n30017), .D(n26597), .Y(n30191)
         );
  OAI21X1 U24736 ( .A(n29977), .B(n30103), .C(n30195), .Y(n30189) );
  AOI21X1 U24737 ( .A(n26267), .B(n30196), .C(n30197), .Y(n30187) );
  OAI22X1 U24738 ( .A(n30094), .B(n30198), .C(n26145), .D(n30199), .Y(n30197)
         );
  AOI21X1 U24739 ( .A(n30200), .B(n30201), .C(n30202), .Y(n30094) );
  INVX1 U24740 ( .A(n30203), .Y(n30202) );
  AOI22X1 U24741 ( .A(n30024), .B(n30204), .C(reg_B[62]), .D(n30205), .Y(
        n30203) );
  NAND2X1 U24742 ( .A(n30206), .B(n30207), .Y(n30204) );
  AOI22X1 U24743 ( .A(n30111), .B(reg_A[38]), .C(n30112), .D(reg_A[46]), .Y(
        n30207) );
  AOI22X1 U24744 ( .A(reg_A[62]), .B(n30117), .C(n30208), .D(reg_A[54]), .Y(
        n30206) );
  OAI21X1 U24745 ( .A(n30209), .B(n30210), .C(n30211), .Y(n30196) );
  AOI22X1 U24746 ( .A(n30102), .B(n30028), .C(n30212), .D(n30213), .Y(n30211)
         );
  NAND2X1 U24747 ( .A(n30214), .B(n30215), .Y(n30102) );
  MUX2X1 U24748 ( .B(n30216), .A(n30217), .S(reg_B[62]), .Y(n30215) );
  INVX1 U24749 ( .A(n30218), .Y(n30217) );
  NOR2X1 U24750 ( .A(n30219), .B(n30220), .Y(n30216) );
  AOI22X1 U24751 ( .A(reg_B[60]), .B(n30221), .C(n30222), .D(reg_A[62]), .Y(
        n30214) );
  OAI22X1 U24752 ( .A(n30223), .B(n30168), .C(n30008), .D(n30021), .Y(n30221)
         );
  NOR2X1 U24753 ( .A(n30224), .B(n30225), .Y(n30125) );
  OAI22X1 U24754 ( .A(n26525), .B(n30123), .C(n30226), .D(n26107), .Y(n30225)
         );
  OAI21X1 U24755 ( .A(n30227), .B(n26030), .C(n30228), .Y(n30123) );
  AOI22X1 U24756 ( .A(n26032), .B(n30229), .C(n25025), .D(n30230), .Y(n30228)
         );
  OAI21X1 U24757 ( .A(reg_A[62]), .B(n25063), .C(n30231), .Y(n30229) );
  AOI22X1 U24758 ( .A(n26038), .B(n30168), .C(reg_B[0]), .D(n30232), .Y(n30231) );
  OAI21X1 U24759 ( .A(n30233), .B(n30234), .C(n30235), .Y(n30224) );
  AOI22X1 U24760 ( .A(reg_A[63]), .B(n26408), .C(n30236), .D(n30121), .Y(
        n30235) );
  AOI21X1 U24761 ( .A(n30237), .B(n30201), .C(n30238), .Y(n30121) );
  INVX1 U24762 ( .A(n30239), .Y(n30238) );
  AOI22X1 U24763 ( .A(n30024), .B(n30240), .C(reg_B[62]), .D(n30241), .Y(
        n30239) );
  OAI21X1 U24764 ( .A(reg_A[54]), .B(n30109), .C(n30242), .Y(n30240) );
  AOI22X1 U24765 ( .A(reg_B[59]), .B(n30243), .C(n30117), .D(n30016), .Y(
        n30242) );
  NOR2X1 U24766 ( .A(n30244), .B(n30245), .Y(n30124) );
  NAND2X1 U24767 ( .A(n30246), .B(n30247), .Y(n30245) );
  MUX2X1 U24768 ( .B(n30042), .A(n30248), .S(reg_B[63]), .Y(n30246) );
  NOR2X1 U24769 ( .A(n28213), .B(n30249), .Y(n30248) );
  OAI21X1 U24770 ( .A(n30021), .B(n30250), .C(n30251), .Y(n30042) );
  OAI21X1 U24771 ( .A(n30252), .B(n30253), .C(n26186), .Y(n30251) );
  OAI22X1 U24772 ( .A(n30223), .B(n30016), .C(n30254), .D(n30255), .Y(n30253)
         );
  OAI22X1 U24773 ( .A(n30219), .B(n30021), .C(n30015), .D(n30256), .Y(n30252)
         );
  NAND2X1 U24774 ( .A(reg_A[58]), .B(n26504), .Y(n30250) );
  OAI21X1 U24775 ( .A(n30257), .B(n30258), .C(n30259), .Y(n30244) );
  AOI22X1 U24776 ( .A(n30260), .B(n26260), .C(n30261), .D(n30262), .Y(n30259)
         );
  OR2X1 U24777 ( .A(n30263), .B(n30264), .Y(result[61]) );
  NAND3X1 U24778 ( .A(n30265), .B(n30266), .C(n30267), .Y(n30264) );
  NOR2X1 U24779 ( .A(n30268), .B(n30269), .Y(n30267) );
  NAND2X1 U24780 ( .A(n30270), .B(n30247), .Y(n30269) );
  INVX1 U24781 ( .A(n30271), .Y(n30247) );
  OAI22X1 U24782 ( .A(n30255), .B(n30272), .C(n29998), .D(n30091), .Y(n30271)
         );
  MUX2X1 U24783 ( .B(n30031), .A(n30273), .S(reg_B[62]), .Y(n30270) );
  NOR2X1 U24784 ( .A(n25032), .B(n30274), .Y(n30273) );
  OAI22X1 U24785 ( .A(n30275), .B(n30276), .C(n25342), .D(n30277), .Y(n30031)
         );
  MUX2X1 U24786 ( .B(n30278), .A(n30279), .S(reg_B[61]), .Y(n30277) );
  MUX2X1 U24787 ( .B(n29990), .A(n30254), .S(reg_B[63]), .Y(n30279) );
  OAI21X1 U24788 ( .A(n30280), .B(n29973), .C(n25188), .Y(n30276) );
  OAI22X1 U24789 ( .A(n30281), .B(n30136), .C(n30278), .D(n29975), .Y(n30275)
         );
  MUX2X1 U24790 ( .B(n29989), .A(n30015), .S(reg_B[63]), .Y(n30278) );
  OAI21X1 U24791 ( .A(n30282), .B(n29989), .C(n30283), .Y(n30268) );
  AOI22X1 U24792 ( .A(n30284), .B(n26262), .C(n30285), .D(n30286), .Y(n30283)
         );
  AOI21X1 U24793 ( .A(reg_A[58]), .B(n30287), .C(n30288), .Y(n30266) );
  OAI22X1 U24794 ( .A(n30233), .B(n30289), .C(n30290), .D(n30234), .Y(n30288)
         );
  OAI21X1 U24795 ( .A(n30291), .B(n30255), .C(n30292), .Y(n30234) );
  AOI22X1 U24796 ( .A(n30037), .B(n30293), .C(n30141), .D(n30033), .Y(n30292)
         );
  NAND2X1 U24797 ( .A(n30294), .B(n30295), .Y(n30037) );
  AOI22X1 U24798 ( .A(n30041), .B(n30296), .C(reg_B[61]), .D(n30297), .Y(
        n30295) );
  AOI22X1 U24799 ( .A(n30298), .B(n29989), .C(n30039), .D(n30299), .Y(n30294)
         );
  AOI22X1 U24800 ( .A(n30260), .B(n26028), .C(n30300), .D(n26260), .Y(n30265)
         );
  INVX1 U24801 ( .A(n30301), .Y(n30260) );
  OAI21X1 U24802 ( .A(n30302), .B(n26208), .C(n30303), .Y(n30301) );
  AOI22X1 U24803 ( .A(n25026), .B(n29965), .C(n30304), .D(n26030), .Y(n30303)
         );
  INVX1 U24804 ( .A(n29962), .Y(n30304) );
  MUX2X1 U24805 ( .B(n30305), .A(n30306), .S(reg_B[2]), .Y(n29962) );
  OAI21X1 U24806 ( .A(reg_A[61]), .B(n25063), .C(n30307), .Y(n30305) );
  AOI22X1 U24807 ( .A(n26038), .B(n30299), .C(reg_B[0]), .D(n30308), .Y(n30307) );
  NAND3X1 U24808 ( .A(n30309), .B(n30310), .C(n30311), .Y(n30263) );
  NOR2X1 U24809 ( .A(n30312), .B(n30313), .Y(n30311) );
  OAI21X1 U24810 ( .A(n30314), .B(n30315), .C(n30316), .Y(n30313) );
  OAI21X1 U24811 ( .A(n30317), .B(n30318), .C(n26267), .Y(n30316) );
  OAI22X1 U24812 ( .A(n30319), .B(n30210), .C(n30209), .D(n30038), .Y(n30318)
         );
  OAI22X1 U24813 ( .A(n30218), .B(n30320), .C(n30099), .D(n29970), .Y(n30317)
         );
  INVX1 U24814 ( .A(n30213), .Y(n30099) );
  NAND2X1 U24815 ( .A(n30321), .B(n30322), .Y(n30213) );
  AOI22X1 U24816 ( .A(n30323), .B(reg_A[49]), .C(n30324), .D(reg_A[53]), .Y(
        n30322) );
  AOI22X1 U24817 ( .A(n30325), .B(reg_A[61]), .C(n30326), .D(reg_A[57]), .Y(
        n30321) );
  OAI21X1 U24818 ( .A(n30327), .B(n30328), .C(n30329), .Y(n30312) );
  AOI22X1 U24819 ( .A(n30330), .B(n30331), .C(n30332), .D(n26186), .Y(n30329)
         );
  NOR2X1 U24820 ( .A(reg_B[63]), .B(n30249), .Y(n30332) );
  INVX1 U24821 ( .A(n30333), .Y(n30249) );
  OAI21X1 U24822 ( .A(n30223), .B(n29989), .C(n30334), .Y(n30333) );
  AOI22X1 U24823 ( .A(n30141), .B(reg_A[59]), .C(n30201), .D(reg_A[57]), .Y(
        n30334) );
  MUX2X1 U24824 ( .B(n29984), .A(n30219), .S(reg_B[63]), .Y(n30331) );
  NOR2X1 U24825 ( .A(n25031), .B(n30256), .Y(n30330) );
  NAND2X1 U24826 ( .A(n25170), .B(n30262), .Y(n30328) );
  NAND2X1 U24827 ( .A(n30335), .B(n30336), .Y(n30262) );
  AOI22X1 U24828 ( .A(n30115), .B(n30293), .C(n30141), .D(n30116), .Y(n30336)
         );
  NAND2X1 U24829 ( .A(n30337), .B(n30338), .Y(n30115) );
  AOI22X1 U24830 ( .A(n30339), .B(n30324), .C(n30340), .D(reg_A[45]), .Y(
        n30338) );
  NOR2X1 U24831 ( .A(n30057), .B(n30341), .Y(n30339) );
  AOI22X1 U24832 ( .A(n30298), .B(reg_A[61]), .C(n30039), .D(reg_A[53]), .Y(
        n30337) );
  AOI22X1 U24833 ( .A(n30201), .B(n30114), .C(n30342), .D(n30343), .Y(n30335)
         );
  AOI21X1 U24834 ( .A(n30344), .B(n25150), .C(n30345), .Y(n30310) );
  OAI21X1 U24835 ( .A(n30346), .B(n29998), .C(n30347), .Y(n30345) );
  OAI21X1 U24836 ( .A(n30348), .B(n30349), .C(n26045), .Y(n30347) );
  NAND3X1 U24837 ( .A(n30350), .B(n30351), .C(n30352), .Y(n30349) );
  NOR2X1 U24838 ( .A(n30353), .B(n30354), .Y(n30352) );
  OAI22X1 U24839 ( .A(n27218), .B(n30015), .C(n30355), .D(n25884), .Y(n30354)
         );
  OAI21X1 U24840 ( .A(n30179), .B(n25855), .C(n30356), .Y(n30353) );
  AOI22X1 U24841 ( .A(reg_A[51]), .B(n25439), .C(reg_A[55]), .D(n25440), .Y(
        n30356) );
  AOI22X1 U24842 ( .A(reg_A[58]), .B(n25442), .C(reg_A[57]), .D(n27387), .Y(
        n30351) );
  AOI22X1 U24843 ( .A(reg_A[67]), .B(n30357), .C(reg_A[61]), .D(n25434), .Y(
        n30350) );
  NAND3X1 U24844 ( .A(n30358), .B(n30359), .C(n30360), .Y(n30348) );
  NOR2X1 U24845 ( .A(n30361), .B(n30362), .Y(n30360) );
  OAI22X1 U24846 ( .A(n25449), .B(n30254), .C(n25451), .D(n30174), .Y(n30362)
         );
  OAI21X1 U24847 ( .A(n25453), .B(n29655), .C(n30363), .Y(n30361) );
  AND2X1 U24848 ( .A(n30364), .B(n30365), .Y(n30363) );
  OAI21X1 U24849 ( .A(n30366), .B(n30367), .C(n25044), .Y(n30365) );
  NAND3X1 U24850 ( .A(n30368), .B(n30369), .C(n30370), .Y(n30367) );
  NOR2X1 U24851 ( .A(n30371), .B(n30372), .Y(n30370) );
  OAI21X1 U24852 ( .A(n25043), .B(n29989), .C(n30373), .Y(n30372) );
  AOI22X1 U24853 ( .A(reg_A[60]), .B(n25135), .C(reg_A[59]), .D(n25252), .Y(
        n30373) );
  NAND2X1 U24854 ( .A(n30374), .B(n30375), .Y(n30371) );
  AOI22X1 U24855 ( .A(reg_A[58]), .B(n25136), .C(reg_A[55]), .D(n25253), .Y(
        n30375) );
  AOI22X1 U24856 ( .A(reg_A[57]), .B(n25071), .C(reg_A[56]), .D(n25123), .Y(
        n30374) );
  NOR2X1 U24857 ( .A(n30376), .B(n30377), .Y(n30369) );
  OAI22X1 U24858 ( .A(n25034), .B(n30299), .C(n25030), .D(n30168), .Y(n30377)
         );
  OAI22X1 U24859 ( .A(n25036), .B(n30009), .C(n25037), .D(n30378), .Y(n30376)
         );
  NOR2X1 U24860 ( .A(n30379), .B(n30380), .Y(n30368) );
  OAI22X1 U24861 ( .A(n25064), .B(n30174), .C(n25473), .D(n30008), .Y(n30380)
         );
  OAI22X1 U24862 ( .A(n25039), .B(n29655), .C(n25475), .D(n30068), .Y(n30379)
         );
  NAND3X1 U24863 ( .A(n30381), .B(n30382), .C(n30383), .Y(n30366) );
  NOR2X1 U24864 ( .A(n30384), .B(n30385), .Y(n30383) );
  OAI21X1 U24865 ( .A(n25065), .B(n30069), .C(n30386), .Y(n30385) );
  AOI22X1 U24866 ( .A(reg_A[44]), .B(n25246), .C(reg_A[45]), .D(n25247), .Y(
        n30386) );
  NAND2X1 U24867 ( .A(n30387), .B(n30388), .Y(n30384) );
  AOI22X1 U24868 ( .A(reg_A[42]), .B(n25487), .C(reg_A[43]), .D(n25241), .Y(
        n30388) );
  AOI22X1 U24869 ( .A(reg_A[41]), .B(n25339), .C(reg_A[40]), .D(n25257), .Y(
        n30387) );
  NOR2X1 U24870 ( .A(n30389), .B(n30390), .Y(n30382) );
  OAI22X1 U24871 ( .A(n25491), .B(n30060), .C(n25492), .D(n30059), .Y(n30390)
         );
  OAI22X1 U24872 ( .A(n25057), .B(n30057), .C(n25322), .D(n30058), .Y(n30389)
         );
  NOR2X1 U24873 ( .A(n30391), .B(n30392), .Y(n30381) );
  OAI22X1 U24874 ( .A(n25059), .B(n30393), .C(n25318), .D(n30394), .Y(n30392)
         );
  OAI22X1 U24875 ( .A(n25498), .B(n30395), .C(n25499), .D(n30170), .Y(n30391)
         );
  OAI21X1 U24876 ( .A(n28312), .B(n27388), .C(reg_A[59]), .Y(n30364) );
  AOI22X1 U24877 ( .A(reg_A[52]), .B(n25500), .C(reg_A[53]), .D(n25501), .Y(
        n30359) );
  AOI22X1 U24878 ( .A(reg_A[54]), .B(n25502), .C(reg_A[50]), .D(n25503), .Y(
        n30358) );
  AOI21X1 U24879 ( .A(n30194), .B(n26597), .C(n30396), .Y(n30346) );
  INVX1 U24880 ( .A(n30397), .Y(n30396) );
  AOI22X1 U24881 ( .A(n27012), .B(n30017), .C(n26601), .D(n30398), .Y(n30397)
         );
  MUX2X1 U24882 ( .B(n29989), .A(n25851), .S(reg_B[2]), .Y(n30017) );
  INVX1 U24883 ( .A(n30118), .Y(n30344) );
  NAND2X1 U24884 ( .A(n30399), .B(n30400), .Y(n30118) );
  AOI22X1 U24885 ( .A(n26313), .B(n30015), .C(n26314), .D(n29989), .Y(n30400)
         );
  AOI22X1 U24886 ( .A(reg_B[1]), .B(n30401), .C(reg_B[2]), .D(n30402), .Y(
        n30399) );
  INVX1 U24887 ( .A(n30403), .Y(n30401) );
  AOI22X1 U24888 ( .A(reg_A[63]), .B(n26310), .C(reg_A[62]), .D(n26408), .Y(
        n30309) );
  NAND3X1 U24889 ( .A(n30404), .B(n30405), .C(n30406), .Y(result[60]) );
  NOR2X1 U24890 ( .A(n30407), .B(n30408), .Y(n30406) );
  NAND2X1 U24891 ( .A(n30409), .B(n30410), .Y(n30408) );
  AOI21X1 U24892 ( .A(reg_A[60]), .B(n30411), .C(n30412), .Y(n30410) );
  OAI21X1 U24893 ( .A(n29973), .B(n30272), .C(n30413), .Y(n30412) );
  OAI21X1 U24894 ( .A(n30414), .B(n30415), .C(n26267), .Y(n30413) );
  OAI22X1 U24895 ( .A(n30416), .B(n30210), .C(n30319), .D(n30038), .Y(n30415)
         );
  OAI22X1 U24896 ( .A(n30209), .B(n30320), .C(n30218), .D(n29970), .Y(n30414)
         );
  NOR2X1 U24897 ( .A(n30417), .B(n30418), .Y(n30218) );
  OAI22X1 U24898 ( .A(n30378), .B(n30136), .C(n30254), .D(n30220), .Y(n30418)
         );
  OAI21X1 U24899 ( .A(n30015), .B(n29975), .C(n30419), .Y(n30417) );
  OAI21X1 U24900 ( .A(n29977), .B(n30103), .C(n30420), .Y(n30411) );
  AOI21X1 U24901 ( .A(n27008), .B(n27012), .C(n26179), .Y(n30420) );
  INVX1 U24902 ( .A(n30421), .Y(n29977) );
  AOI21X1 U24903 ( .A(reg_A[57]), .B(n26161), .C(n30422), .Y(n30409) );
  NAND2X1 U24904 ( .A(n30423), .B(n30424), .Y(n30422) );
  OAI21X1 U24905 ( .A(n30425), .B(n30426), .C(n30427), .Y(n30424) );
  INVX1 U24906 ( .A(n30428), .Y(n30426) );
  AOI22X1 U24907 ( .A(n26597), .B(n30398), .C(n27012), .D(n30194), .Y(n30428)
         );
  MUX2X1 U24908 ( .B(n30015), .A(n25884), .S(reg_B[2]), .Y(n30194) );
  OAI21X1 U24909 ( .A(n27575), .B(n30429), .C(n30091), .Y(n30425) );
  NAND2X1 U24910 ( .A(reg_A[56]), .B(n26002), .Y(n30091) );
  OAI21X1 U24911 ( .A(n30430), .B(n30431), .C(n26045), .Y(n30423) );
  NAND3X1 U24912 ( .A(n30432), .B(n30433), .C(n30434), .Y(n30431) );
  NOR2X1 U24913 ( .A(n30435), .B(n30436), .Y(n30434) );
  OAI22X1 U24914 ( .A(n30437), .B(n29990), .C(n27218), .D(n29984), .Y(n30436)
         );
  OAI22X1 U24915 ( .A(n30355), .B(n25855), .C(n30179), .D(n25853), .Y(n30435)
         );
  AOI22X1 U24916 ( .A(reg_A[56]), .B(n27387), .C(reg_A[66]), .D(n30357), .Y(
        n30433) );
  AOI22X1 U24917 ( .A(reg_A[58]), .B(n28312), .C(reg_A[60]), .D(n25434), .Y(
        n30432) );
  NAND3X1 U24918 ( .A(n30438), .B(n30439), .C(n30440), .Y(n30430) );
  NOR2X1 U24919 ( .A(n30441), .B(n30442), .Y(n30440) );
  OAI22X1 U24920 ( .A(n30443), .B(n30299), .C(n30444), .D(n30378), .Y(n30442)
         );
  OAI21X1 U24921 ( .A(n26229), .B(n30009), .C(n30445), .Y(n30441) );
  AOI22X1 U24922 ( .A(reg_A[48]), .B(n28364), .C(reg_A[55]), .D(n30446), .Y(
        n30445) );
  AOI22X1 U24923 ( .A(reg_A[49]), .B(n25503), .C(reg_A[50]), .D(n25439), .Y(
        n30439) );
  AOI22X1 U24924 ( .A(reg_A[54]), .B(n25440), .C(n25097), .D(n30447), .Y(
        n30438) );
  NAND3X1 U24925 ( .A(n30448), .B(n30449), .C(n30450), .Y(n30447) );
  NOR2X1 U24926 ( .A(n30451), .B(n30452), .Y(n30450) );
  NAND3X1 U24927 ( .A(n30453), .B(n30454), .C(n30455), .Y(n30452) );
  AOI21X1 U24928 ( .A(reg_A[57]), .B(n25136), .C(n30456), .Y(n30455) );
  OAI22X1 U24929 ( .A(n25042), .B(n29984), .C(n25499), .D(n30395), .Y(n30456)
         );
  AOI22X1 U24930 ( .A(reg_A[35]), .B(n25857), .C(reg_A[36]), .D(n25647), .Y(
        n30454) );
  AOI22X1 U24931 ( .A(reg_A[33]), .B(n25648), .C(reg_A[34]), .D(n26432), .Y(
        n30453) );
  NAND3X1 U24932 ( .A(n30457), .B(n30458), .C(n30459), .Y(n30451) );
  NOR2X1 U24933 ( .A(n30460), .B(n30461), .Y(n30459) );
  OAI22X1 U24934 ( .A(n25051), .B(n30462), .C(n25243), .D(n30463), .Y(n30461)
         );
  OAI22X1 U24935 ( .A(n25334), .B(n30067), .C(n25336), .D(n30160), .Y(n30460)
         );
  AOI22X1 U24936 ( .A(reg_A[38]), .B(n25242), .C(reg_A[37]), .D(n25338), .Y(
        n30458) );
  AOI22X1 U24937 ( .A(reg_A[40]), .B(n25339), .C(reg_A[39]), .D(n25257), .Y(
        n30457) );
  NOR2X1 U24938 ( .A(n30464), .B(n30465), .Y(n30449) );
  OAI21X1 U24939 ( .A(n25034), .B(n30378), .C(n30466), .Y(n30465) );
  AOI22X1 U24940 ( .A(reg_A[55]), .B(n25123), .C(reg_A[51]), .D(n25629), .Y(
        n30466) );
  NAND2X1 U24941 ( .A(n30467), .B(n30468), .Y(n30464) );
  AOI22X1 U24942 ( .A(reg_A[58]), .B(n25252), .C(reg_A[54]), .D(n25253), .Y(
        n30468) );
  AOI22X1 U24943 ( .A(reg_A[53]), .B(n25628), .C(reg_A[56]), .D(n25068), .Y(
        n30467) );
  NOR2X1 U24944 ( .A(n30469), .B(n30470), .Y(n30448) );
  OAI21X1 U24945 ( .A(n25043), .B(n30015), .C(n30471), .Y(n30470) );
  AOI22X1 U24946 ( .A(reg_A[48]), .B(n25635), .C(reg_A[47]), .D(n25325), .Y(
        n30471) );
  NAND2X1 U24947 ( .A(n30472), .B(n30473), .Y(n30469) );
  AOI22X1 U24948 ( .A(reg_A[49]), .B(n25222), .C(reg_A[50]), .D(n25637), .Y(
        n30473) );
  AOI22X1 U24949 ( .A(reg_A[46]), .B(n25234), .C(reg_A[45]), .D(n25235), .Y(
        n30472) );
  NAND2X1 U24950 ( .A(n30474), .B(n30475), .Y(n30407) );
  AOI21X1 U24951 ( .A(reg_A[58]), .B(n30476), .C(n30477), .Y(n30475) );
  OAI21X1 U24952 ( .A(n30478), .B(n25794), .C(n30479), .Y(n30477) );
  NAND3X1 U24953 ( .A(reg_B[63]), .B(n30421), .C(n30480), .Y(n30479) );
  AOI22X1 U24954 ( .A(n30481), .B(n30324), .C(n30482), .D(n30326), .Y(n30478)
         );
  INVX1 U24955 ( .A(n30483), .Y(n30482) );
  INVX1 U24956 ( .A(n30484), .Y(n30476) );
  AOI21X1 U24957 ( .A(n26262), .B(n26314), .C(n30193), .Y(n30484) );
  OAI21X1 U24958 ( .A(n30256), .B(n30485), .C(n30486), .Y(n30193) );
  NAND2X1 U24959 ( .A(n30421), .B(n30028), .Y(n30485) );
  AOI21X1 U24960 ( .A(n30487), .B(n30488), .C(n30489), .Y(n30474) );
  OAI22X1 U24961 ( .A(n30314), .B(n30490), .C(n30491), .D(n29984), .Y(n30489)
         );
  AOI22X1 U24962 ( .A(n27008), .B(n26597), .C(n30492), .D(n30421), .Y(n30491)
         );
  OAI21X1 U24963 ( .A(reg_B[60]), .B(n25794), .C(n25031), .Y(n30421) );
  INVX1 U24964 ( .A(n30493), .Y(n30314) );
  OAI21X1 U24965 ( .A(n30494), .B(n30256), .C(n30495), .Y(n30493) );
  AOI22X1 U24966 ( .A(n25097), .B(n30496), .C(n25589), .D(n30497), .Y(n30495)
         );
  OAI22X1 U24967 ( .A(n30223), .B(n30015), .C(n30254), .D(n30021), .Y(n30497)
         );
  INVX1 U24968 ( .A(n30498), .Y(n30496) );
  AOI22X1 U24969 ( .A(n30499), .B(n30342), .C(n30293), .D(n30205), .Y(n30498)
         );
  NAND2X1 U24970 ( .A(n30500), .B(n30501), .Y(n30205) );
  AOI21X1 U24971 ( .A(n30340), .B(reg_A[44]), .C(n30502), .Y(n30501) );
  OAI21X1 U24972 ( .A(n30503), .B(n29973), .C(n30504), .Y(n30502) );
  NAND3X1 U24973 ( .A(reg_B[59]), .B(reg_A[36]), .C(n30324), .Y(n30504) );
  INVX1 U24974 ( .A(n30505), .Y(n30503) );
  AOI22X1 U24975 ( .A(n30298), .B(reg_A[60]), .C(n30039), .D(reg_A[52]), .Y(
        n30500) );
  NOR2X1 U24976 ( .A(n30506), .B(n30507), .Y(n30405) );
  OAI21X1 U24977 ( .A(n30290), .B(n30289), .C(n30508), .Y(n30507) );
  AOI22X1 U24978 ( .A(reg_A[62]), .B(n26310), .C(reg_A[61]), .D(n26408), .Y(
        n30508) );
  OAI21X1 U24979 ( .A(n30509), .B(n30255), .C(n30510), .Y(n30289) );
  AOI22X1 U24980 ( .A(n30241), .B(n30293), .C(n30141), .D(n30237), .Y(n30510)
         );
  NAND2X1 U24981 ( .A(n30511), .B(n30512), .Y(n30241) );
  AOI22X1 U24982 ( .A(n30041), .B(n30513), .C(reg_B[61]), .D(n30514), .Y(
        n30512) );
  NOR2X1 U24983 ( .A(n30341), .B(reg_B[61]), .Y(n30041) );
  AOI22X1 U24984 ( .A(n30298), .B(n30015), .C(n30039), .D(n30378), .Y(n30511)
         );
  OAI21X1 U24985 ( .A(n26418), .B(n30007), .C(n30515), .Y(n30506) );
  AOI22X1 U24986 ( .A(n30516), .B(n26139), .C(n30517), .D(n28575), .Y(n30515)
         );
  INVX1 U24987 ( .A(n30518), .Y(n30516) );
  NOR2X1 U24988 ( .A(n30519), .B(n30520), .Y(n30404) );
  OAI21X1 U24989 ( .A(n30258), .B(n30521), .C(n30522), .Y(n30520) );
  INVX1 U24990 ( .A(n30523), .Y(n30522) );
  INVX1 U24991 ( .A(n30286), .Y(n30258) );
  NAND2X1 U24992 ( .A(n30524), .B(n30525), .Y(n30286) );
  OAI21X1 U24993 ( .A(n26012), .B(n30526), .C(n30527), .Y(n30519) );
  AOI22X1 U24994 ( .A(n30528), .B(n30120), .C(n30300), .D(n26028), .Y(n30527)
         );
  INVX1 U24995 ( .A(n30529), .Y(n30300) );
  OAI21X1 U24996 ( .A(n30530), .B(n26208), .C(n30531), .Y(n30529) );
  AOI22X1 U24997 ( .A(n25026), .B(n30230), .C(n30532), .D(n26030), .Y(n30531)
         );
  INVX1 U24998 ( .A(n30227), .Y(n30532) );
  MUX2X1 U24999 ( .B(n30533), .A(n30534), .S(reg_B[2]), .Y(n30227) );
  OAI21X1 U25000 ( .A(reg_A[60]), .B(n25063), .C(n30535), .Y(n30533) );
  AOI22X1 U25001 ( .A(n26038), .B(n30378), .C(reg_B[0]), .D(n30536), .Y(n30535) );
  INVX1 U25002 ( .A(n30537), .Y(n30528) );
  NAND3X1 U25003 ( .A(n30538), .B(n30539), .C(n30540), .Y(result[5]) );
  NOR2X1 U25004 ( .A(n30541), .B(n30542), .Y(n30540) );
  NAND3X1 U25005 ( .A(n30543), .B(n26754), .C(n30544), .Y(n30542) );
  AOI21X1 U25006 ( .A(n29361), .B(reg_A[7]), .C(n30545), .Y(n30544) );
  OAI22X1 U25007 ( .A(n26677), .B(n25719), .C(n30546), .D(n30547), .Y(n30545)
         );
  INVX1 U25008 ( .A(n27969), .Y(n26754) );
  OAI21X1 U25009 ( .A(n30548), .B(n25794), .C(n25157), .Y(n27969) );
  MUX2X1 U25010 ( .B(n30549), .A(n30550), .S(reg_B[15]), .Y(n30543) );
  NOR2X1 U25011 ( .A(n27354), .B(n29301), .Y(n30549) );
  AOI22X1 U25012 ( .A(n29256), .B(n26735), .C(reg_A[3]), .D(n30551), .Y(n29301) );
  OAI22X1 U25013 ( .A(n29304), .B(n29265), .C(n30552), .D(n25177), .Y(n26735)
         );
  NAND3X1 U25014 ( .A(n30553), .B(n30554), .C(n30555), .Y(n30541) );
  AOI21X1 U25015 ( .A(n25730), .B(n30556), .C(n30557), .Y(n30555) );
  OAI21X1 U25016 ( .A(n30558), .B(n30559), .C(n30560), .Y(n30557) );
  OAI21X1 U25017 ( .A(n30561), .B(n30562), .C(n27358), .Y(n30560) );
  OAI21X1 U25018 ( .A(n29339), .B(n29265), .C(n30563), .Y(n30562) );
  AOI22X1 U25019 ( .A(reg_A[1]), .B(n25650), .C(reg_A[4]), .D(n29341), .Y(
        n30563) );
  NAND2X1 U25020 ( .A(n30564), .B(n30565), .Y(n30561) );
  AOI22X1 U25021 ( .A(n30566), .B(n29345), .C(reg_A[2]), .D(n29346), .Y(n30565) );
  INVX1 U25022 ( .A(n27963), .Y(n30566) );
  NAND2X1 U25023 ( .A(n30567), .B(n30568), .Y(n27963) );
  AOI22X1 U25024 ( .A(n26292), .B(n25177), .C(n26293), .D(n29265), .Y(n30568)
         );
  AOI22X1 U25025 ( .A(n26294), .B(n26742), .C(n26295), .D(n30569), .Y(n30567)
         );
  AOI22X1 U25026 ( .A(reg_A[3]), .B(n29349), .C(reg_A[0]), .D(n29350), .Y(
        n30564) );
  INVX1 U25027 ( .A(n30570), .Y(n30558) );
  NAND3X1 U25028 ( .A(n30571), .B(n30572), .C(n30573), .Y(n30556) );
  NOR2X1 U25029 ( .A(n30574), .B(n30575), .Y(n30573) );
  OAI21X1 U25030 ( .A(n25146), .B(n26801), .C(n30576), .Y(n30575) );
  AOI22X1 U25031 ( .A(reg_A[11]), .B(n26878), .C(n25613), .D(reg_A[12]), .Y(
        n30576) );
  OAI21X1 U25032 ( .A(n25132), .B(n25746), .C(n30577), .Y(n30574) );
  AOI22X1 U25033 ( .A(reg_A[6]), .B(n26803), .C(n26804), .D(reg_A[8]), .Y(
        n30577) );
  AOI21X1 U25034 ( .A(n25615), .B(reg_A[13]), .C(n30578), .Y(n30572) );
  OAI22X1 U25035 ( .A(n25208), .B(n27253), .C(n26800), .D(n25147), .Y(n30578)
         );
  AOI22X1 U25036 ( .A(n25607), .B(reg_A[15]), .C(n26924), .D(reg_A[5]), .Y(
        n30571) );
  OAI21X1 U25037 ( .A(n30579), .B(n30580), .C(n25310), .Y(n30554) );
  NAND3X1 U25038 ( .A(n30581), .B(n30582), .C(n30583), .Y(n30580) );
  NOR2X1 U25039 ( .A(n30584), .B(n30585), .Y(n30583) );
  OAI21X1 U25040 ( .A(n29265), .B(n25043), .C(n30586), .Y(n30585) );
  AOI22X1 U25041 ( .A(n25635), .B(reg_A[17]), .C(n25325), .D(reg_A[18]), .Y(
        n30586) );
  OAI21X1 U25042 ( .A(n30587), .B(n25482), .C(n30588), .Y(n30584) );
  AOI22X1 U25043 ( .A(n25637), .B(reg_A[15]), .C(n25234), .D(reg_A[19]), .Y(
        n30588) );
  NOR2X1 U25044 ( .A(n30589), .B(n30590), .Y(n30582) );
  OAI22X1 U25045 ( .A(n25147), .B(n26703), .C(n25146), .D(n26431), .Y(n30590)
         );
  OAI22X1 U25046 ( .A(n25255), .B(n25129), .C(n27967), .D(n25131), .Y(n30589)
         );
  AOI21X1 U25047 ( .A(n25222), .B(reg_A[16]), .C(n30591), .Y(n30581) );
  OAI22X1 U25048 ( .A(n25206), .B(n25467), .C(n25208), .D(n25223), .Y(n30591)
         );
  NAND3X1 U25049 ( .A(n30592), .B(n30593), .C(n30594), .Y(n30579) );
  NOR2X1 U25050 ( .A(n30595), .B(n30596), .Y(n30594) );
  OAI21X1 U25051 ( .A(n27960), .B(n25238), .C(n30597), .Y(n30596) );
  AOI22X1 U25052 ( .A(n25242), .B(reg_A[27]), .C(n25338), .D(reg_A[28]), .Y(
        n30597) );
  NAND2X1 U25053 ( .A(n30598), .B(n30599), .Y(n30595) );
  AOI22X1 U25054 ( .A(reg_A[22]), .B(n25246), .C(reg_A[21]), .D(n25247), .Y(
        n30599) );
  AOI22X1 U25055 ( .A(reg_A[24]), .B(n25487), .C(reg_A[23]), .D(n25241), .Y(
        n30598) );
  NOR2X1 U25056 ( .A(n30600), .B(n30601), .Y(n30593) );
  OAI22X1 U25057 ( .A(n27954), .B(n25316), .C(n25239), .D(n25320), .Y(n30601)
         );
  OAI22X1 U25058 ( .A(n29286), .B(n25322), .C(n27961), .D(n25049), .Y(n30600)
         );
  AOI21X1 U25059 ( .A(n25252), .B(reg_A[7]), .C(n30602), .Y(n30592) );
  OAI22X1 U25060 ( .A(n26701), .B(n25254), .C(n26677), .D(n25784), .Y(n30602)
         );
  AOI22X1 U25061 ( .A(reg_B[7]), .B(n30603), .C(reg_A[5]), .D(n29393), .Y(
        n30553) );
  NOR2X1 U25062 ( .A(n30604), .B(n30605), .Y(n30539) );
  OAI21X1 U25063 ( .A(n25177), .B(n29397), .C(n30606), .Y(n30605) );
  AOI22X1 U25064 ( .A(reg_A[3]), .B(n30607), .C(n30608), .D(n29314), .Y(n30606) );
  OAI21X1 U25065 ( .A(n25130), .B(n30609), .C(n30610), .Y(n29314) );
  AOI22X1 U25066 ( .A(n30611), .B(reg_B[5]), .C(n30612), .D(reg_A[5]), .Y(
        n30610) );
  NOR2X1 U25067 ( .A(reg_B[6]), .B(n25177), .Y(n30611) );
  NAND2X1 U25068 ( .A(n29513), .B(n29322), .Y(n30607) );
  NAND3X1 U25069 ( .A(n26504), .B(n28041), .C(n30613), .Y(n29322) );
  NAND3X1 U25070 ( .A(n30614), .B(n29312), .C(n30615), .Y(n30604) );
  OAI21X1 U25071 ( .A(n30616), .B(n30617), .C(n29306), .Y(n30615) );
  MUX2X1 U25072 ( .B(n30618), .A(n30619), .S(reg_B[30]), .Y(n29306) );
  NAND2X1 U25073 ( .A(n25110), .B(reg_A[3]), .Y(n30619) );
  INVX1 U25074 ( .A(n26762), .Y(n30618) );
  OAI21X1 U25075 ( .A(n28033), .B(n25177), .C(n30620), .Y(n26762) );
  NAND3X1 U25076 ( .A(reg_B[5]), .B(reg_A[0]), .C(n30621), .Y(n29312) );
  NAND3X1 U25077 ( .A(n26504), .B(n28005), .C(n28011), .Y(n30614) );
  MUX2X1 U25078 ( .B(n30622), .A(n30623), .S(reg_B[7]), .Y(n28011) );
  MUX2X1 U25079 ( .B(reg_A[5]), .A(reg_A[1]), .S(reg_B[5]), .Y(n30622) );
  NOR2X1 U25080 ( .A(n30624), .B(n30625), .Y(n30538) );
  OAI21X1 U25081 ( .A(n30626), .B(n25128), .C(n30627), .Y(n30625) );
  OAI21X1 U25082 ( .A(n30628), .B(n30629), .C(n25382), .Y(n30627) );
  OAI22X1 U25083 ( .A(n25092), .B(n28026), .C(n30630), .D(n30631), .Y(n30629)
         );
  INVX1 U25084 ( .A(n30632), .Y(n30628) );
  AOI22X1 U25085 ( .A(n30633), .B(n27984), .C(n25090), .D(n28038), .Y(n30632)
         );
  AOI21X1 U25086 ( .A(n30634), .B(n25110), .C(n30635), .Y(n30626) );
  OAI21X1 U25087 ( .A(n25194), .B(n26727), .C(n30636), .Y(n30635) );
  NAND3X1 U25088 ( .A(n30637), .B(n30638), .C(n30639), .Y(n30624) );
  INVX1 U25089 ( .A(n30640), .Y(n30639) );
  AOI21X1 U25090 ( .A(n30641), .B(n30642), .C(n26996), .Y(n30640) );
  AOI22X1 U25091 ( .A(n30643), .B(n26772), .C(n25102), .D(n30644), .Y(n30642)
         );
  AOI22X1 U25092 ( .A(n25111), .B(n25101), .C(n30645), .D(reg_B[27]), .Y(
        n30641) );
  OAI21X1 U25093 ( .A(n30646), .B(n30647), .C(reg_A[0]), .Y(n30638) );
  OAI21X1 U25094 ( .A(n27438), .B(n30648), .C(n30649), .Y(n30647) );
  NOR2X1 U25095 ( .A(n25116), .B(n28057), .Y(n30646) );
  OAI21X1 U25096 ( .A(n30650), .B(n30651), .C(reg_A[4]), .Y(n30637) );
  OR2X1 U25097 ( .A(n25173), .B(n29502), .Y(n30651) );
  NAND3X1 U25098 ( .A(n30652), .B(n30653), .C(n30654), .Y(result[59]) );
  NOR2X1 U25099 ( .A(n30655), .B(n30656), .Y(n30654) );
  NAND3X1 U25100 ( .A(n30657), .B(n30658), .C(n30659), .Y(n30656) );
  AOI22X1 U25101 ( .A(n30427), .B(n30660), .C(reg_A[59]), .D(n30661), .Y(
        n30659) );
  OAI21X1 U25102 ( .A(n27454), .B(n30429), .C(n30662), .Y(n30660) );
  AOI22X1 U25103 ( .A(n30663), .B(n26601), .C(n30398), .D(n27012), .Y(n30662)
         );
  MUX2X1 U25104 ( .B(n29984), .A(n25855), .S(reg_B[2]), .Y(n30398) );
  INVX1 U25105 ( .A(n30664), .Y(n30429) );
  OAI21X1 U25106 ( .A(n30665), .B(n30666), .C(n26267), .Y(n30658) );
  OAI22X1 U25107 ( .A(n30667), .B(n30210), .C(n30416), .D(n30038), .Y(n30666)
         );
  OAI22X1 U25108 ( .A(n30319), .B(n30320), .C(n30209), .D(n29970), .Y(n30665)
         );
  INVX1 U25109 ( .A(n30668), .Y(n30209) );
  OAI21X1 U25110 ( .A(n30043), .B(n30220), .C(n30669), .Y(n30668) );
  AOI22X1 U25111 ( .A(n30324), .B(reg_A[51]), .C(n30325), .D(reg_A[59]), .Y(
        n30669) );
  AOI22X1 U25112 ( .A(reg_A[63]), .B(n26482), .C(n26504), .D(n30670), .Y(
        n30657) );
  OAI21X1 U25113 ( .A(n30219), .B(n29978), .C(n30671), .Y(n30670) );
  AOI22X1 U25114 ( .A(n30480), .B(n30028), .C(reg_A[56]), .D(n30672), .Y(
        n30671) );
  NAND2X1 U25115 ( .A(n30673), .B(n30674), .Y(n30655) );
  AOI21X1 U25116 ( .A(n30675), .B(n25188), .C(n30676), .Y(n30674) );
  OAI21X1 U25117 ( .A(n30677), .B(n30678), .C(n30679), .Y(n30676) );
  AOI22X1 U25118 ( .A(n25382), .B(n30680), .C(n30117), .D(n26480), .Y(n30678)
         );
  MUX2X1 U25119 ( .B(n30274), .A(n30681), .S(reg_B[62]), .Y(n30675) );
  OAI21X1 U25120 ( .A(n30023), .B(n30220), .C(n30682), .Y(n30274) );
  AOI21X1 U25121 ( .A(n30020), .B(n29973), .C(n30683), .Y(n30682) );
  INVX1 U25122 ( .A(n30684), .Y(n30020) );
  MUX2X1 U25123 ( .B(n30685), .A(n30686), .S(reg_B[63]), .Y(n30684) );
  MUX2X1 U25124 ( .B(reg_A[59]), .A(reg_A[51]), .S(reg_B[60]), .Y(n30685) );
  AOI22X1 U25125 ( .A(n30687), .B(n30488), .C(n30487), .D(n30688), .Y(n30673)
         );
  INVX1 U25126 ( .A(n30315), .Y(n30487) );
  NAND2X1 U25127 ( .A(reg_B[63]), .B(n25170), .Y(n30315) );
  OAI21X1 U25128 ( .A(n30689), .B(n26999), .C(n30690), .Y(n30488) );
  INVX1 U25129 ( .A(n30691), .Y(n30690) );
  AOI21X1 U25130 ( .A(n30692), .B(n30693), .C(n25403), .Y(n30691) );
  AOI22X1 U25131 ( .A(n30694), .B(n30342), .C(n30343), .D(n30201), .Y(n30693)
         );
  AOI22X1 U25132 ( .A(n30114), .B(n30141), .C(n30116), .D(n30024), .Y(n30692)
         );
  NAND2X1 U25133 ( .A(n30695), .B(n30696), .Y(n30116) );
  AOI22X1 U25134 ( .A(n30111), .B(reg_A[35]), .C(n30112), .D(reg_A[43]), .Y(
        n30696) );
  AOI22X1 U25135 ( .A(n30117), .B(reg_A[59]), .C(n30208), .D(reg_A[51]), .Y(
        n30695) );
  AOI21X1 U25136 ( .A(n30024), .B(reg_A[59]), .C(n30480), .Y(n30689) );
  NOR2X1 U25137 ( .A(n30256), .B(n29990), .Y(n30480) );
  NOR2X1 U25138 ( .A(n30697), .B(n30698), .Y(n30653) );
  OAI22X1 U25139 ( .A(n30290), .B(n30537), .C(n26136), .D(n30015), .Y(n30698)
         );
  NAND2X1 U25140 ( .A(n30699), .B(n30700), .Y(n30537) );
  AOI22X1 U25141 ( .A(n30024), .B(n30033), .C(n30141), .D(n30297), .Y(n30700)
         );
  OAI21X1 U25142 ( .A(reg_A[51]), .B(n30109), .C(n30701), .Y(n30033) );
  AOI22X1 U25143 ( .A(reg_B[59]), .B(n30702), .C(n30117), .D(n29984), .Y(
        n30701) );
  AOI22X1 U25144 ( .A(n30201), .B(n30703), .C(n30342), .D(n30704), .Y(n30699)
         );
  OAI21X1 U25145 ( .A(n26812), .B(n29989), .C(n30705), .Y(n30697) );
  AOI22X1 U25146 ( .A(reg_A[62]), .B(n26451), .C(n30284), .D(n25150), .Y(
        n30705) );
  INVX1 U25147 ( .A(n30706), .Y(n30284) );
  OAI21X1 U25148 ( .A(reg_B[2]), .B(n29961), .C(n30707), .Y(n30706) );
  AOI22X1 U25149 ( .A(n26455), .B(n29655), .C(n26456), .D(n29959), .Y(n30707)
         );
  AND2X1 U25150 ( .A(n30708), .B(n30709), .Y(n29961) );
  AOI22X1 U25151 ( .A(n26460), .B(n30009), .C(n26461), .D(n29984), .Y(n30709)
         );
  AOI22X1 U25152 ( .A(n26462), .B(n30219), .C(n26463), .D(n30008), .Y(n30708)
         );
  NOR2X1 U25153 ( .A(n30710), .B(n30711), .Y(n30652) );
  OAI21X1 U25154 ( .A(n25994), .B(n30712), .C(n30713), .Y(n30711) );
  OAI21X1 U25155 ( .A(n30714), .B(n30715), .C(n26045), .Y(n30713) );
  NAND3X1 U25156 ( .A(n30716), .B(n30717), .C(n30718), .Y(n30715) );
  NOR2X1 U25157 ( .A(n30719), .B(n30720), .Y(n30718) );
  OAI22X1 U25158 ( .A(n27755), .B(n30299), .C(n27756), .D(n30043), .Y(n30720)
         );
  OAI22X1 U25159 ( .A(n30149), .B(n30219), .C(n25619), .D(n29984), .Y(n30719)
         );
  INVX1 U25160 ( .A(n25617), .Y(n30149) );
  AOI22X1 U25161 ( .A(reg_A[54]), .B(n30721), .C(reg_A[63]), .D(n30722), .Y(
        n30717) );
  AOI22X1 U25162 ( .A(reg_A[64]), .B(n30177), .C(reg_A[65]), .D(n30357), .Y(
        n30716) );
  NAND3X1 U25163 ( .A(n30723), .B(n30724), .C(n30725), .Y(n30714) );
  NOR2X1 U25164 ( .A(n30726), .B(n30727), .Y(n30725) );
  OAI21X1 U25165 ( .A(n28362), .B(n30174), .C(n30728), .Y(n30727) );
  OAI21X1 U25166 ( .A(n30729), .B(n30730), .C(n25044), .Y(n30728) );
  NAND3X1 U25167 ( .A(n30731), .B(n30732), .C(n30733), .Y(n30730) );
  NOR2X1 U25168 ( .A(n30734), .B(n30735), .Y(n30733) );
  OAI22X1 U25169 ( .A(n25473), .B(n29655), .C(n25467), .D(n30009), .Y(n30735)
         );
  OAI21X1 U25170 ( .A(n25037), .B(n30008), .C(n30736), .Y(n30734) );
  AOI22X1 U25171 ( .A(reg_A[33]), .B(n26432), .C(reg_A[52]), .D(n25628), .Y(
        n30736) );
  AOI21X1 U25172 ( .A(reg_A[44]), .B(n25235), .C(n30737), .Y(n30732) );
  OAI22X1 U25173 ( .A(n25035), .B(n30066), .C(n25219), .D(n30174), .Y(n30737)
         );
  AOI22X1 U25174 ( .A(reg_A[47]), .B(n25635), .C(reg_A[46]), .D(n25325), .Y(
        n30731) );
  NAND3X1 U25175 ( .A(n30738), .B(n30739), .C(n30740), .Y(n30729) );
  NOR2X1 U25176 ( .A(n30741), .B(n30742), .Y(n30740) );
  OAI21X1 U25177 ( .A(n25491), .B(n30058), .C(n30743), .Y(n30742) );
  AOI22X1 U25178 ( .A(reg_A[41]), .B(n25241), .C(reg_A[37]), .D(n25242), .Y(
        n30743) );
  OAI21X1 U25179 ( .A(n25038), .B(n30744), .C(n30745), .Y(n30741) );
  AOI22X1 U25180 ( .A(reg_A[42]), .B(n25246), .C(reg_A[43]), .D(n25247), .Y(
        n30745) );
  AOI21X1 U25181 ( .A(reg_A[34]), .B(n25857), .C(n30746), .Y(n30739) );
  OAI22X1 U25182 ( .A(n26719), .B(n30060), .C(n25238), .D(n30059), .Y(n30746)
         );
  AOI22X1 U25183 ( .A(reg_A[35]), .B(n25647), .C(reg_A[32]), .D(n25648), .Y(
        n30738) );
  OAI22X1 U25184 ( .A(n28363), .B(n29655), .C(n30443), .D(n30378), .Y(n30726)
         );
  AOI22X1 U25185 ( .A(reg_A[56]), .B(n29346), .C(reg_A[57]), .D(n29349), .Y(
        n30724) );
  AOI22X1 U25186 ( .A(reg_A[50]), .B(n25500), .C(reg_A[51]), .D(n25501), .Y(
        n30723) );
  OAI21X1 U25187 ( .A(n26012), .B(n30747), .C(n30748), .Y(n30710) );
  INVX1 U25188 ( .A(n30749), .Y(n30748) );
  OAI22X1 U25189 ( .A(n30750), .B(n30233), .C(n30526), .D(n26525), .Y(n30749)
         );
  NAND2X1 U25190 ( .A(n30751), .B(n30752), .Y(n30526) );
  AOI22X1 U25191 ( .A(n25025), .B(n30753), .C(n25026), .D(n30306), .Y(n30752)
         );
  AOI22X1 U25192 ( .A(n26032), .B(n29965), .C(n26530), .D(n30754), .Y(n30751)
         );
  OAI21X1 U25193 ( .A(reg_A[59]), .B(n25063), .C(n30755), .Y(n29965) );
  AOI22X1 U25194 ( .A(n26038), .B(n30009), .C(reg_B[0]), .D(n30756), .Y(n30755) );
  OR2X1 U25195 ( .A(n30757), .B(n30758), .Y(result[58]) );
  NAND3X1 U25196 ( .A(n30759), .B(n30760), .C(n30761), .Y(n30758) );
  NOR2X1 U25197 ( .A(n30762), .B(n30763), .Y(n30761) );
  OAI21X1 U25198 ( .A(n26136), .B(n29984), .C(n30764), .Y(n30763) );
  AOI22X1 U25199 ( .A(reg_A[61]), .B(n26451), .C(reg_A[60]), .D(n26310), .Y(
        n30764) );
  OAI21X1 U25200 ( .A(n26420), .B(n30765), .C(n30766), .Y(n30762) );
  AOI22X1 U25201 ( .A(reg_A[58]), .B(n30661), .C(reg_A[62]), .D(n30767), .Y(
        n30766) );
  OAI21X1 U25202 ( .A(n25031), .B(n30103), .C(n30282), .Y(n30661) );
  AOI21X1 U25203 ( .A(n30768), .B(n26028), .C(n30769), .Y(n30760) );
  OAI22X1 U25204 ( .A(n30233), .B(n30770), .C(n30290), .D(n30750), .Y(n30769)
         );
  NAND2X1 U25205 ( .A(n30771), .B(n30772), .Y(n30750) );
  AOI22X1 U25206 ( .A(n30024), .B(n30237), .C(n30141), .D(n30514), .Y(n30772)
         );
  NAND2X1 U25207 ( .A(n30773), .B(n30774), .Y(n30237) );
  AOI22X1 U25208 ( .A(n30111), .B(n30394), .C(n30112), .D(n30462), .Y(n30774)
         );
  AOI22X1 U25209 ( .A(n30117), .B(n30219), .C(n30208), .D(n30008), .Y(n30773)
         );
  AOI22X1 U25210 ( .A(n30201), .B(n30775), .C(n30342), .D(n30776), .Y(n30771)
         );
  INVX1 U25211 ( .A(n30747), .Y(n30768) );
  NAND2X1 U25212 ( .A(n30777), .B(n30778), .Y(n30747) );
  AOI22X1 U25213 ( .A(n25025), .B(n30779), .C(n25026), .D(n30534), .Y(n30778)
         );
  AOI22X1 U25214 ( .A(n26032), .B(n30230), .C(n26530), .D(n30780), .Y(n30777)
         );
  NAND2X1 U25215 ( .A(n30781), .B(n30782), .Y(n30230) );
  AOI22X1 U25216 ( .A(n26662), .B(n30394), .C(n26663), .D(n30462), .Y(n30782)
         );
  AOI22X1 U25217 ( .A(n26038), .B(n30008), .C(n26664), .D(n30219), .Y(n30781)
         );
  NOR2X1 U25218 ( .A(n30523), .B(n30783), .Y(n30759) );
  OAI21X1 U25219 ( .A(n26012), .B(n30784), .C(n30785), .Y(n30783) );
  OAI21X1 U25220 ( .A(n30786), .B(n30787), .C(n26045), .Y(n30785) );
  NAND2X1 U25221 ( .A(n30788), .B(n30789), .Y(n30787) );
  AOI22X1 U25222 ( .A(reg_A[57]), .B(n30790), .C(reg_A[64]), .D(n30357), .Y(
        n30789) );
  INVX1 U25223 ( .A(n30791), .Y(n30790) );
  AOI22X1 U25224 ( .A(reg_A[56]), .B(n27388), .C(reg_A[58]), .D(n30792), .Y(
        n30788) );
  NAND2X1 U25225 ( .A(n30793), .B(n30794), .Y(n30786) );
  AOI22X1 U25226 ( .A(n25097), .B(n30795), .C(n25604), .D(n30796), .Y(n30794)
         );
  NAND3X1 U25227 ( .A(n30797), .B(n30798), .C(n30799), .Y(n30796) );
  NOR2X1 U25228 ( .A(n30800), .B(n30801), .Y(n30799) );
  OAI21X1 U25229 ( .A(n26801), .B(n30168), .C(n30802), .Y(n30801) );
  AOI22X1 U25230 ( .A(reg_A[52]), .B(n26878), .C(reg_A[51]), .D(n25613), .Y(
        n30802) );
  OAI21X1 U25231 ( .A(n25746), .B(n30254), .C(n30803), .Y(n30800) );
  AOI22X1 U25232 ( .A(reg_A[57]), .B(n26803), .C(reg_A[55]), .D(n26804), .Y(
        n30803) );
  AOI21X1 U25233 ( .A(reg_A[50]), .B(n25615), .C(n30804), .Y(n30798) );
  OAI22X1 U25234 ( .A(n27253), .B(n30174), .C(n26800), .D(n30299), .Y(n30804)
         );
  AOI22X1 U25235 ( .A(reg_A[48]), .B(n25607), .C(reg_A[58]), .D(n26924), .Y(
        n30797) );
  NAND3X1 U25236 ( .A(n30805), .B(n30806), .C(n30807), .Y(n30795) );
  NOR2X1 U25237 ( .A(n30808), .B(n30809), .Y(n30807) );
  NAND3X1 U25238 ( .A(n30810), .B(n30811), .C(n30812), .Y(n30809) );
  AOI21X1 U25239 ( .A(reg_A[56]), .B(n25252), .C(n30813), .Y(n30812) );
  OAI22X1 U25240 ( .A(n25041), .B(n30043), .C(n25042), .D(n29990), .Y(n30813)
         );
  AOI22X1 U25241 ( .A(reg_A[37]), .B(n25257), .C(reg_A[33]), .D(n25857), .Y(
        n30811) );
  AOI22X1 U25242 ( .A(reg_A[34]), .B(n25647), .C(reg_A[32]), .D(n26432), .Y(
        n30810) );
  NAND3X1 U25243 ( .A(n30814), .B(n30815), .C(n30816), .Y(n30808) );
  AOI21X1 U25244 ( .A(reg_A[38]), .B(n25339), .C(n30817), .Y(n30816) );
  OAI22X1 U25245 ( .A(n25491), .B(n30393), .C(n25492), .D(n30058), .Y(n30817)
         );
  AOI22X1 U25246 ( .A(reg_A[41]), .B(n25246), .C(reg_A[42]), .D(n25247), .Y(
        n30815) );
  AOI22X1 U25247 ( .A(reg_A[39]), .B(n25487), .C(reg_A[40]), .D(n25241), .Y(
        n30814) );
  NOR2X1 U25248 ( .A(n30818), .B(n30819), .Y(n30806) );
  OAI21X1 U25249 ( .A(n25473), .B(n30068), .C(n30820), .Y(n30819) );
  AOI22X1 U25250 ( .A(reg_A[49]), .B(n25629), .C(reg_A[50]), .D(n25124), .Y(
        n30820) );
  NAND2X1 U25251 ( .A(n30821), .B(n30822), .Y(n30818) );
  AOI22X1 U25252 ( .A(reg_A[52]), .B(n25253), .C(reg_A[51]), .D(n25628), .Y(
        n30822) );
  AOI22X1 U25253 ( .A(reg_A[54]), .B(n25071), .C(reg_A[53]), .D(n25123), .Y(
        n30821) );
  NOR2X1 U25254 ( .A(n30823), .B(n30824), .Y(n30805) );
  OAI21X1 U25255 ( .A(n25043), .B(n30219), .C(n30825), .Y(n30824) );
  AOI22X1 U25256 ( .A(reg_A[46]), .B(n25635), .C(reg_A[45]), .D(n25325), .Y(
        n30825) );
  OAI21X1 U25257 ( .A(n25065), .B(n30160), .C(n30826), .Y(n30823) );
  AOI22X1 U25258 ( .A(reg_A[48]), .B(n25637), .C(reg_A[44]), .D(n25234), .Y(
        n30826) );
  AOI22X1 U25259 ( .A(reg_A[62]), .B(n30722), .C(reg_A[63]), .D(n30177), .Y(
        n30793) );
  OAI22X1 U25260 ( .A(n25794), .B(n30419), .C(n29655), .D(n30827), .Y(n30523)
         );
  NAND2X1 U25261 ( .A(n30828), .B(reg_B[61]), .Y(n30419) );
  NAND3X1 U25262 ( .A(n30829), .B(n30830), .C(n30831), .Y(n30757) );
  NOR2X1 U25263 ( .A(n30832), .B(n30833), .Y(n30831) );
  OAI21X1 U25264 ( .A(n26584), .B(n30199), .C(n30834), .Y(n30833) );
  AOI22X1 U25265 ( .A(n25188), .B(n30835), .C(n30687), .D(n30688), .Y(n30834)
         );
  OAI21X1 U25266 ( .A(n30494), .B(n30223), .C(n30836), .Y(n30688) );
  AOI22X1 U25267 ( .A(n30837), .B(n30141), .C(n25097), .D(n30838), .Y(n30836)
         );
  OAI21X1 U25268 ( .A(n30839), .B(n30255), .C(n30840), .Y(n30838) );
  AOI22X1 U25269 ( .A(n30141), .B(n30505), .C(n30201), .D(n30499), .Y(n30840)
         );
  INVX1 U25270 ( .A(n30841), .Y(n30839) );
  NOR2X1 U25271 ( .A(n26999), .B(n30254), .Y(n30837) );
  AOI22X1 U25272 ( .A(n25589), .B(reg_A[58]), .C(n30200), .D(n25097), .Y(
        n30494) );
  NAND2X1 U25273 ( .A(n30842), .B(n30843), .Y(n30200) );
  AOI22X1 U25274 ( .A(n30111), .B(reg_A[34]), .C(reg_A[58]), .D(n30117), .Y(
        n30843) );
  AOI22X1 U25275 ( .A(n30208), .B(reg_A[50]), .C(n30112), .D(reg_A[42]), .Y(
        n30842) );
  INVX1 U25276 ( .A(n30490), .Y(n30687) );
  NAND2X1 U25277 ( .A(n25170), .B(n30028), .Y(n30490) );
  OAI22X1 U25278 ( .A(reg_B[61]), .B(n30135), .C(n30220), .D(n30137), .Y(
        n30835) );
  NAND2X1 U25279 ( .A(n30844), .B(n30845), .Y(n30137) );
  AOI22X1 U25280 ( .A(n30846), .B(n30168), .C(n30212), .D(n30299), .Y(n30845)
         );
  AOI22X1 U25281 ( .A(n29987), .B(n30378), .C(n30847), .D(n30009), .Y(n30844)
         );
  NAND2X1 U25282 ( .A(n30848), .B(n30849), .Y(n30135) );
  MUX2X1 U25283 ( .B(n30850), .A(n30851), .S(reg_B[60]), .Y(n30849) );
  NOR2X1 U25284 ( .A(reg_A[48]), .B(n30293), .Y(n30851) );
  OAI22X1 U25285 ( .A(reg_A[55]), .B(n30210), .C(reg_A[56]), .D(n30038), .Y(
        n30850) );
  AOI22X1 U25286 ( .A(n30846), .B(n30686), .C(n30212), .D(n30852), .Y(n30848)
         );
  MUX2X1 U25287 ( .B(reg_A[50]), .A(reg_A[58]), .S(n30853), .Y(n30686) );
  NAND2X1 U25288 ( .A(n30854), .B(n30855), .Y(n30199) );
  AOI22X1 U25289 ( .A(n26593), .B(n30008), .C(n26594), .D(n29655), .Y(n30855)
         );
  AOI22X1 U25290 ( .A(n30856), .B(n26596), .C(n26597), .D(n30857), .Y(n30854)
         );
  OAI21X1 U25291 ( .A(reg_A[58]), .B(n26599), .C(n30858), .Y(n30856) );
  AOI22X1 U25292 ( .A(n26601), .B(n30254), .C(n26602), .D(n30043), .Y(n30858)
         );
  OAI21X1 U25293 ( .A(n29978), .B(n30859), .C(n30860), .Y(n30832) );
  AOI21X1 U25294 ( .A(n30861), .B(n30862), .C(n30863), .Y(n30860) );
  INVX1 U25295 ( .A(n30679), .Y(n30863) );
  AND2X1 U25296 ( .A(n30864), .B(n25170), .Y(n30861) );
  NAND2X1 U25297 ( .A(reg_A[57]), .B(n29315), .Y(n30859) );
  AOI21X1 U25298 ( .A(reg_A[63]), .B(n30865), .C(n30866), .Y(n30830) );
  OAI22X1 U25299 ( .A(n30024), .B(n30272), .C(n30257), .D(n30867), .Y(n30866)
         );
  NAND2X1 U25300 ( .A(reg_A[56]), .B(n26504), .Y(n30272) );
  AOI21X1 U25301 ( .A(n30427), .B(n30868), .C(n30869), .Y(n30829) );
  OAI21X1 U25302 ( .A(n30870), .B(n30871), .C(n30872), .Y(n30869) );
  OAI21X1 U25303 ( .A(n30873), .B(n30874), .C(n26267), .Y(n30872) );
  OAI22X1 U25304 ( .A(n30875), .B(n30210), .C(n30667), .D(n30038), .Y(n30874)
         );
  OAI22X1 U25305 ( .A(n30416), .B(n30320), .C(n30319), .D(n29970), .Y(n30873)
         );
  INVX1 U25306 ( .A(n30876), .Y(n30319) );
  OAI21X1 U25307 ( .A(n30168), .B(n30220), .C(n30877), .Y(n30876) );
  AOI22X1 U25308 ( .A(n30324), .B(reg_A[50]), .C(n30325), .D(reg_A[58]), .Y(
        n30877) );
  OAI21X1 U25309 ( .A(n27454), .B(n30878), .C(n30879), .Y(n30868) );
  AOI22X1 U25310 ( .A(reg_A[56]), .B(n25026), .C(n30664), .D(n27012), .Y(
        n30879) );
  MUX2X1 U25311 ( .B(n30219), .A(n25853), .S(reg_B[2]), .Y(n30664) );
  NAND3X1 U25312 ( .A(n30880), .B(n30881), .C(n30882), .Y(result[57]) );
  NOR2X1 U25313 ( .A(n30883), .B(n30884), .Y(n30882) );
  NAND2X1 U25314 ( .A(n30885), .B(n30886), .Y(n30884) );
  NOR2X1 U25315 ( .A(n30887), .B(n30888), .Y(n30886) );
  OAI21X1 U25316 ( .A(n30871), .B(n30889), .C(n30890), .Y(n30888) );
  OAI21X1 U25317 ( .A(n30891), .B(n30892), .C(n25188), .Y(n30890) );
  OAI21X1 U25318 ( .A(n30038), .B(n30893), .C(n30894), .Y(n30892) );
  INVX1 U25319 ( .A(n30895), .Y(n30894) );
  MUX2X1 U25320 ( .B(n30681), .A(n30896), .S(reg_B[62]), .Y(n30895) );
  OAI21X1 U25321 ( .A(reg_B[61]), .B(n30280), .C(n30897), .Y(n30681) );
  AOI21X1 U25322 ( .A(n30326), .B(n30898), .C(n30683), .Y(n30897) );
  AND2X1 U25323 ( .A(n30323), .B(n29655), .Y(n30683) );
  INVX1 U25324 ( .A(n30281), .Y(n30898) );
  MUX2X1 U25325 ( .B(n30299), .A(n30378), .S(reg_B[63]), .Y(n30281) );
  AOI21X1 U25326 ( .A(n30254), .B(n30140), .C(n30899), .Y(n30280) );
  INVX1 U25327 ( .A(n30900), .Y(n30899) );
  MUX2X1 U25328 ( .B(n30852), .A(n30901), .S(reg_B[63]), .Y(n30900) );
  NOR2X1 U25329 ( .A(reg_A[48]), .B(n30853), .Y(n30901) );
  MUX2X1 U25330 ( .B(reg_A[49]), .A(reg_A[57]), .S(n30853), .Y(n30852) );
  OAI21X1 U25331 ( .A(n30255), .B(n30902), .C(n30903), .Y(n30891) );
  NAND3X1 U25332 ( .A(n30023), .B(n30853), .C(n30141), .Y(n30903) );
  MUX2X1 U25333 ( .B(n30043), .A(n30168), .S(reg_B[63]), .Y(n30023) );
  NAND2X1 U25334 ( .A(n30140), .B(reg_A[50]), .Y(n30902) );
  NOR2X1 U25335 ( .A(n30028), .B(reg_B[60]), .Y(n30140) );
  INVX1 U25336 ( .A(n30904), .Y(n30871) );
  OAI21X1 U25337 ( .A(n26881), .B(n29959), .C(n30905), .Y(n30887) );
  OAI21X1 U25338 ( .A(n30906), .B(n30907), .C(reg_A[57]), .Y(n30905) );
  NAND2X1 U25339 ( .A(n30908), .B(n30282), .Y(n30907) );
  NOR2X1 U25340 ( .A(n28213), .B(n30103), .Y(n30906) );
  INVX1 U25341 ( .A(n30909), .Y(n29959) );
  AOI21X1 U25342 ( .A(n30910), .B(n30911), .C(n30912), .Y(n30885) );
  OAI21X1 U25343 ( .A(n30913), .B(n29655), .C(n30914), .Y(n30912) );
  OAI21X1 U25344 ( .A(n30915), .B(n30916), .C(reg_A[56]), .Y(n30914) );
  OAI22X1 U25345 ( .A(n27523), .B(n30791), .C(n30107), .D(n25342), .Y(n30916)
         );
  OAI21X1 U25346 ( .A(n26151), .B(n29978), .C(n30917), .Y(n30915) );
  OAI21X1 U25347 ( .A(n26295), .B(n25026), .C(n30427), .Y(n30917) );
  NAND2X1 U25348 ( .A(n30918), .B(n30919), .Y(n30883) );
  NOR2X1 U25349 ( .A(n30920), .B(n30921), .Y(n30919) );
  OAI21X1 U25350 ( .A(n30922), .B(n29989), .C(n30923), .Y(n30921) );
  OAI21X1 U25351 ( .A(n30865), .B(n28282), .C(reg_A[62]), .Y(n30923) );
  AOI21X1 U25352 ( .A(n30722), .B(n26045), .C(n30767), .Y(n30922) );
  OAI21X1 U25353 ( .A(n25754), .B(n29998), .C(n30924), .Y(n30767) );
  OAI21X1 U25354 ( .A(n30878), .B(n30925), .C(n30679), .Y(n30920) );
  NAND2X1 U25355 ( .A(n27012), .B(n30427), .Y(n30925) );
  INVX1 U25356 ( .A(n30663), .Y(n30878) );
  MUX2X1 U25357 ( .B(n29990), .A(n30007), .S(reg_B[2]), .Y(n30663) );
  AOI21X1 U25358 ( .A(n30926), .B(n30285), .C(n30927), .Y(n30918) );
  OAI21X1 U25359 ( .A(n30928), .B(n25697), .C(n30929), .Y(n30927) );
  NAND2X1 U25360 ( .A(reg_A[63]), .B(n30930), .Y(n30929) );
  OAI21X1 U25361 ( .A(n26894), .B(n30931), .C(n30932), .Y(n30930) );
  AOI21X1 U25362 ( .A(n30933), .B(n30864), .C(n30934), .Y(n30928) );
  OAI21X1 U25363 ( .A(n30935), .B(n30095), .C(n30936), .Y(n30934) );
  OAI21X1 U25364 ( .A(n30937), .B(n30938), .C(n25604), .Y(n30936) );
  OAI22X1 U25365 ( .A(n30939), .B(n30210), .C(n30875), .D(n30038), .Y(n30938)
         );
  OAI22X1 U25366 ( .A(n30667), .B(n30320), .C(n30416), .D(n29970), .Y(n30937)
         );
  INVX1 U25367 ( .A(n30940), .Y(n30416) );
  OAI21X1 U25368 ( .A(n30299), .B(n30220), .C(n30941), .Y(n30940) );
  AOI22X1 U25369 ( .A(n30324), .B(reg_A[49]), .C(n30325), .D(reg_A[57]), .Y(
        n30941) );
  INVX1 U25370 ( .A(n30942), .Y(n30935) );
  NAND2X1 U25371 ( .A(n30943), .B(n30944), .Y(n30864) );
  AOI22X1 U25372 ( .A(n30024), .B(n30114), .C(n30141), .D(n30343), .Y(n30944)
         );
  NAND2X1 U25373 ( .A(n30945), .B(n30946), .Y(n30114) );
  AOI22X1 U25374 ( .A(n30111), .B(reg_A[33]), .C(n30112), .D(reg_A[41]), .Y(
        n30946) );
  AOI22X1 U25375 ( .A(reg_A[57]), .B(n30117), .C(n30208), .D(reg_A[49]), .Y(
        n30945) );
  AOI22X1 U25376 ( .A(n30201), .B(n30694), .C(n30342), .D(n30947), .Y(n30943)
         );
  NOR2X1 U25377 ( .A(n30948), .B(n30949), .Y(n30881) );
  OAI21X1 U25378 ( .A(n30950), .B(n30951), .C(n30952), .Y(n30949) );
  INVX1 U25379 ( .A(n30953), .Y(n30952) );
  OAI22X1 U25380 ( .A(n30770), .B(n30290), .C(n30954), .D(n30233), .Y(n30953)
         );
  NAND2X1 U25381 ( .A(n30955), .B(n30956), .Y(n30770) );
  AOI22X1 U25382 ( .A(n30024), .B(n30297), .C(n30141), .D(n30703), .Y(n30956)
         );
  INVX1 U25383 ( .A(n30291), .Y(n30703) );
  NAND2X1 U25384 ( .A(n30957), .B(n30958), .Y(n30297) );
  AOI22X1 U25385 ( .A(n30111), .B(n30170), .C(n30112), .D(n30463), .Y(n30958)
         );
  AOI22X1 U25386 ( .A(n30117), .B(n29990), .C(n30208), .D(n30174), .Y(n30957)
         );
  AOI22X1 U25387 ( .A(n30201), .B(n30704), .C(n30342), .D(n30959), .Y(n30955)
         );
  INVX1 U25388 ( .A(n30960), .Y(n30959) );
  NOR2X1 U25389 ( .A(n30961), .B(n30962), .Y(n30950) );
  NAND3X1 U25390 ( .A(n30963), .B(n30964), .C(n30965), .Y(n30962) );
  NOR2X1 U25391 ( .A(n30966), .B(n30967), .Y(n30965) );
  OAI21X1 U25392 ( .A(n25037), .B(n29655), .C(n30968), .Y(n30967) );
  AOI22X1 U25393 ( .A(reg_A[53]), .B(n25072), .C(reg_A[52]), .D(n25123), .Y(
        n30968) );
  OAI21X1 U25394 ( .A(n25030), .B(n30008), .C(n30969), .Y(n30966) );
  AOI22X1 U25395 ( .A(reg_A[55]), .B(n25252), .C(reg_A[51]), .D(n25253), .Y(
        n30969) );
  AOI21X1 U25396 ( .A(reg_A[43]), .B(n25234), .C(n30970), .Y(n30964) );
  OAI22X1 U25397 ( .A(n25036), .B(n30068), .C(n25467), .D(n30174), .Y(n30970)
         );
  AOI22X1 U25398 ( .A(reg_A[44]), .B(n25325), .C(reg_A[57]), .D(n25125), .Y(
        n30963) );
  NAND2X1 U25399 ( .A(n30971), .B(n30972), .Y(n30961) );
  NOR2X1 U25400 ( .A(n30973), .B(n30974), .Y(n30972) );
  OAI21X1 U25401 ( .A(n25050), .B(n30394), .C(n30975), .Y(n30974) );
  AOI22X1 U25402 ( .A(reg_A[39]), .B(n25241), .C(reg_A[35]), .D(n25242), .Y(
        n30975) );
  OAI21X1 U25403 ( .A(n25038), .B(n30060), .C(n30976), .Y(n30973) );
  AOI22X1 U25404 ( .A(reg_A[40]), .B(n25246), .C(reg_A[41]), .D(n25247), .Y(
        n30976) );
  NOR2X1 U25405 ( .A(n30977), .B(n30978), .Y(n30971) );
  OAI21X1 U25406 ( .A(n25041), .B(n30168), .C(n30979), .Y(n30978) );
  AOI22X1 U25407 ( .A(reg_A[33]), .B(n25647), .C(reg_A[56]), .D(n25135), .Y(
        n30979) );
  OAI21X1 U25408 ( .A(n25054), .B(n30395), .C(n30980), .Y(n30977) );
  AOI22X1 U25409 ( .A(reg_A[37]), .B(n25339), .C(reg_A[36]), .D(n25257), .Y(
        n30980) );
  NAND2X1 U25410 ( .A(n30981), .B(n30982), .Y(n30948) );
  AOI22X1 U25411 ( .A(reg_A[60]), .B(n26451), .C(n30983), .D(n25150), .Y(
        n30982) );
  INVX1 U25412 ( .A(n30712), .Y(n30983) );
  NAND2X1 U25413 ( .A(n30984), .B(n30985), .Y(n30712) );
  AOI22X1 U25414 ( .A(n26859), .B(n30378), .C(n26860), .D(n30299), .Y(n30985)
         );
  AOI22X1 U25415 ( .A(n26455), .B(n29655), .C(n30402), .D(n26452), .Y(n30984)
         );
  OAI21X1 U25416 ( .A(reg_A[48]), .B(n26861), .C(n30986), .Y(n30402) );
  AOI22X1 U25417 ( .A(n30857), .B(n26863), .C(n26462), .D(n30254), .Y(n30986)
         );
  MUX2X1 U25418 ( .B(reg_A[49]), .A(reg_A[57]), .S(n26596), .Y(n30857) );
  AOI22X1 U25419 ( .A(reg_A[59]), .B(n26310), .C(reg_A[58]), .D(n26408), .Y(
        n30981) );
  NOR2X1 U25420 ( .A(n30987), .B(n30988), .Y(n30880) );
  OAI21X1 U25421 ( .A(n30989), .B(n30990), .C(n30991), .Y(n30988) );
  AOI22X1 U25422 ( .A(reg_A[45]), .B(n26519), .C(reg_A[42]), .D(n26349), .Y(
        n30991) );
  AND2X1 U25423 ( .A(n30992), .B(n30993), .Y(n30989) );
  NOR2X1 U25424 ( .A(n30994), .B(n30995), .Y(n30993) );
  OAI22X1 U25425 ( .A(n26800), .B(n30378), .C(n26801), .D(n30299), .Y(n30995)
         );
  OAI21X1 U25426 ( .A(n25062), .B(n30043), .C(n30996), .Y(n30994) );
  AOI22X1 U25427 ( .A(reg_A[56]), .B(n26803), .C(reg_A[54]), .D(n26804), .Y(
        n30996) );
  NOR2X1 U25428 ( .A(n30997), .B(n30998), .Y(n30992) );
  OAI21X1 U25429 ( .A(n25060), .B(n29990), .C(n30999), .Y(n30998) );
  INVX1 U25430 ( .A(n30911), .Y(n30999) );
  OAI22X1 U25431 ( .A(n26936), .B(n30008), .C(n25745), .D(n30009), .Y(n30911)
         );
  OAI22X1 U25432 ( .A(n27252), .B(n30174), .C(n27253), .D(n29655), .Y(n30997)
         );
  OAI21X1 U25433 ( .A(n31000), .B(n30069), .C(n31001), .Y(n30987) );
  AOI22X1 U25434 ( .A(n31002), .B(n26028), .C(n31003), .D(n26260), .Y(n31001)
         );
  INVX1 U25435 ( .A(n30784), .Y(n31002) );
  NAND2X1 U25436 ( .A(n31004), .B(n31005), .Y(n30784) );
  AOI22X1 U25437 ( .A(n25025), .B(n30754), .C(n25026), .D(n30753), .Y(n31005)
         );
  AOI22X1 U25438 ( .A(n26032), .B(n30306), .C(n26530), .D(n31006), .Y(n31004)
         );
  NAND2X1 U25439 ( .A(n31007), .B(n31008), .Y(n30306) );
  AOI22X1 U25440 ( .A(n26662), .B(n30170), .C(n26663), .D(n30463), .Y(n31008)
         );
  AOI22X1 U25441 ( .A(n26038), .B(n30174), .C(n26664), .D(n29990), .Y(n31007)
         );
  NAND3X1 U25442 ( .A(n31009), .B(n31010), .C(n31011), .Y(result[56]) );
  NOR2X1 U25443 ( .A(n31012), .B(n31013), .Y(n31011) );
  NAND3X1 U25444 ( .A(n31014), .B(n31015), .C(n31016), .Y(n31013) );
  AOI21X1 U25445 ( .A(n31017), .B(n30120), .C(n31018), .Y(n31016) );
  OAI22X1 U25446 ( .A(n30290), .B(n30954), .C(n26420), .D(n30518), .Y(n31018)
         );
  NAND2X1 U25447 ( .A(n31019), .B(n31020), .Y(n30954) );
  AOI22X1 U25448 ( .A(n30024), .B(n30514), .C(n30141), .D(n30775), .Y(n31020)
         );
  OR2X1 U25449 ( .A(n31021), .B(n31022), .Y(n30514) );
  OAI22X1 U25450 ( .A(reg_A[48]), .B(n30109), .C(reg_A[56]), .D(n29994), .Y(
        n31022) );
  OAI21X1 U25451 ( .A(reg_A[40]), .B(n31023), .C(n31024), .Y(n31021) );
  AOI22X1 U25452 ( .A(n30201), .B(n30776), .C(n30342), .D(n31025), .Y(n31019)
         );
  OAI21X1 U25453 ( .A(n31026), .B(n31027), .C(n25310), .Y(n31015) );
  NAND2X1 U25454 ( .A(n31028), .B(n31029), .Y(n31027) );
  AOI22X1 U25455 ( .A(reg_A[63]), .B(n25628), .C(reg_A[60]), .D(n25068), .Y(
        n31029) );
  AOI22X1 U25456 ( .A(reg_A[61]), .B(n25123), .C(reg_A[56]), .D(n25125), .Y(
        n31028) );
  NAND2X1 U25457 ( .A(n31030), .B(n31031), .Y(n31026) );
  AOI22X1 U25458 ( .A(reg_A[57]), .B(n25135), .C(reg_A[59]), .D(n25136), .Y(
        n31031) );
  AOI22X1 U25459 ( .A(reg_A[58]), .B(n25252), .C(reg_A[62]), .D(n25253), .Y(
        n31030) );
  AOI22X1 U25460 ( .A(n31032), .B(n30904), .C(n25188), .D(n31033), .Y(n31014)
         );
  OAI21X1 U25461 ( .A(n29975), .B(n30483), .C(n31034), .Y(n31033) );
  AOI21X1 U25462 ( .A(n30481), .B(n30326), .C(n30828), .Y(n31034) );
  INVX1 U25463 ( .A(n30896), .Y(n30828) );
  AND2X1 U25464 ( .A(n31035), .B(n31036), .Y(n30481) );
  AOI22X1 U25465 ( .A(n30846), .B(n30378), .C(n30212), .D(n30009), .Y(n31036)
         );
  AOI22X1 U25466 ( .A(n29987), .B(n30008), .C(n30847), .D(n30174), .Y(n31035)
         );
  NAND2X1 U25467 ( .A(n31037), .B(n31038), .Y(n30483) );
  AOI22X1 U25468 ( .A(n30846), .B(n30254), .C(n30212), .D(n30043), .Y(n31038)
         );
  AOI22X1 U25469 ( .A(n29987), .B(n30168), .C(n30847), .D(n30299), .Y(n31037)
         );
  OAI21X1 U25470 ( .A(n31039), .B(n31040), .C(n30525), .Y(n30904) );
  NAND3X1 U25471 ( .A(n30680), .B(n29973), .C(n25382), .Y(n30525) );
  NAND2X1 U25472 ( .A(n30325), .B(n25382), .Y(n31040) );
  NAND3X1 U25473 ( .A(n31041), .B(n31042), .C(n31043), .Y(n31012) );
  AOI21X1 U25474 ( .A(n30926), .B(n31044), .C(n31045), .Y(n31043) );
  OAI21X1 U25475 ( .A(n31046), .B(n30254), .C(n30679), .Y(n31045) );
  NAND3X1 U25476 ( .A(n30427), .B(n26602), .C(reg_A[56]), .Y(n30679) );
  NOR2X1 U25477 ( .A(n31047), .B(n31048), .Y(n31046) );
  OAI21X1 U25478 ( .A(n26151), .B(n30103), .C(n27190), .Y(n31048) );
  NAND2X1 U25479 ( .A(n30908), .B(n25031), .Y(n31047) );
  INVX1 U25480 ( .A(n30867), .Y(n30926) );
  NAND2X1 U25481 ( .A(n25382), .B(n31049), .Y(n30867) );
  OAI22X1 U25482 ( .A(n30220), .B(n31039), .C(n29993), .D(n29973), .Y(n31049)
         );
  INVX1 U25483 ( .A(n30680), .Y(n29993) );
  OAI21X1 U25484 ( .A(reg_B[60]), .B(n25415), .C(n26999), .Y(n30680) );
  OAI21X1 U25485 ( .A(n31050), .B(n31051), .C(n26267), .Y(n31042) );
  OAI22X1 U25486 ( .A(n31052), .B(n30210), .C(n30939), .D(n30038), .Y(n31051)
         );
  INVX1 U25487 ( .A(n31053), .Y(n30939) );
  OAI22X1 U25488 ( .A(n30875), .B(n30320), .C(n30667), .D(n29970), .Y(n31050)
         );
  INVX1 U25489 ( .A(n31054), .Y(n30667) );
  OAI21X1 U25490 ( .A(n30378), .B(n30220), .C(n31055), .Y(n31054) );
  AOI22X1 U25491 ( .A(n30324), .B(reg_A[48]), .C(n30325), .D(reg_A[56]), .Y(
        n31055) );
  INVX1 U25492 ( .A(n31056), .Y(n30875) );
  AOI22X1 U25493 ( .A(n30517), .B(n27008), .C(n31057), .D(n29565), .Y(n31041)
         );
  OAI21X1 U25494 ( .A(n31058), .B(n30016), .C(n31059), .Y(n31057) );
  AOI22X1 U25495 ( .A(reg_A[60]), .B(n30722), .C(reg_A[61]), .D(n30177), .Y(
        n31059) );
  AND2X1 U25496 ( .A(n31060), .B(n31061), .Y(n30517) );
  AOI22X1 U25497 ( .A(n26601), .B(n30168), .C(n26602), .D(n30299), .Y(n31061)
         );
  AOI22X1 U25498 ( .A(n27012), .B(n30254), .C(n26597), .D(n30043), .Y(n31060)
         );
  NOR2X1 U25499 ( .A(n31062), .B(n31063), .Y(n31010) );
  OAI21X1 U25500 ( .A(n26985), .B(n29655), .C(n31064), .Y(n31063) );
  AOI22X1 U25501 ( .A(n31003), .B(n26028), .C(n31065), .D(n26260), .Y(n31064)
         );
  INVX1 U25502 ( .A(n31066), .Y(n31065) );
  AND2X1 U25503 ( .A(n31067), .B(n31068), .Y(n31003) );
  AOI22X1 U25504 ( .A(n25025), .B(n30780), .C(n25026), .D(n30779), .Y(n31068)
         );
  AOI22X1 U25505 ( .A(n26032), .B(n30534), .C(n26530), .D(n31069), .Y(n31067)
         );
  OR2X1 U25506 ( .A(n31070), .B(n31071), .Y(n30534) );
  OAI22X1 U25507 ( .A(reg_A[56]), .B(n26036), .C(reg_A[48]), .D(n26981), .Y(
        n31071) );
  OAI21X1 U25508 ( .A(reg_A[40]), .B(n26982), .C(n31072), .Y(n31070) );
  OAI21X1 U25509 ( .A(n31073), .B(n30951), .C(n31074), .Y(n31062) );
  AOI22X1 U25510 ( .A(n30261), .B(n31075), .C(n31076), .D(n30942), .Y(n31074)
         );
  NAND2X1 U25511 ( .A(n31077), .B(n31078), .Y(n30942) );
  AOI22X1 U25512 ( .A(n30024), .B(n30505), .C(n30141), .D(n30499), .Y(n31078)
         );
  NAND2X1 U25513 ( .A(n31079), .B(n31080), .Y(n30505) );
  AOI22X1 U25514 ( .A(n30111), .B(reg_A[32]), .C(n30112), .D(reg_A[40]), .Y(
        n31080) );
  AOI22X1 U25515 ( .A(reg_A[56]), .B(n30117), .C(n30208), .D(reg_A[48]), .Y(
        n31079) );
  AOI22X1 U25516 ( .A(n30201), .B(n30841), .C(n30342), .D(n31081), .Y(n31077)
         );
  NOR2X1 U25517 ( .A(n31082), .B(n31083), .Y(n31073) );
  NAND3X1 U25518 ( .A(n31084), .B(n31085), .C(n31086), .Y(n31083) );
  NOR2X1 U25519 ( .A(n31087), .B(n31088), .Y(n31086) );
  OAI21X1 U25520 ( .A(n25037), .B(n30068), .C(n31089), .Y(n31088) );
  AOI22X1 U25521 ( .A(reg_A[52]), .B(n25072), .C(reg_A[51]), .D(n25123), .Y(
        n31089) );
  OAI21X1 U25522 ( .A(n25030), .B(n30174), .C(n31090), .Y(n31087) );
  AOI22X1 U25523 ( .A(reg_A[54]), .B(n25252), .C(reg_A[50]), .D(n25253), .Y(
        n31090) );
  AOI21X1 U25524 ( .A(reg_A[42]), .B(n25234), .C(n31091), .Y(n31085) );
  OAI22X1 U25525 ( .A(n25036), .B(n30069), .C(n25467), .D(n29655), .Y(n31091)
         );
  AOI22X1 U25526 ( .A(reg_A[43]), .B(n25325), .C(reg_A[56]), .D(n25125), .Y(
        n31084) );
  NAND3X1 U25527 ( .A(n31092), .B(n31093), .C(n31094), .Y(n31082) );
  NOR2X1 U25528 ( .A(n31095), .B(n31096), .Y(n31094) );
  OAI21X1 U25529 ( .A(n25050), .B(n30170), .C(n31097), .Y(n31096) );
  AOI22X1 U25530 ( .A(reg_A[38]), .B(n25241), .C(reg_A[34]), .D(n25242), .Y(
        n31097) );
  OAI21X1 U25531 ( .A(n25038), .B(n30057), .C(n31098), .Y(n31095) );
  AOI22X1 U25532 ( .A(reg_A[39]), .B(n25246), .C(reg_A[40]), .D(n25247), .Y(
        n31098) );
  AOI21X1 U25533 ( .A(reg_A[32]), .B(n25647), .C(n31099), .Y(n31093) );
  OAI22X1 U25534 ( .A(n26719), .B(n30393), .C(n25238), .D(n30058), .Y(n31099)
         );
  AOI22X1 U25535 ( .A(reg_A[55]), .B(n25135), .C(reg_A[53]), .D(n25136), .Y(
        n31092) );
  NOR2X1 U25536 ( .A(n31100), .B(n31101), .Y(n31009) );
  OAI21X1 U25537 ( .A(n31102), .B(n27152), .C(n31103), .Y(n31101) );
  AOI22X1 U25538 ( .A(n26928), .B(n31104), .C(n25918), .D(n31105), .Y(n31103)
         );
  NAND3X1 U25539 ( .A(n31106), .B(n31107), .C(n31108), .Y(n31105) );
  NOR2X1 U25540 ( .A(n31109), .B(n31110), .Y(n31108) );
  OAI22X1 U25541 ( .A(n26936), .B(n30174), .C(n25745), .D(n30008), .Y(n31110)
         );
  OAI21X1 U25542 ( .A(n25062), .B(n30168), .C(n31111), .Y(n31109) );
  AOI22X1 U25543 ( .A(reg_A[55]), .B(n26803), .C(reg_A[53]), .D(n26804), .Y(
        n31111) );
  AOI22X1 U25544 ( .A(reg_A[52]), .B(n25749), .C(reg_A[51]), .D(n25750), .Y(
        n31107) );
  AOI22X1 U25545 ( .A(reg_A[48]), .B(n25615), .C(reg_A[56]), .D(n26924), .Y(
        n31106) );
  NAND3X1 U25546 ( .A(n31112), .B(n31113), .C(n31114), .Y(n31104) );
  NOR2X1 U25547 ( .A(n31115), .B(n31116), .Y(n31114) );
  OAI22X1 U25548 ( .A(n26943), .B(n30254), .C(n26944), .D(n29989), .Y(n31116)
         );
  OAI22X1 U25549 ( .A(n26945), .B(n30015), .C(n25753), .D(n30007), .Y(n31115)
         );
  AOI22X1 U25550 ( .A(reg_A[57]), .B(n26007), .C(reg_A[59]), .D(n26008), .Y(
        n31113) );
  AOI22X1 U25551 ( .A(reg_A[58]), .B(n26009), .C(reg_A[62]), .D(n26010), .Y(
        n31112) );
  NOR2X1 U25552 ( .A(n31117), .B(n31118), .Y(n31102) );
  NAND2X1 U25553 ( .A(n31119), .B(n31120), .Y(n31118) );
  AOI22X1 U25554 ( .A(reg_A[63]), .B(n25613), .C(reg_A[60]), .D(n25749), .Y(
        n31120) );
  AOI22X1 U25555 ( .A(reg_A[61]), .B(n25750), .C(reg_A[56]), .D(n26924), .Y(
        n31119) );
  NAND2X1 U25556 ( .A(n31121), .B(n31122), .Y(n31117) );
  AOI22X1 U25557 ( .A(reg_A[57]), .B(n26803), .C(reg_A[59]), .D(n26804), .Y(
        n31122) );
  AOI22X1 U25558 ( .A(reg_A[58]), .B(n26927), .C(reg_A[62]), .D(n26878), .Y(
        n31121) );
  OAI21X1 U25559 ( .A(n26625), .B(n30463), .C(n31123), .Y(n31100) );
  AOI22X1 U25560 ( .A(reg_A[45]), .B(n26627), .C(reg_A[44]), .D(n26519), .Y(
        n31123) );
  NAND3X1 U25561 ( .A(n31124), .B(n31125), .C(n31126), .Y(result[55]) );
  NOR2X1 U25562 ( .A(n31127), .B(n31128), .Y(n31126) );
  NAND3X1 U25563 ( .A(n31129), .B(n31130), .C(n31131), .Y(n31128) );
  AOI22X1 U25564 ( .A(n26504), .B(n31132), .C(reg_A[51]), .D(n27132), .Y(
        n31131) );
  NAND2X1 U25565 ( .A(n31133), .B(n31134), .Y(n31132) );
  AOI22X1 U25566 ( .A(n31135), .B(n31136), .C(n31137), .D(n31138), .Y(n31134)
         );
  AOI22X1 U25567 ( .A(reg_B[55]), .B(n31139), .C(n31140), .D(reg_B[54]), .Y(
        n31133) );
  INVX1 U25568 ( .A(n31141), .Y(n31139) );
  OAI21X1 U25569 ( .A(n31142), .B(n31143), .C(n25999), .Y(n31130) );
  OAI22X1 U25570 ( .A(n25754), .B(n30174), .C(n31144), .D(n30299), .Y(n31143)
         );
  OAI22X1 U25571 ( .A(n30090), .B(n30378), .C(n27925), .D(n30168), .Y(n31142)
         );
  AOI22X1 U25572 ( .A(n30909), .B(n27110), .C(reg_A[50]), .D(n28050), .Y(
        n31129) );
  MUX2X1 U25573 ( .B(n30043), .A(n30168), .S(reg_B[4]), .Y(n30909) );
  NAND3X1 U25574 ( .A(n31145), .B(n31146), .C(n31147), .Y(n31127) );
  AOI21X1 U25575 ( .A(n31148), .B(n27067), .C(n31149), .Y(n31147) );
  OAI21X1 U25576 ( .A(n31150), .B(n31151), .C(n31152), .Y(n31149) );
  OAI21X1 U25577 ( .A(n31153), .B(n31154), .C(n25840), .Y(n31152) );
  NAND2X1 U25578 ( .A(n31155), .B(n31156), .Y(n31154) );
  NOR2X1 U25579 ( .A(n31157), .B(n31158), .Y(n31156) );
  OAI21X1 U25580 ( .A(n25043), .B(n30043), .C(n31159), .Y(n31158) );
  AOI22X1 U25581 ( .A(reg_A[54]), .B(n25135), .C(reg_A[53]), .D(n25252), .Y(
        n31159) );
  OAI21X1 U25582 ( .A(n25028), .B(n30008), .C(n31160), .Y(n31157) );
  AOI22X1 U25583 ( .A(reg_A[52]), .B(n25136), .C(reg_A[51]), .D(n25069), .Y(
        n31160) );
  NOR2X1 U25584 ( .A(n31161), .B(n31162), .Y(n31155) );
  OAI21X1 U25585 ( .A(n25034), .B(n30068), .C(n31163), .Y(n31162) );
  AOI22X1 U25586 ( .A(reg_A[49]), .B(n25253), .C(reg_A[48]), .D(n25628), .Y(
        n31163) );
  OAI21X1 U25587 ( .A(n25036), .B(n30066), .C(n31164), .Y(n31161) );
  AOI22X1 U25588 ( .A(reg_A[46]), .B(n25629), .C(reg_A[44]), .D(n25222), .Y(
        n31164) );
  NAND2X1 U25589 ( .A(n31165), .B(n31166), .Y(n31153) );
  NOR2X1 U25590 ( .A(n31167), .B(n31168), .Y(n31166) );
  OAI21X1 U25591 ( .A(n25039), .B(n30462), .C(n31169), .Y(n31168) );
  AOI22X1 U25592 ( .A(reg_A[41]), .B(n25234), .C(reg_A[43]), .D(n25635), .Y(
        n31169) );
  OAI21X1 U25593 ( .A(n25065), .B(n30744), .C(n31170), .Y(n31167) );
  AOI22X1 U25594 ( .A(reg_A[38]), .B(n25246), .C(reg_A[39]), .D(n25247), .Y(
        n31170) );
  NOR2X1 U25595 ( .A(n31171), .B(n31172), .Y(n31165) );
  OAI21X1 U25596 ( .A(n25238), .B(n30393), .C(n31173), .Y(n31172) );
  AOI22X1 U25597 ( .A(reg_A[36]), .B(n25487), .C(reg_A[37]), .D(n25241), .Y(
        n31173) );
  OAI21X1 U25598 ( .A(n26719), .B(n30394), .C(n31174), .Y(n31171) );
  AOI22X1 U25599 ( .A(reg_A[33]), .B(n25242), .C(reg_A[32]), .D(n25338), .Y(
        n31174) );
  NAND2X1 U25600 ( .A(n31137), .B(n25382), .Y(n31151) );
  NAND3X1 U25601 ( .A(n31175), .B(n31176), .C(n31177), .Y(n31148) );
  AOI21X1 U25602 ( .A(reg_A[55]), .B(n26924), .C(n31178), .Y(n31177) );
  OAI22X1 U25603 ( .A(n26800), .B(n30008), .C(n26801), .D(n30009), .Y(n31178)
         );
  AOI22X1 U25604 ( .A(reg_A[54]), .B(n26803), .C(reg_A[52]), .D(n26804), .Y(
        n31176) );
  AOI22X1 U25605 ( .A(reg_A[53]), .B(n26927), .C(reg_A[49]), .D(n26878), .Y(
        n31175) );
  OAI21X1 U25606 ( .A(n31179), .B(n31180), .C(n25188), .Y(n31146) );
  OAI21X1 U25607 ( .A(n31181), .B(n30210), .C(n30896), .Y(n31180) );
  AOI21X1 U25608 ( .A(reg_B[61]), .B(reg_A[48]), .C(n31182), .Y(n31181) );
  OAI21X1 U25609 ( .A(n31183), .B(n31184), .C(n25170), .Y(n31145) );
  OAI21X1 U25610 ( .A(n31185), .B(n30327), .C(n31186), .Y(n31184) );
  MUX2X1 U25611 ( .B(n31187), .A(n31188), .S(reg_B[55]), .Y(n31186) );
  NOR2X1 U25612 ( .A(n31189), .B(n26999), .Y(n31188) );
  OAI21X1 U25613 ( .A(n30299), .B(n31190), .C(n31191), .Y(n31187) );
  AOI22X1 U25614 ( .A(n31192), .B(n31193), .C(n31194), .D(reg_A[55]), .Y(
        n31191) );
  MUX2X1 U25615 ( .B(n30009), .A(n30174), .S(reg_B[54]), .Y(n31192) );
  INVX1 U25616 ( .A(n31075), .Y(n31185) );
  NAND2X1 U25617 ( .A(n31195), .B(n31196), .Y(n31075) );
  AOI22X1 U25618 ( .A(n30024), .B(n30343), .C(n30141), .D(n30694), .Y(n31196)
         );
  OAI21X1 U25619 ( .A(n30068), .B(n30109), .C(n31197), .Y(n30343) );
  AOI22X1 U25620 ( .A(n30112), .B(reg_A[39]), .C(reg_A[55]), .D(n30117), .Y(
        n31197) );
  AOI22X1 U25621 ( .A(n30201), .B(n30947), .C(n30342), .D(n31198), .Y(n31195)
         );
  OAI21X1 U25622 ( .A(n31199), .B(n30095), .C(n31200), .Y(n31183) );
  OAI21X1 U25623 ( .A(n31201), .B(n31179), .C(n25604), .Y(n31200) );
  OAI21X1 U25624 ( .A(n31052), .B(n30038), .C(n31202), .Y(n31179) );
  AOI22X1 U25625 ( .A(n30846), .B(n31056), .C(n30212), .D(n31053), .Y(n31202)
         );
  OAI21X1 U25626 ( .A(n30043), .B(n29975), .C(n30893), .Y(n31056) );
  NAND2X1 U25627 ( .A(n30326), .B(reg_A[51]), .Y(n30893) );
  NOR2X1 U25628 ( .A(n31203), .B(n30210), .Y(n31201) );
  INVX1 U25629 ( .A(n31204), .Y(n31199) );
  NOR2X1 U25630 ( .A(n31205), .B(n31206), .Y(n31125) );
  INVX1 U25631 ( .A(n31207), .Y(n31206) );
  AOI22X1 U25632 ( .A(n30120), .B(n31208), .C(n30236), .D(n31017), .Y(n31207)
         );
  NOR2X1 U25633 ( .A(n31209), .B(n31210), .Y(n31017) );
  OAI22X1 U25634 ( .A(n30223), .B(n30291), .C(n30256), .D(n31211), .Y(n31210)
         );
  NOR2X1 U25635 ( .A(n31212), .B(n31213), .Y(n30291) );
  OAI22X1 U25636 ( .A(reg_A[47]), .B(n30109), .C(reg_A[55]), .D(n29994), .Y(
        n31213) );
  OAI21X1 U25637 ( .A(reg_A[39]), .B(n31023), .C(n31024), .Y(n31212) );
  OAI22X1 U25638 ( .A(n30021), .B(n30960), .C(n30255), .D(n31214), .Y(n31209)
         );
  OAI21X1 U25639 ( .A(n25945), .B(n31215), .C(n31216), .Y(n31205) );
  AOI22X1 U25640 ( .A(reg_A[48]), .B(n27051), .C(reg_A[55]), .D(n27046), .Y(
        n31216) );
  AND2X1 U25641 ( .A(n31217), .B(n31218), .Y(n31124) );
  AOI21X1 U25642 ( .A(n25730), .B(n31219), .C(n31220), .Y(n31218) );
  OAI22X1 U25643 ( .A(n26012), .B(n31221), .C(n26525), .D(n31066), .Y(n31220)
         );
  NAND2X1 U25644 ( .A(n31222), .B(n31223), .Y(n31066) );
  AOI22X1 U25645 ( .A(n25025), .B(n31006), .C(n25026), .D(n30754), .Y(n31223)
         );
  INVX1 U25646 ( .A(n31224), .Y(n31006) );
  AOI22X1 U25647 ( .A(n26032), .B(n30753), .C(n26530), .D(n31225), .Y(n31222)
         );
  INVX1 U25648 ( .A(n30302), .Y(n30753) );
  NOR2X1 U25649 ( .A(n31226), .B(n31227), .Y(n30302) );
  OAI22X1 U25650 ( .A(reg_A[55]), .B(n26036), .C(reg_A[47]), .D(n26981), .Y(
        n31227) );
  OAI21X1 U25651 ( .A(reg_A[39]), .B(n26982), .C(n31072), .Y(n31226) );
  NAND3X1 U25652 ( .A(n31228), .B(n31229), .C(n31230), .Y(n31219) );
  NOR2X1 U25653 ( .A(n31231), .B(n31232), .Y(n31230) );
  OAI22X1 U25654 ( .A(n26936), .B(n30016), .C(n25745), .D(n29989), .Y(n31232)
         );
  OAI21X1 U25655 ( .A(n25062), .B(n29990), .C(n31233), .Y(n31231) );
  AOI22X1 U25656 ( .A(reg_A[56]), .B(n26803), .C(reg_A[58]), .D(n26804), .Y(
        n31233) );
  AOI22X1 U25657 ( .A(reg_A[59]), .B(n25749), .C(reg_A[60]), .D(n25750), .Y(
        n31229) );
  AOI22X1 U25658 ( .A(reg_A[63]), .B(n25615), .C(reg_A[55]), .D(n26924), .Y(
        n31228) );
  AOI22X1 U25659 ( .A(n25310), .B(n31234), .C(n31235), .D(n31236), .Y(n31217)
         );
  NAND3X1 U25660 ( .A(n31237), .B(n31238), .C(n31239), .Y(n31234) );
  NOR2X1 U25661 ( .A(n31240), .B(n31241), .Y(n31239) );
  OAI22X1 U25662 ( .A(n25030), .B(n30016), .C(n25033), .D(n29989), .Y(n31241)
         );
  OAI21X1 U25663 ( .A(n25040), .B(n29990), .C(n31242), .Y(n31240) );
  AOI22X1 U25664 ( .A(reg_A[56]), .B(n25135), .C(reg_A[58]), .D(n25136), .Y(
        n31242) );
  AOI22X1 U25665 ( .A(reg_A[59]), .B(n25072), .C(reg_A[60]), .D(n25123), .Y(
        n31238) );
  AOI22X1 U25666 ( .A(reg_A[63]), .B(n25124), .C(reg_A[55]), .D(n25125), .Y(
        n31237) );
  NAND3X1 U25667 ( .A(n31243), .B(n31244), .C(n31245), .Y(result[54]) );
  NOR2X1 U25668 ( .A(n31246), .B(n31247), .Y(n31245) );
  NAND3X1 U25669 ( .A(n31248), .B(n31249), .C(n31250), .Y(n31247) );
  AOI21X1 U25670 ( .A(n30261), .B(n31251), .C(n31252), .Y(n31250) );
  OAI21X1 U25671 ( .A(n31189), .B(n31253), .C(n31254), .Y(n31252) );
  OAI21X1 U25672 ( .A(n31255), .B(n31256), .C(n25310), .Y(n31254) );
  OR2X1 U25673 ( .A(n31257), .B(n31258), .Y(n31256) );
  OAI22X1 U25674 ( .A(n25043), .B(n30168), .C(n25467), .D(n30016), .Y(n31258)
         );
  OAI21X1 U25675 ( .A(n25037), .B(n30007), .C(n31259), .Y(n31257) );
  AOI22X1 U25676 ( .A(reg_A[58]), .B(n25072), .C(reg_A[59]), .D(n25123), .Y(
        n31259) );
  OR2X1 U25677 ( .A(n31260), .B(n31261), .Y(n31255) );
  OAI22X1 U25678 ( .A(n25030), .B(n29989), .C(n25033), .D(n30015), .Y(n31261)
         );
  OAI21X1 U25679 ( .A(n25040), .B(n30254), .C(n31262), .Y(n31260) );
  AOI22X1 U25680 ( .A(reg_A[55]), .B(n25135), .C(reg_A[57]), .D(n25136), .Y(
        n31262) );
  AOI21X1 U25681 ( .A(reg_B[54]), .B(n31263), .C(n31264), .Y(n31189) );
  AOI22X1 U25682 ( .A(n31265), .B(n31235), .C(reg_A[55]), .D(n27402), .Y(
        n31248) );
  NAND3X1 U25683 ( .A(n31266), .B(n31267), .C(n31268), .Y(n31246) );
  AOI21X1 U25684 ( .A(n25730), .B(n31269), .C(n31270), .Y(n31268) );
  OAI21X1 U25685 ( .A(n26012), .B(n31271), .C(n31272), .Y(n31270) );
  OAI21X1 U25686 ( .A(n31273), .B(n31274), .C(n26045), .Y(n31272) );
  NAND2X1 U25687 ( .A(n31275), .B(n31276), .Y(n31274) );
  AOI22X1 U25688 ( .A(reg_A[51]), .B(n27241), .C(reg_A[50]), .D(n27242), .Y(
        n31276) );
  AOI22X1 U25689 ( .A(reg_A[52]), .B(n27243), .C(reg_A[54]), .D(n25434), .Y(
        n31275) );
  OR2X1 U25690 ( .A(n31277), .B(n31278), .Y(n31273) );
  OAI22X1 U25691 ( .A(n27218), .B(n30299), .C(n25207), .D(n30174), .Y(n31278)
         );
  OAI21X1 U25692 ( .A(n27219), .B(n29655), .C(n31279), .Y(n31277) );
  OAI21X1 U25693 ( .A(n31280), .B(n31281), .C(n25044), .Y(n31279) );
  NAND3X1 U25694 ( .A(n31282), .B(n31283), .C(n31284), .Y(n31281) );
  NOR2X1 U25695 ( .A(n31285), .B(n31286), .Y(n31284) );
  OAI21X1 U25696 ( .A(n25036), .B(n30067), .C(n31287), .Y(n31286) );
  AOI22X1 U25697 ( .A(reg_A[46]), .B(n25124), .C(reg_A[43]), .D(n25222), .Y(
        n31287) );
  OAI21X1 U25698 ( .A(n25037), .B(n30066), .C(n31288), .Y(n31285) );
  AOI22X1 U25699 ( .A(reg_A[50]), .B(n25072), .C(reg_A[49]), .D(n25123), .Y(
        n31288) );
  AOI21X1 U25700 ( .A(reg_A[42]), .B(n25635), .C(n31289), .Y(n31283) );
  OAI22X1 U25701 ( .A(n25065), .B(n30059), .C(n25035), .D(n30744), .Y(n31289)
         );
  AOI22X1 U25702 ( .A(reg_A[41]), .B(n25325), .C(reg_A[54]), .D(n25125), .Y(
        n31282) );
  NAND2X1 U25703 ( .A(n31290), .B(n31291), .Y(n31280) );
  NOR2X1 U25704 ( .A(n31292), .B(n31293), .Y(n31291) );
  OAI21X1 U25705 ( .A(n25238), .B(n30394), .C(n31294), .Y(n31293) );
  AOI22X1 U25706 ( .A(reg_A[36]), .B(n25241), .C(reg_A[32]), .D(n25242), .Y(
        n31294) );
  OAI21X1 U25707 ( .A(n25038), .B(n30393), .C(n31295), .Y(n31292) );
  AOI22X1 U25708 ( .A(reg_A[37]), .B(n25246), .C(reg_A[38]), .D(n25247), .Y(
        n31295) );
  NOR2X1 U25709 ( .A(n31296), .B(n31297), .Y(n31290) );
  OAI21X1 U25710 ( .A(n25030), .B(n30068), .C(n31298), .Y(n31297) );
  AOI22X1 U25711 ( .A(reg_A[52]), .B(n25252), .C(reg_A[48]), .D(n25253), .Y(
        n31298) );
  OAI21X1 U25712 ( .A(n25041), .B(n30009), .C(n31299), .Y(n31296) );
  AOI22X1 U25713 ( .A(reg_A[33]), .B(n25257), .C(reg_A[53]), .D(n25135), .Y(
        n31299) );
  NAND3X1 U25714 ( .A(n31300), .B(n31301), .C(n31302), .Y(n31269) );
  NOR2X1 U25715 ( .A(n31303), .B(n31304), .Y(n31302) );
  OAI22X1 U25716 ( .A(n26936), .B(n29989), .C(n25745), .D(n30015), .Y(n31304)
         );
  OAI21X1 U25717 ( .A(n25062), .B(n30254), .C(n31305), .Y(n31303) );
  AOI22X1 U25718 ( .A(reg_A[55]), .B(n26803), .C(reg_A[57]), .D(n26804), .Y(
        n31305) );
  AOI21X1 U25719 ( .A(reg_A[63]), .B(n25614), .C(n31306), .Y(n31301) );
  OAI22X1 U25720 ( .A(n26800), .B(n29984), .C(n26801), .D(n30219), .Y(n31306)
         );
  AOI22X1 U25721 ( .A(reg_A[62]), .B(n25615), .C(reg_A[54]), .D(n26924), .Y(
        n31300) );
  AOI22X1 U25722 ( .A(reg_A[50]), .B(n31307), .C(n31076), .D(n31204), .Y(
        n31267) );
  NAND2X1 U25723 ( .A(n31308), .B(n31309), .Y(n31204) );
  AOI22X1 U25724 ( .A(n30024), .B(n30499), .C(n30141), .D(n30841), .Y(n31309)
         );
  OAI21X1 U25725 ( .A(n30069), .B(n30109), .C(n31310), .Y(n30499) );
  AOI22X1 U25726 ( .A(n30112), .B(reg_A[38]), .C(reg_A[54]), .D(n30117), .Y(
        n31310) );
  AOI22X1 U25727 ( .A(n30201), .B(n31081), .C(n30342), .D(n31311), .Y(n31308)
         );
  AOI22X1 U25728 ( .A(reg_A[49]), .B(n27256), .C(n31312), .D(n26028), .Y(
        n31266) );
  INVX1 U25729 ( .A(n31221), .Y(n31312) );
  NAND2X1 U25730 ( .A(n31313), .B(n31314), .Y(n31221) );
  AOI22X1 U25731 ( .A(n25025), .B(n31069), .C(n25026), .D(n30780), .Y(n31314)
         );
  INVX1 U25732 ( .A(n31315), .Y(n31069) );
  AOI22X1 U25733 ( .A(n26032), .B(n30779), .C(n26530), .D(n31316), .Y(n31313)
         );
  INVX1 U25734 ( .A(n30530), .Y(n30779) );
  NOR2X1 U25735 ( .A(n31317), .B(n31318), .Y(n30530) );
  OAI22X1 U25736 ( .A(reg_A[54]), .B(n26036), .C(reg_A[46]), .D(n26981), .Y(
        n31318) );
  OAI21X1 U25737 ( .A(reg_A[38]), .B(n26982), .C(n31072), .Y(n31317) );
  NOR2X1 U25738 ( .A(n31319), .B(n31320), .Y(n31244) );
  OAI21X1 U25739 ( .A(n31321), .B(n31322), .C(n31323), .Y(n31320) );
  AOI22X1 U25740 ( .A(reg_A[48]), .B(n31324), .C(reg_A[51]), .D(n27204), .Y(
        n31323) );
  OAI21X1 U25741 ( .A(n25032), .B(n30255), .C(n31325), .Y(n31324) );
  OR2X1 U25742 ( .A(n31326), .B(n31327), .Y(n31319) );
  OAI21X1 U25743 ( .A(n31328), .B(n30038), .C(n31329), .Y(n31327) );
  OAI21X1 U25744 ( .A(n31330), .B(n31331), .C(n31332), .Y(n31329) );
  INVX1 U25745 ( .A(n31333), .Y(n31331) );
  INVX1 U25746 ( .A(n31334), .Y(n31330) );
  AOI22X1 U25747 ( .A(n26267), .B(n31335), .C(n31182), .D(n25188), .Y(n31328)
         );
  INVX1 U25748 ( .A(n31203), .Y(n31335) );
  OAI21X1 U25749 ( .A(n27354), .B(n31336), .C(n31337), .Y(n31326) );
  NAND3X1 U25750 ( .A(n31264), .B(n31338), .C(n26504), .Y(n31337) );
  OAI21X1 U25751 ( .A(n30378), .B(n31339), .C(n31141), .Y(n31264) );
  AOI22X1 U25752 ( .A(reg_A[54]), .B(n31138), .C(reg_A[50]), .D(n31136), .Y(
        n31141) );
  AOI22X1 U25753 ( .A(n30846), .B(n31053), .C(reg_B[63]), .D(n31340), .Y(
        n31336) );
  OAI22X1 U25754 ( .A(n30168), .B(n29975), .C(n30008), .D(n30220), .Y(n31053)
         );
  NOR2X1 U25755 ( .A(n31341), .B(n31342), .Y(n31243) );
  OAI21X1 U25756 ( .A(n30233), .B(n31343), .C(n31344), .Y(n31342) );
  AOI22X1 U25757 ( .A(reg_A[54]), .B(n27184), .C(n31208), .D(n30236), .Y(
        n31344) );
  AND2X1 U25758 ( .A(n31345), .B(n31346), .Y(n31208) );
  AOI22X1 U25759 ( .A(n30024), .B(n30775), .C(n30141), .D(n30776), .Y(n31346)
         );
  INVX1 U25760 ( .A(n30509), .Y(n30775) );
  NOR2X1 U25761 ( .A(n31347), .B(n31348), .Y(n30509) );
  OAI22X1 U25762 ( .A(reg_A[46]), .B(n30109), .C(reg_A[54]), .D(n29994), .Y(
        n31348) );
  OAI21X1 U25763 ( .A(reg_A[38]), .B(n31023), .C(n31024), .Y(n31347) );
  AOI22X1 U25764 ( .A(n30342), .B(n31349), .C(n30201), .D(n31025), .Y(n31345)
         );
  INVX1 U25765 ( .A(n31350), .Y(n31025) );
  OAI21X1 U25766 ( .A(n31351), .B(n30378), .C(n31352), .Y(n31341) );
  AOI22X1 U25767 ( .A(n30132), .B(n29209), .C(reg_A[53]), .D(n27188), .Y(
        n31352) );
  INVX1 U25768 ( .A(n30765), .Y(n30132) );
  NAND2X1 U25769 ( .A(n31353), .B(n31354), .Y(n30765) );
  AOI22X1 U25770 ( .A(n26601), .B(n30378), .C(n26602), .D(n30009), .Y(n31354)
         );
  AOI22X1 U25771 ( .A(n27012), .B(n30168), .C(n26597), .D(n30299), .Y(n31353)
         );
  OR2X1 U25772 ( .A(n31355), .B(n31356), .Y(result[53]) );
  NAND3X1 U25773 ( .A(n31357), .B(n31358), .C(n31359), .Y(n31356) );
  NOR2X1 U25774 ( .A(n31360), .B(n31361), .Y(n31359) );
  OAI21X1 U25775 ( .A(n31362), .B(n31363), .C(n31364), .Y(n31361) );
  AOI22X1 U25776 ( .A(n31076), .B(n31251), .C(n31365), .D(n31332), .Y(n31364)
         );
  OAI21X1 U25777 ( .A(n30299), .B(n31366), .C(n31367), .Y(n31332) );
  AOI22X1 U25778 ( .A(n31136), .B(reg_A[49]), .C(n31368), .D(reg_A[51]), .Y(
        n31367) );
  NOR2X1 U25779 ( .A(n31369), .B(reg_B[54]), .Y(n31136) );
  NAND2X1 U25780 ( .A(n31370), .B(n31371), .Y(n31251) );
  AOI22X1 U25781 ( .A(n30024), .B(n30694), .C(n30141), .D(n30947), .Y(n31371)
         );
  OAI21X1 U25782 ( .A(n30066), .B(n30109), .C(n31372), .Y(n30694) );
  AOI22X1 U25783 ( .A(n30112), .B(reg_A[37]), .C(reg_A[53]), .D(n30117), .Y(
        n31372) );
  AOI22X1 U25784 ( .A(n30201), .B(n31198), .C(n30342), .D(n31373), .Y(n31370)
         );
  OAI21X1 U25785 ( .A(n31374), .B(n27152), .C(n31375), .Y(n31360) );
  AOI22X1 U25786 ( .A(reg_A[52]), .B(n27513), .C(n27358), .D(n31376), .Y(
        n31375) );
  NAND3X1 U25787 ( .A(n31377), .B(n31378), .C(n31379), .Y(n31376) );
  NOR2X1 U25788 ( .A(n31380), .B(n31381), .Y(n31379) );
  OAI22X1 U25789 ( .A(n27374), .B(n31215), .C(n27375), .D(n29655), .Y(n31381)
         );
  NAND2X1 U25790 ( .A(n31382), .B(n30403), .Y(n31215) );
  AOI22X1 U25791 ( .A(n30378), .B(n26295), .C(n30299), .D(n26293), .Y(n30403)
         );
  AOI22X1 U25792 ( .A(n26292), .B(n30174), .C(n26294), .D(n29655), .Y(n31382)
         );
  OAI22X1 U25793 ( .A(n27377), .B(n31271), .C(n27379), .D(n31383), .Y(n31380)
         );
  OAI21X1 U25794 ( .A(n31384), .B(n26030), .C(n31385), .Y(n31271) );
  AOI22X1 U25795 ( .A(n25025), .B(n31225), .C(n26032), .D(n30754), .Y(n31385)
         );
  OR2X1 U25796 ( .A(n31386), .B(n31387), .Y(n30754) );
  OAI22X1 U25797 ( .A(reg_A[53]), .B(n26036), .C(reg_A[45]), .D(n26981), .Y(
        n31387) );
  OAI21X1 U25798 ( .A(reg_A[37]), .B(n26982), .C(n31072), .Y(n31386) );
  INVX1 U25799 ( .A(n31388), .Y(n31225) );
  INVX1 U25800 ( .A(n31389), .Y(n31384) );
  AOI22X1 U25801 ( .A(reg_A[50]), .B(n27386), .C(reg_A[49]), .D(n27387), .Y(
        n31378) );
  AOI22X1 U25802 ( .A(reg_A[51]), .B(n27388), .C(reg_A[53]), .D(n27389), .Y(
        n31377) );
  AND2X1 U25803 ( .A(n31390), .B(n31391), .Y(n31374) );
  NOR2X1 U25804 ( .A(n31392), .B(n31393), .Y(n31391) );
  OAI21X1 U25805 ( .A(n26801), .B(n29990), .C(n31394), .Y(n31393) );
  AOI22X1 U25806 ( .A(reg_A[59]), .B(n26878), .C(reg_A[60]), .D(n25613), .Y(
        n31394) );
  OAI21X1 U25807 ( .A(n25062), .B(n30043), .C(n31395), .Y(n31392) );
  AOI22X1 U25808 ( .A(reg_A[54]), .B(n26803), .C(reg_A[56]), .D(n26804), .Y(
        n31395) );
  NOR2X1 U25809 ( .A(n31396), .B(n31397), .Y(n31390) );
  OAI22X1 U25810 ( .A(n25736), .B(n30299), .C(n31398), .D(n30007), .Y(n31397)
         );
  OAI21X1 U25811 ( .A(n27252), .B(n29989), .C(n31399), .Y(n31396) );
  AOI22X1 U25812 ( .A(reg_A[58]), .B(n25750), .C(reg_A[62]), .D(n25614), .Y(
        n31399) );
  AOI21X1 U25813 ( .A(reg_A[54]), .B(n27402), .C(n31400), .Y(n31358) );
  OAI22X1 U25814 ( .A(n31401), .B(n31402), .C(n31403), .D(n31333), .Y(n31400)
         );
  NOR2X1 U25815 ( .A(n31404), .B(n31405), .Y(n31357) );
  OAI21X1 U25816 ( .A(n25717), .B(n30043), .C(n31249), .Y(n31405) );
  INVX1 U25817 ( .A(n31406), .Y(n31249) );
  OAI21X1 U25818 ( .A(n25032), .B(n30896), .C(n31407), .Y(n31406) );
  NAND3X1 U25819 ( .A(reg_B[54]), .B(n26504), .C(n31263), .Y(n31407) );
  NAND2X1 U25820 ( .A(reg_B[60]), .B(reg_A[48]), .Y(n30896) );
  MUX2X1 U25821 ( .B(n31408), .A(n31409), .S(reg_B[63]), .Y(n31404) );
  NAND2X1 U25822 ( .A(n26267), .B(n31410), .Y(n31409) );
  NAND2X1 U25823 ( .A(n31340), .B(n27155), .Y(n31408) );
  OAI22X1 U25824 ( .A(reg_B[62]), .B(n31052), .C(n30009), .D(n31411), .Y(
        n31340) );
  AOI22X1 U25825 ( .A(reg_A[53]), .B(n30325), .C(reg_A[49]), .D(n30326), .Y(
        n31052) );
  NAND3X1 U25826 ( .A(n31412), .B(n31413), .C(n31414), .Y(n31355) );
  NOR2X1 U25827 ( .A(n31415), .B(n31416), .Y(n31414) );
  OAI21X1 U25828 ( .A(n27418), .B(n30009), .C(n31417), .Y(n31416) );
  AOI22X1 U25829 ( .A(reg_A[53]), .B(n27303), .C(reg_A[50]), .D(n27396), .Y(
        n31417) );
  OAI21X1 U25830 ( .A(n30233), .B(n31418), .C(n31419), .Y(n31415) );
  AOI22X1 U25831 ( .A(reg_A[48]), .B(n27316), .C(n31420), .D(n30236), .Y(
        n31419) );
  INVX1 U25832 ( .A(n31343), .Y(n31420) );
  OAI21X1 U25833 ( .A(n31214), .B(n30021), .C(n31421), .Y(n31343) );
  AOI22X1 U25834 ( .A(n30024), .B(n30704), .C(reg_B[62]), .D(n31422), .Y(
        n31421) );
  INVX1 U25835 ( .A(n31211), .Y(n30704) );
  NOR2X1 U25836 ( .A(n31423), .B(n31424), .Y(n31211) );
  OAI22X1 U25837 ( .A(reg_A[45]), .B(n30109), .C(reg_A[53]), .D(n29994), .Y(
        n31424) );
  OAI21X1 U25838 ( .A(reg_A[37]), .B(n31023), .C(n31024), .Y(n31423) );
  AOI21X1 U25839 ( .A(n31425), .B(n31426), .C(n31427), .Y(n31413) );
  OAI21X1 U25840 ( .A(n31428), .B(n25342), .C(n31429), .Y(n31427) );
  OAI21X1 U25841 ( .A(n31430), .B(n31431), .C(n25840), .Y(n31429) );
  NAND3X1 U25842 ( .A(n31432), .B(n31433), .C(n31434), .Y(n31431) );
  NOR2X1 U25843 ( .A(n31435), .B(n31436), .Y(n31434) );
  OAI21X1 U25844 ( .A(n25036), .B(n30160), .C(n31437), .Y(n31436) );
  AOI22X1 U25845 ( .A(reg_A[45]), .B(n25124), .C(reg_A[42]), .D(n25222), .Y(
        n31437) );
  OAI21X1 U25846 ( .A(n25037), .B(n30067), .C(n31438), .Y(n31435) );
  AOI22X1 U25847 ( .A(reg_A[49]), .B(n25072), .C(reg_A[48]), .D(n25123), .Y(
        n31438) );
  AOI21X1 U25848 ( .A(reg_A[41]), .B(n25635), .C(n31439), .Y(n31433) );
  OAI22X1 U25849 ( .A(n25065), .B(n30060), .C(n25475), .D(n30059), .Y(n31439)
         );
  AOI22X1 U25850 ( .A(reg_A[40]), .B(n25325), .C(reg_A[53]), .D(n25125), .Y(
        n31432) );
  NAND3X1 U25851 ( .A(n31440), .B(n31441), .C(n31442), .Y(n31430) );
  NOR2X1 U25852 ( .A(n31443), .B(n31444), .Y(n31442) );
  OAI21X1 U25853 ( .A(n26719), .B(n30395), .C(n31445), .Y(n31444) );
  AOI22X1 U25854 ( .A(reg_A[35]), .B(n25241), .C(reg_A[33]), .D(n25339), .Y(
        n31445) );
  OAI21X1 U25855 ( .A(n25038), .B(n30394), .C(n31446), .Y(n31443) );
  AOI22X1 U25856 ( .A(reg_A[36]), .B(n25246), .C(reg_A[37]), .D(n25247), .Y(
        n31446) );
  AOI21X1 U25857 ( .A(reg_A[51]), .B(n25252), .C(n31447), .Y(n31441) );
  OAI22X1 U25858 ( .A(n25041), .B(n30008), .C(n25042), .D(n30378), .Y(n31447)
         );
  AOI22X1 U25859 ( .A(reg_A[47]), .B(n25253), .C(reg_A[46]), .D(n25628), .Y(
        n31440) );
  AOI22X1 U25860 ( .A(n31368), .B(n31448), .C(n31140), .D(n31449), .Y(n31428)
         );
  MUX2X1 U25861 ( .B(n31450), .A(n31451), .S(reg_B[55]), .Y(n31140) );
  MUX2X1 U25862 ( .B(reg_A[52]), .A(reg_A[48]), .S(reg_B[53]), .Y(n31451) );
  MUX2X1 U25863 ( .B(reg_A[53]), .A(reg_A[49]), .S(reg_B[53]), .Y(n31450) );
  OAI21X1 U25864 ( .A(n30008), .B(n31338), .C(n31452), .Y(n31448) );
  INVX1 U25865 ( .A(n31453), .Y(n31426) );
  AOI21X1 U25866 ( .A(n25310), .B(n31454), .C(n31455), .Y(n31412) );
  OAI21X1 U25867 ( .A(n27431), .B(n30174), .C(n31456), .Y(n31455) );
  OAI21X1 U25868 ( .A(n31457), .B(n31458), .C(n25188), .Y(n31456) );
  OAI21X1 U25869 ( .A(n29655), .B(n31459), .C(n31460), .Y(n31458) );
  NAND3X1 U25870 ( .A(n30325), .B(reg_A[50]), .C(n30847), .Y(n31460) );
  NOR2X1 U25871 ( .A(n30378), .B(n30138), .Y(n31457) );
  NAND3X1 U25872 ( .A(n31461), .B(n31462), .C(n31463), .Y(n31454) );
  NOR2X1 U25873 ( .A(n31464), .B(n31465), .Y(n31463) );
  OAI22X1 U25874 ( .A(n25036), .B(n30007), .C(n25467), .D(n29989), .Y(n31465)
         );
  OAI21X1 U25875 ( .A(n25037), .B(n30016), .C(n31466), .Y(n31464) );
  AOI22X1 U25876 ( .A(reg_A[57]), .B(n25072), .C(reg_A[58]), .D(n25123), .Y(
        n31466) );
  AOI21X1 U25877 ( .A(reg_A[55]), .B(n25252), .C(n31467), .Y(n31462) );
  OAI22X1 U25878 ( .A(n25041), .B(n30254), .C(n25042), .D(n30168), .Y(n31467)
         );
  AOI22X1 U25879 ( .A(reg_A[59]), .B(n25253), .C(reg_A[60]), .D(n25628), .Y(
        n31461) );
  NAND3X1 U25880 ( .A(n31468), .B(n31469), .C(n31470), .Y(result[52]) );
  NOR2X1 U25881 ( .A(n31471), .B(n31472), .Y(n31470) );
  NAND3X1 U25882 ( .A(n31473), .B(n31474), .C(n31475), .Y(n31472) );
  NOR2X1 U25883 ( .A(n31476), .B(n31477), .Y(n31475) );
  OAI22X1 U25884 ( .A(n31401), .B(n31478), .C(n31403), .D(n31253), .Y(n31477)
         );
  INVX1 U25885 ( .A(n31479), .Y(n31403) );
  OAI21X1 U25886 ( .A(n30378), .B(n31366), .C(n31480), .Y(n31479) );
  AOI22X1 U25887 ( .A(n31368), .B(reg_A[50]), .C(n31263), .D(n31449), .Y(
        n31480) );
  INVX1 U25888 ( .A(n31235), .Y(n31401) );
  OAI21X1 U25889 ( .A(reg_B[59]), .B(n26996), .C(n27500), .Y(n31235) );
  OAI21X1 U25890 ( .A(n31362), .B(n30198), .C(n31481), .Y(n31476) );
  OAI21X1 U25891 ( .A(n31482), .B(n31483), .C(n27358), .Y(n31481) );
  OAI21X1 U25892 ( .A(n27442), .B(n30378), .C(n31484), .Y(n31483) );
  OAI21X1 U25893 ( .A(n31485), .B(n31486), .C(n25044), .Y(n31484) );
  OAI22X1 U25894 ( .A(n27454), .B(n31389), .C(n27455), .D(n31487), .Y(n31486)
         );
  NOR2X1 U25895 ( .A(reg_B[4]), .B(n31383), .Y(n31485) );
  OAI21X1 U25896 ( .A(n31488), .B(n26030), .C(n31489), .Y(n31383) );
  AOI22X1 U25897 ( .A(n25025), .B(n31316), .C(n26032), .D(n30780), .Y(n31489)
         );
  OR2X1 U25898 ( .A(n31490), .B(n31491), .Y(n30780) );
  OAI22X1 U25899 ( .A(reg_A[52]), .B(n26036), .C(reg_A[44]), .D(n26981), .Y(
        n31491) );
  OAI21X1 U25900 ( .A(reg_A[36]), .B(n26982), .C(n31072), .Y(n31490) );
  OAI22X1 U25901 ( .A(n27449), .B(n30518), .C(n27448), .D(n29655), .Y(n31482)
         );
  NAND2X1 U25902 ( .A(n31492), .B(n31493), .Y(n30518) );
  AOI22X1 U25903 ( .A(n26601), .B(n30008), .C(n26602), .D(n30174), .Y(n31493)
         );
  AOI22X1 U25904 ( .A(n27012), .B(n30378), .C(n26597), .D(n30009), .Y(n31492)
         );
  AND2X1 U25905 ( .A(n31494), .B(n31495), .Y(n31362) );
  AOI22X1 U25906 ( .A(n30024), .B(n30841), .C(n30141), .D(n31081), .Y(n31495)
         );
  OAI21X1 U25907 ( .A(n30067), .B(n30109), .C(n31496), .Y(n30841) );
  AOI22X1 U25908 ( .A(n30112), .B(reg_A[36]), .C(reg_A[52]), .D(n30117), .Y(
        n31496) );
  AOI22X1 U25909 ( .A(n30201), .B(n31311), .C(n30342), .D(n31497), .Y(n31494)
         );
  MUX2X1 U25910 ( .B(n31498), .A(n31499), .S(reg_B[63]), .Y(n31474) );
  AND2X1 U25911 ( .A(n27155), .B(n31500), .Y(n31499) );
  AND2X1 U25912 ( .A(n31410), .B(n26267), .Y(n31498) );
  OAI22X1 U25913 ( .A(reg_B[62]), .B(n31203), .C(n30008), .D(n31411), .Y(
        n31410) );
  AOI21X1 U25914 ( .A(reg_A[48]), .B(n30326), .C(n31182), .Y(n31203) );
  NOR2X1 U25915 ( .A(n29975), .B(n30378), .Y(n31182) );
  INVX1 U25916 ( .A(n31501), .Y(n31473) );
  OAI22X1 U25917 ( .A(n31363), .B(n31502), .C(n31333), .D(n31503), .Y(n31501)
         );
  NAND3X1 U25918 ( .A(n31504), .B(n31505), .C(n31506), .Y(n31471) );
  AOI21X1 U25919 ( .A(reg_A[53]), .B(n25282), .C(n31507), .Y(n31506) );
  OAI22X1 U25920 ( .A(n27971), .B(n29984), .C(n25295), .D(n30219), .Y(n31507)
         );
  AOI22X1 U25921 ( .A(reg_A[61]), .B(n25301), .C(reg_A[60]), .D(n25302), .Y(
        n31505) );
  AOI22X1 U25922 ( .A(reg_A[56]), .B(n29029), .C(reg_A[57]), .D(n29030), .Y(
        n31504) );
  NOR2X1 U25923 ( .A(n31508), .B(n31509), .Y(n31469) );
  OR2X1 U25924 ( .A(n31510), .B(n31511), .Y(n31509) );
  OAI22X1 U25925 ( .A(n31512), .B(n25342), .C(n31513), .D(n31514), .Y(n31511)
         );
  AOI21X1 U25926 ( .A(n31138), .B(n31515), .C(n31263), .Y(n31512) );
  NOR2X1 U25927 ( .A(n31369), .B(n29655), .Y(n31263) );
  OAI21X1 U25928 ( .A(reg_B[55]), .B(n30378), .C(n31516), .Y(n31515) );
  OAI21X1 U25929 ( .A(n31517), .B(n31321), .C(n31518), .Y(n31510) );
  OAI21X1 U25930 ( .A(n31519), .B(n31520), .C(reg_A[52]), .Y(n31518) );
  INVX1 U25931 ( .A(n31521), .Y(n31519) );
  INVX1 U25932 ( .A(n31425), .Y(n31321) );
  NOR2X1 U25933 ( .A(n25523), .B(reg_B[53]), .Y(n31425) );
  NAND3X1 U25934 ( .A(n31522), .B(n31523), .C(n31524), .Y(n31508) );
  AOI22X1 U25935 ( .A(reg_A[48]), .B(n31525), .C(reg_A[49]), .D(n31526), .Y(
        n31524) );
  OAI21X1 U25936 ( .A(n31190), .B(n31527), .C(n27419), .Y(n31526) );
  NAND2X1 U25937 ( .A(reg_B[55]), .B(n25372), .Y(n31527) );
  OAI21X1 U25938 ( .A(n30325), .B(n25794), .C(n31528), .Y(n31525) );
  INVX1 U25939 ( .A(n31529), .Y(n31528) );
  NAND3X1 U25940 ( .A(n30212), .B(n25932), .C(n31530), .Y(n31523) );
  INVX1 U25941 ( .A(n31422), .Y(n31530) );
  OAI21X1 U25942 ( .A(n31531), .B(n31532), .C(n25840), .Y(n31522) );
  NAND3X1 U25943 ( .A(n31533), .B(n31534), .C(n31535), .Y(n31532) );
  NOR2X1 U25944 ( .A(n31536), .B(n31537), .Y(n31535) );
  OAI22X1 U25945 ( .A(n25043), .B(n30378), .C(n25039), .D(n30059), .Y(n31537)
         );
  OAI21X1 U25946 ( .A(n25064), .B(n30744), .C(n31538), .Y(n31536) );
  AOI22X1 U25947 ( .A(reg_A[38]), .B(n25234), .C(reg_A[37]), .D(n25235), .Y(
        n31538) );
  AOI21X1 U25948 ( .A(reg_A[44]), .B(n25124), .C(n31539), .Y(n31534) );
  OAI22X1 U25949 ( .A(n25037), .B(n30160), .C(n25028), .D(n30068), .Y(n31539)
         );
  AOI22X1 U25950 ( .A(reg_A[41]), .B(n25222), .C(reg_A[42]), .D(n25637), .Y(
        n31533) );
  NAND3X1 U25951 ( .A(n31540), .B(n31541), .C(n31542), .Y(n31531) );
  NOR2X1 U25952 ( .A(n31543), .B(n31544), .Y(n31542) );
  OAI21X1 U25953 ( .A(n25042), .B(n30009), .C(n31545), .Y(n31544) );
  AOI22X1 U25954 ( .A(reg_A[34]), .B(n25241), .C(reg_A[32]), .D(n25339), .Y(
        n31545) );
  OAI21X1 U25955 ( .A(n25038), .B(n30170), .C(n31546), .Y(n31543) );
  AOI22X1 U25956 ( .A(reg_A[35]), .B(n25246), .C(reg_A[36]), .D(n25247), .Y(
        n31546) );
  AOI21X1 U25957 ( .A(reg_A[46]), .B(n25253), .C(n31547), .Y(n31541) );
  OAI22X1 U25958 ( .A(n25040), .B(n30008), .C(n25254), .D(n30174), .Y(n31547)
         );
  AOI22X1 U25959 ( .A(reg_A[45]), .B(n25628), .C(reg_A[48]), .D(n25069), .Y(
        n31540) );
  NOR2X1 U25960 ( .A(n31548), .B(n31549), .Y(n31468) );
  OAI21X1 U25961 ( .A(n31550), .B(n30007), .C(n31551), .Y(n31549) );
  AOI22X1 U25962 ( .A(reg_A[51]), .B(n27513), .C(reg_A[62]), .D(n25299), .Y(
        n31551) );
  INVX1 U25963 ( .A(n25300), .Y(n31550) );
  OR2X1 U25964 ( .A(n31552), .B(n31553), .Y(n31548) );
  OAI22X1 U25965 ( .A(n25360), .B(n30043), .C(n27420), .D(n30168), .Y(n31553)
         );
  OAI21X1 U25966 ( .A(n30290), .B(n31418), .C(n31554), .Y(n31552) );
  OAI21X1 U25967 ( .A(n27397), .B(n31555), .C(reg_A[50]), .Y(n31554) );
  OAI21X1 U25968 ( .A(n29975), .B(n31556), .C(n31557), .Y(n31555) );
  NAND3X1 U25969 ( .A(n25372), .B(n31338), .C(n31558), .Y(n31557) );
  INVX1 U25970 ( .A(n31190), .Y(n31558) );
  NAND2X1 U25971 ( .A(n29987), .B(n25188), .Y(n31556) );
  OAI21X1 U25972 ( .A(n31559), .B(n30293), .C(n31560), .Y(n31418) );
  AOI22X1 U25973 ( .A(n30024), .B(n30776), .C(n30201), .D(n31349), .Y(n31560)
         );
  OR2X1 U25974 ( .A(n31561), .B(n31562), .Y(n30776) );
  OAI22X1 U25975 ( .A(reg_A[44]), .B(n30109), .C(reg_A[52]), .D(n29994), .Y(
        n31562) );
  OAI21X1 U25976 ( .A(reg_A[36]), .B(n31023), .C(n31024), .Y(n31561) );
  INVX1 U25977 ( .A(n31563), .Y(n31559) );
  NAND3X1 U25978 ( .A(n31564), .B(n31565), .C(n31566), .Y(result[51]) );
  NOR2X1 U25979 ( .A(n31567), .B(n31568), .Y(n31566) );
  NAND3X1 U25980 ( .A(n31569), .B(n31570), .C(n31571), .Y(n31568) );
  NOR2X1 U25981 ( .A(n31572), .B(n31573), .Y(n31571) );
  OAI22X1 U25982 ( .A(n31574), .B(n31333), .C(n31502), .D(n30198), .Y(n31573)
         );
  AND2X1 U25983 ( .A(n31575), .B(n31576), .Y(n31502) );
  AOI22X1 U25984 ( .A(n30024), .B(n30947), .C(n30141), .D(n31198), .Y(n31576)
         );
  OAI21X1 U25985 ( .A(n30160), .B(n30109), .C(n31577), .Y(n30947) );
  AOI22X1 U25986 ( .A(n30112), .B(reg_A[35]), .C(reg_A[51]), .D(n30117), .Y(
        n31577) );
  AOI22X1 U25987 ( .A(n30201), .B(n31373), .C(n30342), .D(n31578), .Y(n31575)
         );
  MUX2X1 U25988 ( .B(n31579), .A(n31580), .S(reg_B[63]), .Y(n31572) );
  NAND2X1 U25989 ( .A(n26267), .B(n31581), .Y(n31580) );
  NAND2X1 U25990 ( .A(n31500), .B(n27155), .Y(n31579) );
  OAI22X1 U25991 ( .A(n30174), .B(n31411), .C(n30009), .D(n31582), .Y(n31500)
         );
  AOI22X1 U25992 ( .A(reg_A[58]), .B(n25293), .C(reg_A[52]), .D(n25282), .Y(
        n31570) );
  AOI22X1 U25993 ( .A(reg_A[51]), .B(n25283), .C(n31583), .D(n29565), .Y(
        n31569) );
  OAI21X1 U25994 ( .A(n25204), .B(n30009), .C(n31584), .Y(n31583) );
  AOI22X1 U25995 ( .A(reg_A[50]), .B(n25441), .C(reg_A[49]), .D(n27243), .Y(
        n31584) );
  NAND3X1 U25996 ( .A(n31585), .B(n31586), .C(n31587), .Y(n31567) );
  NOR2X1 U25997 ( .A(n31588), .B(n31589), .Y(n31587) );
  OAI22X1 U25998 ( .A(n25295), .B(n29990), .C(n25297), .D(n30254), .Y(n31589)
         );
  OAI22X1 U25999 ( .A(n27512), .B(n29984), .C(n31590), .D(n30015), .Y(n31588)
         );
  AOI22X1 U26000 ( .A(reg_A[53]), .B(n25364), .C(reg_A[54]), .D(n27622), .Y(
        n31586) );
  AOI22X1 U26001 ( .A(reg_A[61]), .B(n25299), .C(reg_A[62]), .D(n25300), .Y(
        n31585) );
  AND2X1 U26002 ( .A(n31591), .B(n31592), .Y(n31565) );
  NOR2X1 U26003 ( .A(n31593), .B(n31594), .Y(n31592) );
  OAI21X1 U26004 ( .A(n31503), .B(n31595), .C(n31596), .Y(n31594) );
  OAI21X1 U26005 ( .A(n31597), .B(n31598), .C(n25840), .Y(n31596) );
  NAND3X1 U26006 ( .A(n31599), .B(n31600), .C(n31601), .Y(n31598) );
  NOR2X1 U26007 ( .A(n31602), .B(n31603), .Y(n31601) );
  OAI22X1 U26008 ( .A(n25043), .B(n30009), .C(n25039), .D(n30060), .Y(n31603)
         );
  OAI21X1 U26009 ( .A(n25064), .B(n30059), .C(n31604), .Y(n31602) );
  AOI22X1 U26010 ( .A(reg_A[37]), .B(n25234), .C(reg_A[36]), .D(n25235), .Y(
        n31604) );
  AOI21X1 U26011 ( .A(reg_A[43]), .B(n25124), .C(n31605), .Y(n31600) );
  OAI22X1 U26012 ( .A(n25037), .B(n30462), .C(n25028), .D(n30069), .Y(n31605)
         );
  AOI22X1 U26013 ( .A(reg_A[40]), .B(n25222), .C(reg_A[41]), .D(n25637), .Y(
        n31599) );
  NAND3X1 U26014 ( .A(n31606), .B(n31607), .C(n31608), .Y(n31597) );
  NOR2X1 U26015 ( .A(n31609), .B(n31610), .Y(n31608) );
  OAI22X1 U26016 ( .A(n25042), .B(n30008), .C(n25331), .D(n30170), .Y(n31610)
         );
  OAI21X1 U26017 ( .A(n25038), .B(n30395), .C(n31611), .Y(n31609) );
  AOI22X1 U26018 ( .A(reg_A[34]), .B(n25246), .C(reg_A[35]), .D(n25247), .Y(
        n31611) );
  AOI21X1 U26019 ( .A(reg_A[45]), .B(n25253), .C(n31612), .Y(n31607) );
  OAI22X1 U26020 ( .A(n25040), .B(n30174), .C(n25041), .D(n29655), .Y(n31612)
         );
  AOI22X1 U26021 ( .A(reg_A[44]), .B(n25628), .C(reg_A[47]), .D(n25069), .Y(
        n31606) );
  AOI21X1 U26022 ( .A(n26504), .B(n31338), .C(n31365), .Y(n31595) );
  INVX1 U26023 ( .A(n31253), .Y(n31365) );
  AOI22X1 U26024 ( .A(reg_A[51]), .B(n31138), .C(reg_A[49]), .D(n31368), .Y(
        n31503) );
  OAI21X1 U26025 ( .A(n31613), .B(n31614), .C(n31615), .Y(n31593) );
  NAND3X1 U26026 ( .A(n27921), .B(n26602), .C(n31616), .Y(n31615) );
  NAND2X1 U26027 ( .A(n26597), .B(n27676), .Y(n31614) );
  NOR2X1 U26028 ( .A(n31617), .B(n31618), .Y(n31591) );
  OAI21X1 U26029 ( .A(n27825), .B(n31389), .C(n31619), .Y(n31618) );
  OAI21X1 U26030 ( .A(n31620), .B(n31621), .C(n25382), .Y(n31619) );
  OAI22X1 U26031 ( .A(n31622), .B(n31623), .C(n31624), .D(n31150), .Y(n31621)
         );
  INVX1 U26032 ( .A(n31625), .Y(n31622) );
  OAI21X1 U26033 ( .A(n31626), .B(n31190), .C(n31627), .Y(n31620) );
  NAND3X1 U26034 ( .A(n31137), .B(n31449), .C(n31193), .Y(n31627) );
  INVX1 U26035 ( .A(n31628), .Y(n31193) );
  OAI21X1 U26036 ( .A(reg_B[2]), .B(n31224), .C(n31629), .Y(n31389) );
  AOI21X1 U26037 ( .A(n27570), .B(n31630), .C(n31631), .Y(n31629) );
  NOR2X1 U26038 ( .A(n31632), .B(n31633), .Y(n31224) );
  OAI22X1 U26039 ( .A(reg_A[51]), .B(n26036), .C(reg_A[43]), .D(n26981), .Y(
        n31633) );
  OAI21X1 U26040 ( .A(reg_A[35]), .B(n26982), .C(n31072), .Y(n31632) );
  OAI21X1 U26041 ( .A(n25939), .B(n31487), .C(n31634), .Y(n31617) );
  NAND2X1 U26042 ( .A(reg_A[32]), .B(n31635), .Y(n31634) );
  OAI21X1 U26043 ( .A(n27455), .B(n31636), .C(n25583), .Y(n31635) );
  NOR2X1 U26044 ( .A(n31637), .B(n31638), .Y(n31564) );
  OAI21X1 U26045 ( .A(n27582), .B(n30007), .C(n31639), .Y(n31638) );
  AOI22X1 U26046 ( .A(reg_A[55]), .B(n25368), .C(n30261), .D(n31640), .Y(
        n31639) );
  NAND3X1 U26047 ( .A(n31641), .B(n31642), .C(n31643), .Y(n31637) );
  AOI22X1 U26048 ( .A(reg_A[50]), .B(n31644), .C(n31645), .D(n30847), .Y(
        n31643) );
  OAI21X1 U26049 ( .A(n31646), .B(n31647), .C(n25932), .Y(n31642) );
  OAI22X1 U26050 ( .A(n30038), .B(n31513), .C(n30320), .D(n31563), .Y(n31647)
         );
  OAI21X1 U26051 ( .A(n29970), .B(n31422), .C(n31648), .Y(n31646) );
  NAND3X1 U26052 ( .A(n30847), .B(n30341), .C(n31649), .Y(n31648) );
  OAI21X1 U26053 ( .A(reg_B[61]), .B(n30960), .C(n31650), .Y(n31422) );
  AOI21X1 U26054 ( .A(n31651), .B(n31652), .C(n31653), .Y(n31650) );
  INVX1 U26055 ( .A(n30040), .Y(n31652) );
  NOR2X1 U26056 ( .A(n31654), .B(n31655), .Y(n30960) );
  OAI22X1 U26057 ( .A(reg_A[43]), .B(n30109), .C(reg_A[51]), .D(n29994), .Y(
        n31655) );
  OAI21X1 U26058 ( .A(reg_A[35]), .B(n31023), .C(n31024), .Y(n31654) );
  OAI21X1 U26059 ( .A(n31656), .B(n31657), .C(reg_A[48]), .Y(n31641) );
  OAI22X1 U26060 ( .A(n27564), .B(n31658), .C(n25517), .D(n31628), .Y(n31657)
         );
  OAI21X1 U26061 ( .A(n31449), .B(n31334), .C(n31659), .Y(n31656) );
  AND2X1 U26062 ( .A(n31660), .B(n27587), .Y(n31659) );
  OAI21X1 U26063 ( .A(n30847), .B(n29975), .C(n25188), .Y(n31660) );
  NAND3X1 U26064 ( .A(n31661), .B(n31662), .C(n31663), .Y(result[50]) );
  NOR2X1 U26065 ( .A(n31664), .B(n31665), .Y(n31663) );
  NAND3X1 U26066 ( .A(n31666), .B(n31667), .C(n31668), .Y(n31665) );
  AOI21X1 U26067 ( .A(n30261), .B(n31669), .C(n31670), .Y(n31668) );
  OAI21X1 U26068 ( .A(n31671), .B(n31672), .C(n25203), .Y(n31667) );
  NAND3X1 U26069 ( .A(n31673), .B(n31674), .C(n31675), .Y(n31672) );
  AOI21X1 U26070 ( .A(reg_A[52]), .B(n27637), .C(n31676), .Y(n31675) );
  OAI22X1 U26071 ( .A(n25599), .B(n30299), .C(n25600), .D(n30043), .Y(n31676)
         );
  AOI22X1 U26072 ( .A(reg_A[50]), .B(n27639), .C(reg_A[51]), .D(n25617), .Y(
        n31674) );
  AOI22X1 U26073 ( .A(reg_A[54]), .B(n25650), .C(reg_A[56]), .D(n25651), .Y(
        n31673) );
  NAND3X1 U26074 ( .A(n31677), .B(n31678), .C(n31679), .Y(n31671) );
  AOI21X1 U26075 ( .A(reg_A[61]), .B(n27643), .C(n31680), .Y(n31679) );
  OAI22X1 U26076 ( .A(n27645), .B(n30015), .C(n27646), .D(n29984), .Y(n31680)
         );
  AOI22X1 U26077 ( .A(reg_A[62]), .B(n27647), .C(reg_A[63]), .D(n27648), .Y(
        n31678) );
  AOI22X1 U26078 ( .A(reg_A[57]), .B(n27649), .C(reg_A[58]), .D(n27650), .Y(
        n31677) );
  OAI21X1 U26079 ( .A(n31681), .B(n31682), .C(n25932), .Y(n31666) );
  OAI22X1 U26080 ( .A(n30320), .B(n31513), .C(n29970), .D(n31563), .Y(n31682)
         );
  OAI21X1 U26081 ( .A(reg_B[61]), .B(n31350), .C(n31683), .Y(n31563) );
  AOI21X1 U26082 ( .A(n31651), .B(n30243), .C(n31653), .Y(n31683) );
  NOR2X1 U26083 ( .A(n31684), .B(n31685), .Y(n31350) );
  OAI22X1 U26084 ( .A(reg_A[42]), .B(n30109), .C(reg_A[50]), .D(n29994), .Y(
        n31685) );
  OAI21X1 U26085 ( .A(reg_A[34]), .B(n31023), .C(n31024), .Y(n31684) );
  OAI21X1 U26086 ( .A(n30038), .B(n31686), .C(n31687), .Y(n31681) );
  OAI21X1 U26087 ( .A(n31688), .B(n31689), .C(n30847), .Y(n31687) );
  NOR2X1 U26088 ( .A(reg_B[59]), .B(n31690), .Y(n31688) );
  MUX2X1 U26089 ( .B(n31691), .A(n31692), .S(reg_B[61]), .Y(n31686) );
  OAI21X1 U26090 ( .A(reg_B[59]), .B(n30513), .C(n31693), .Y(n31692) );
  INVX1 U26091 ( .A(n31349), .Y(n31691) );
  OAI21X1 U26092 ( .A(reg_A[32]), .B(n30341), .C(n31694), .Y(n31349) );
  AOI22X1 U26093 ( .A(n30117), .B(n29655), .C(n30208), .D(n30744), .Y(n31694)
         );
  NAND2X1 U26094 ( .A(n31695), .B(n31696), .Y(n31664) );
  INVX1 U26095 ( .A(n31697), .Y(n31696) );
  OAI22X1 U26096 ( .A(n31698), .B(n31699), .C(n31574), .D(n31253), .Y(n31697)
         );
  AOI22X1 U26097 ( .A(reg_A[50]), .B(n31138), .C(reg_A[48]), .D(n31368), .Y(
        n31574) );
  NAND2X1 U26098 ( .A(n31700), .B(n27676), .Y(n31699) );
  AOI22X1 U26099 ( .A(n26597), .B(n31487), .C(n26009), .D(n31316), .Y(n31700)
         );
  OAI21X1 U26100 ( .A(reg_A[32]), .B(n27677), .C(n31701), .Y(n31316) );
  AOI22X1 U26101 ( .A(n26038), .B(n30744), .C(n26664), .D(n29655), .Y(n31701)
         );
  OAI21X1 U26102 ( .A(n31488), .B(n26599), .C(n31702), .Y(n31698) );
  AOI22X1 U26103 ( .A(n27680), .B(n30395), .C(n31703), .D(n27677), .Y(n31702)
         );
  OAI21X1 U26104 ( .A(n31704), .B(n25754), .C(n31705), .Y(n31703) );
  AOI22X1 U26105 ( .A(n26002), .B(n30756), .C(n26008), .D(n31630), .Y(n31705)
         );
  INVX1 U26106 ( .A(n31613), .Y(n31488) );
  OAI21X1 U26107 ( .A(reg_B[2]), .B(n31315), .C(n31706), .Y(n31613) );
  AOI21X1 U26108 ( .A(n27570), .B(n30232), .C(n31631), .Y(n31706) );
  NOR2X1 U26109 ( .A(n31707), .B(n31708), .Y(n31315) );
  OAI22X1 U26110 ( .A(reg_A[50]), .B(n25063), .C(reg_A[42]), .D(n26981), .Y(
        n31708) );
  OAI21X1 U26111 ( .A(reg_A[34]), .B(n26982), .C(n31072), .Y(n31707) );
  AOI22X1 U26112 ( .A(n31640), .B(n31076), .C(n25509), .D(reg_A[55]), .Y(
        n31695) );
  NAND2X1 U26113 ( .A(n31709), .B(n31710), .Y(n31640) );
  AOI22X1 U26114 ( .A(n30024), .B(n31081), .C(n30141), .D(n31311), .Y(n31710)
         );
  OAI21X1 U26115 ( .A(n30462), .B(n30109), .C(n31711), .Y(n31081) );
  AOI22X1 U26116 ( .A(n30112), .B(reg_A[34]), .C(reg_A[50]), .D(n30117), .Y(
        n31711) );
  AOI22X1 U26117 ( .A(n30201), .B(n31497), .C(n30342), .D(n31712), .Y(n31709)
         );
  NOR2X1 U26118 ( .A(n31713), .B(n31714), .Y(n31662) );
  OAI21X1 U26119 ( .A(n27698), .B(n29655), .C(n31715), .Y(n31714) );
  OAI21X1 U26120 ( .A(n31644), .B(n31716), .C(reg_A[49]), .Y(n31715) );
  NAND2X1 U26121 ( .A(n31717), .B(n31718), .Y(n31716) );
  OAI22X1 U26122 ( .A(n25794), .B(n30138), .C(n25517), .D(n31719), .Y(n31644)
         );
  NAND3X1 U26123 ( .A(n31720), .B(n31721), .C(n31722), .Y(n31713) );
  OAI21X1 U26124 ( .A(n31723), .B(n31724), .C(n25382), .Y(n31722) );
  OAI22X1 U26125 ( .A(n31623), .B(n31725), .C(n31628), .D(n31322), .Y(n31724)
         );
  NAND2X1 U26126 ( .A(n31726), .B(n31449), .Y(n31322) );
  INVX1 U26127 ( .A(n31727), .Y(n31725) );
  OAI22X1 U26128 ( .A(n31728), .B(n31190), .C(n31150), .D(n31516), .Y(n31723)
         );
  NAND3X1 U26129 ( .A(n31581), .B(n30028), .C(n26267), .Y(n31721) );
  OAI22X1 U26130 ( .A(n29655), .B(n31411), .C(n30008), .D(n31582), .Y(n31581)
         );
  NAND2X1 U26131 ( .A(n30325), .B(reg_B[62]), .Y(n31411) );
  OAI21X1 U26132 ( .A(n31729), .B(n31730), .C(n25840), .Y(n31720) );
  NAND3X1 U26133 ( .A(n31731), .B(n31732), .C(n31733), .Y(n31730) );
  NOR2X1 U26134 ( .A(n31734), .B(n31735), .Y(n31733) );
  OAI22X1 U26135 ( .A(n25035), .B(n30058), .C(n25219), .D(n30744), .Y(n31735)
         );
  OAI21X1 U26136 ( .A(n25027), .B(n30059), .C(n31736), .Y(n31734) );
  AOI22X1 U26137 ( .A(reg_A[41]), .B(n25629), .C(reg_A[42]), .D(n25124), .Y(
        n31736) );
  AOI22X1 U26138 ( .A(reg_A[35]), .B(n25235), .C(reg_A[38]), .D(n25635), .Y(
        n31732) );
  AOI22X1 U26139 ( .A(reg_A[37]), .B(n25325), .C(reg_A[50]), .D(n25125), .Y(
        n31731) );
  NAND3X1 U26140 ( .A(n31737), .B(n31738), .C(n31739), .Y(n31729) );
  NOR2X1 U26141 ( .A(n31740), .B(n31741), .Y(n31739) );
  OAI22X1 U26142 ( .A(n25041), .B(n30068), .C(n25042), .D(n30174), .Y(n31741)
         );
  OAI21X1 U26143 ( .A(n25051), .B(n30395), .C(n31742), .Y(n31740) );
  AOI22X1 U26144 ( .A(reg_A[33]), .B(n25246), .C(reg_A[34]), .D(n25247), .Y(
        n31742) );
  AOI21X1 U26145 ( .A(reg_A[43]), .B(n25628), .C(n31743), .Y(n31738) );
  OAI22X1 U26146 ( .A(n25033), .B(n30067), .C(n25133), .D(n29655), .Y(n31743)
         );
  AOI22X1 U26147 ( .A(reg_A[46]), .B(n25072), .C(reg_A[45]), .D(n25123), .Y(
        n31737) );
  NOR2X1 U26148 ( .A(n31744), .B(n31745), .Y(n31661) );
  OAI22X1 U26149 ( .A(n29782), .B(n30168), .C(n29765), .D(n30299), .Y(n31745)
         );
  OAI22X1 U26150 ( .A(n29766), .B(n30378), .C(n31746), .D(n30008), .Y(n31744)
         );
  INVX1 U26151 ( .A(n31747), .Y(n31746) );
  NAND3X1 U26152 ( .A(n31748), .B(n31749), .C(n31750), .Y(result[4]) );
  NOR2X1 U26153 ( .A(n31751), .B(n31752), .Y(n31750) );
  NAND3X1 U26154 ( .A(n31753), .B(n31754), .C(n31755), .Y(n31752) );
  AOI21X1 U26155 ( .A(reg_A[14]), .B(n25299), .C(n31756), .Y(n31755) );
  OAI22X1 U26156 ( .A(n25360), .B(n25132), .C(n27420), .D(n26677), .Y(n31756)
         );
  OAI21X1 U26157 ( .A(n31757), .B(n31758), .C(n25310), .Y(n31754) );
  NAND3X1 U26158 ( .A(n31759), .B(n31760), .C(n31761), .Y(n31758) );
  NOR2X1 U26159 ( .A(n31762), .B(n31763), .Y(n31761) );
  OAI22X1 U26160 ( .A(n29286), .B(n25316), .C(n27954), .D(n25318), .Y(n31763)
         );
  OAI22X1 U26161 ( .A(n25244), .B(n25320), .C(n25239), .D(n25322), .Y(n31762)
         );
  AOI22X1 U26162 ( .A(n25234), .B(reg_A[18]), .C(n25235), .D(reg_A[19]), .Y(
        n31760) );
  AOI22X1 U26163 ( .A(n25635), .B(reg_A[16]), .C(n25325), .D(reg_A[17]), .Y(
        n31759) );
  NAND3X1 U26164 ( .A(n31764), .B(n31765), .C(n31766), .Y(n31757) );
  NOR2X1 U26165 ( .A(n31767), .B(n31768), .Y(n31766) );
  OAI22X1 U26166 ( .A(n25331), .B(n25230), .C(n25038), .D(n26714), .Y(n31768)
         );
  OAI22X1 U26167 ( .A(n25334), .B(n30587), .C(n25336), .D(n25232), .Y(n31767)
         );
  AOI22X1 U26168 ( .A(n25242), .B(reg_A[26]), .C(n25338), .D(reg_A[27]), .Y(
        n31765) );
  AOI22X1 U26169 ( .A(reg_A[24]), .B(n25339), .C(n25257), .D(reg_A[25]), .Y(
        n31764) );
  AOI22X1 U26170 ( .A(reg_A[3]), .B(n31769), .C(reg_A[1]), .D(n31770), .Y(
        n31753) );
  NAND3X1 U26171 ( .A(n31771), .B(n31772), .C(n31773), .Y(n31751) );
  NOR2X1 U26172 ( .A(n31774), .B(n31775), .Y(n31773) );
  OAI21X1 U26173 ( .A(n31776), .B(n30569), .C(n31777), .Y(n31775) );
  OAI21X1 U26174 ( .A(n31778), .B(n31779), .C(n26480), .Y(n31777) );
  OAI22X1 U26175 ( .A(n26769), .B(n25106), .C(n31780), .D(n25099), .Y(n31779)
         );
  OAI22X1 U26176 ( .A(n26774), .B(n28033), .C(n31781), .D(n31782), .Y(n31778)
         );
  INVX1 U26177 ( .A(n31783), .Y(n26774) );
  NOR2X1 U26178 ( .A(n31784), .B(n31785), .Y(n31776) );
  OAI21X1 U26179 ( .A(n31786), .B(n31787), .C(n31788), .Y(n31785) );
  NAND2X1 U26180 ( .A(n26504), .B(n31789), .Y(n31787) );
  INVX1 U26181 ( .A(n31790), .Y(n31784) );
  OAI21X1 U26182 ( .A(n26741), .B(n27190), .C(n31791), .Y(n31774) );
  OAI21X1 U26183 ( .A(n31792), .B(n31793), .C(reg_A[2]), .Y(n31791) );
  OAI21X1 U26184 ( .A(n31794), .B(n31795), .C(reg_A[0]), .Y(n31772) );
  OAI21X1 U26185 ( .A(n31796), .B(n25794), .C(n31797), .Y(n31795) );
  OAI22X1 U26186 ( .A(n25110), .B(n27438), .C(n25342), .D(n31789), .Y(n31794)
         );
  AOI21X1 U26187 ( .A(n25372), .B(n31798), .C(n31799), .Y(n31771) );
  AOI21X1 U26188 ( .A(n31800), .B(n31801), .C(n25087), .Y(n31799) );
  AOI22X1 U26189 ( .A(n29245), .B(n26779), .C(n28038), .D(n31802), .Y(n31801)
         );
  AOI22X1 U26190 ( .A(n27984), .B(n31803), .C(n28023), .D(n31804), .Y(n31800)
         );
  OAI21X1 U26191 ( .A(n31805), .B(n31806), .C(n31807), .Y(n31798) );
  AOI22X1 U26192 ( .A(n31808), .B(n28023), .C(n31809), .D(reg_A[4]), .Y(n31807) );
  NOR2X1 U26193 ( .A(n25189), .B(n25128), .Y(n31808) );
  NOR2X1 U26194 ( .A(n31810), .B(n31811), .Y(n31749) );
  OAI21X1 U26195 ( .A(n27971), .B(n27967), .C(n31812), .Y(n31811) );
  AOI22X1 U26196 ( .A(reg_A[9]), .B(n29030), .C(reg_A[10]), .D(n29031), .Y(
        n31812) );
  NAND2X1 U26197 ( .A(n31813), .B(n31814), .Y(n31810) );
  AOI22X1 U26198 ( .A(reg_A[15]), .B(n25300), .C(reg_A[13]), .D(n25301), .Y(
        n31814) );
  AOI22X1 U26199 ( .A(reg_A[12]), .B(n25302), .C(reg_A[8]), .D(n29029), .Y(
        n31813) );
  NOR2X1 U26200 ( .A(n31815), .B(n31816), .Y(n31748) );
  OR2X1 U26201 ( .A(n31817), .B(n31818), .Y(n31816) );
  OAI21X1 U26202 ( .A(n31805), .B(n30547), .C(n31819), .Y(n31818) );
  MUX2X1 U26203 ( .B(n30550), .A(n31820), .S(reg_B[15]), .Y(n31819) );
  NOR2X1 U26204 ( .A(n31821), .B(n25023), .Y(n30550) );
  AOI22X1 U26205 ( .A(n29256), .B(n29257), .C(reg_A[2]), .D(n30551), .Y(n31821) );
  OAI22X1 U26206 ( .A(n30569), .B(n29304), .C(n26742), .D(n30552), .Y(n29257)
         );
  INVX1 U26207 ( .A(n31822), .Y(n31805) );
  MUX2X1 U26208 ( .B(n31823), .A(n31824), .S(reg_B[7]), .Y(n31817) );
  OR2X1 U26209 ( .A(n31825), .B(n28213), .Y(n31824) );
  INVX1 U26210 ( .A(n30603), .Y(n31823) );
  OAI21X1 U26211 ( .A(n30609), .B(n31826), .C(n31827), .Y(n30603) );
  NAND3X1 U26212 ( .A(n29323), .B(n28005), .C(n26186), .Y(n31827) );
  INVX1 U26213 ( .A(n30623), .Y(n29323) );
  MUX2X1 U26214 ( .B(reg_A[4]), .A(reg_A[0]), .S(reg_B[5]), .Y(n30623) );
  OAI21X1 U26215 ( .A(n26504), .B(n26186), .C(reg_A[2]), .Y(n31826) );
  OAI21X1 U26216 ( .A(n30546), .B(n31828), .C(n31829), .Y(n31815) );
  AOI22X1 U26217 ( .A(reg_A[5]), .B(n25282), .C(n31830), .D(n31831), .Y(n31829) );
  INVX1 U26218 ( .A(n31832), .Y(n30546) );
  OAI22X1 U26219 ( .A(reg_B[30]), .B(n27979), .C(n25128), .D(n31833), .Y(
        n31832) );
  AOI21X1 U26220 ( .A(reg_A[0]), .B(n25101), .C(n29317), .Y(n27979) );
  NAND3X1 U26221 ( .A(n31834), .B(n31835), .C(n31836), .Y(result[49]) );
  NOR2X1 U26222 ( .A(n31837), .B(n31838), .Y(n31836) );
  NAND3X1 U26223 ( .A(n31839), .B(n31840), .C(n31841), .Y(n31838) );
  AOI21X1 U26224 ( .A(n31076), .B(n31669), .C(n31842), .Y(n31841) );
  OAI22X1 U26225 ( .A(n31843), .B(n31363), .C(n25652), .D(n30168), .Y(n31842)
         );
  NAND2X1 U26226 ( .A(n31844), .B(n31845), .Y(n31669) );
  AOI22X1 U26227 ( .A(n30024), .B(n31198), .C(n30141), .D(n31373), .Y(n31845)
         );
  OAI21X1 U26228 ( .A(n30463), .B(n30109), .C(n31846), .Y(n31198) );
  AOI22X1 U26229 ( .A(n30112), .B(reg_A[33]), .C(reg_A[49]), .D(n30117), .Y(
        n31846) );
  AOI22X1 U26230 ( .A(n30201), .B(n31578), .C(n30342), .D(n31847), .Y(n31844)
         );
  OAI21X1 U26231 ( .A(n31848), .B(n31849), .C(n25203), .Y(n31840) );
  NAND3X1 U26232 ( .A(n31850), .B(n31851), .C(n31852), .Y(n31849) );
  AOI22X1 U26233 ( .A(reg_A[52]), .B(n27740), .C(reg_A[51]), .D(n27637), .Y(
        n31852) );
  OAI21X1 U26234 ( .A(n31853), .B(n31854), .C(n25044), .Y(n31851) );
  NAND2X1 U26235 ( .A(n31855), .B(n31856), .Y(n31854) );
  AOI22X1 U26236 ( .A(reg_A[59]), .B(n25637), .C(reg_A[63]), .D(n25234), .Y(
        n31856) );
  AOI22X1 U26237 ( .A(reg_A[61]), .B(n25635), .C(reg_A[62]), .D(n25325), .Y(
        n31855) );
  NAND2X1 U26238 ( .A(n31857), .B(n31858), .Y(n31853) );
  AOI22X1 U26239 ( .A(reg_A[56]), .B(n25628), .C(reg_A[58]), .D(n25629), .Y(
        n31858) );
  AOI22X1 U26240 ( .A(reg_A[57]), .B(n25124), .C(reg_A[60]), .D(n25222), .Y(
        n31857) );
  OAI21X1 U26241 ( .A(n31859), .B(n31860), .C(n25604), .Y(n31850) );
  NAND2X1 U26242 ( .A(n31861), .B(n31862), .Y(n31860) );
  AOI22X1 U26243 ( .A(reg_A[59]), .B(n25607), .C(reg_A[63]), .D(n25608), .Y(
        n31862) );
  AOI22X1 U26244 ( .A(reg_A[61]), .B(n25609), .C(reg_A[62]), .D(n25610), .Y(
        n31861) );
  NAND2X1 U26245 ( .A(n31863), .B(n31864), .Y(n31859) );
  AOI22X1 U26246 ( .A(reg_A[56]), .B(n25613), .C(reg_A[58]), .D(n25614), .Y(
        n31864) );
  AOI22X1 U26247 ( .A(reg_A[57]), .B(n25615), .C(reg_A[60]), .D(n25616), .Y(
        n31863) );
  OR2X1 U26248 ( .A(n31865), .B(n31866), .Y(n31848) );
  OAI22X1 U26249 ( .A(n25600), .B(n30168), .C(n27755), .D(n30043), .Y(n31866)
         );
  OAI21X1 U26250 ( .A(n27756), .B(n30299), .C(n31867), .Y(n31865) );
  AOI22X1 U26251 ( .A(reg_A[49]), .B(n27639), .C(reg_A[50]), .D(n25617), .Y(
        n31867) );
  INVX1 U26252 ( .A(n31670), .Y(n31839) );
  OAI22X1 U26253 ( .A(n25583), .B(n30395), .C(n29655), .D(n31868), .Y(n31670)
         );
  OAI21X1 U26254 ( .A(n31869), .B(n31870), .C(n25372), .Y(n31868) );
  OAI21X1 U26255 ( .A(n30222), .B(n25415), .C(n31628), .Y(n31870) );
  INVX1 U26256 ( .A(n31582), .Y(n30222) );
  NAND2X1 U26257 ( .A(n30024), .B(n30853), .Y(n31582) );
  NOR2X1 U26258 ( .A(n26999), .B(n31449), .Y(n31869) );
  NAND2X1 U26259 ( .A(n31871), .B(n31872), .Y(n31837) );
  AOI21X1 U26260 ( .A(reg_A[51]), .B(n25506), .C(n31873), .Y(n31872) );
  OAI21X1 U26261 ( .A(n31874), .B(n30395), .C(n31875), .Y(n31873) );
  OAI21X1 U26262 ( .A(n31876), .B(n31877), .C(reg_A[48]), .Y(n31875) );
  OAI21X1 U26263 ( .A(n25032), .B(n30028), .C(n31717), .Y(n31877) );
  INVX1 U26264 ( .A(n31878), .Y(n31717) );
  OAI21X1 U26265 ( .A(n31366), .B(n31333), .C(n31879), .Y(n31878) );
  AOI21X1 U26266 ( .A(n31880), .B(n26267), .C(n27770), .Y(n31879) );
  INVX1 U26267 ( .A(n30138), .Y(n31880) );
  NAND2X1 U26268 ( .A(n30492), .B(n30853), .Y(n30138) );
  NAND2X1 U26269 ( .A(reg_B[55]), .B(n26186), .Y(n31333) );
  NAND2X1 U26270 ( .A(n31334), .B(n27767), .Y(n31876) );
  NAND2X1 U26271 ( .A(reg_B[55]), .B(n26504), .Y(n31334) );
  INVX1 U26272 ( .A(n27778), .Y(n31874) );
  AOI22X1 U26273 ( .A(reg_A[52]), .B(n25507), .C(reg_A[53]), .D(n25508), .Y(
        n31871) );
  NOR2X1 U26274 ( .A(n31881), .B(n31882), .Y(n31835) );
  OAI21X1 U26275 ( .A(n27820), .B(n30756), .C(n31883), .Y(n31882) );
  OAI21X1 U26276 ( .A(n31884), .B(n31747), .C(reg_A[49]), .Y(n31883) );
  NAND3X1 U26277 ( .A(n31885), .B(n31521), .C(n31886), .Y(n31747) );
  INVX1 U26278 ( .A(n27687), .Y(n31886) );
  NAND3X1 U26279 ( .A(n25188), .B(n30853), .C(n30107), .Y(n31521) );
  NAND3X1 U26280 ( .A(n31887), .B(n31338), .C(n31194), .Y(n31885) );
  INVX1 U26281 ( .A(n31888), .Y(n30756) );
  NAND3X1 U26282 ( .A(n31889), .B(n31890), .C(n31891), .Y(n31881) );
  OAI21X1 U26283 ( .A(n31892), .B(n31893), .C(n25382), .Y(n31891) );
  OAI22X1 U26284 ( .A(n31623), .B(n31894), .C(n31453), .D(n31628), .Y(n31893)
         );
  MUX2X1 U26285 ( .B(n31895), .A(n31137), .S(reg_B[54]), .Y(n31453) );
  NOR2X1 U26286 ( .A(n30043), .B(reg_B[55]), .Y(n31137) );
  INVX1 U26287 ( .A(n31626), .Y(n31895) );
  MUX2X1 U26288 ( .B(reg_A[53]), .A(reg_A[54]), .S(reg_B[55]), .Y(n31626) );
  INVX1 U26289 ( .A(n31896), .Y(n31894) );
  OAI22X1 U26290 ( .A(n31624), .B(n31190), .C(n30008), .D(n31719), .Y(n31892)
         );
  AOI21X1 U26291 ( .A(reg_A[52]), .B(reg_B[55]), .C(n31135), .Y(n31624) );
  INVX1 U26292 ( .A(n31452), .Y(n31135) );
  NAND2X1 U26293 ( .A(reg_A[51]), .B(n31338), .Y(n31452) );
  NAND3X1 U26294 ( .A(n30120), .B(n30341), .C(n31897), .Y(n31890) );
  INVX1 U26295 ( .A(n31898), .Y(n31897) );
  OAI21X1 U26296 ( .A(n31899), .B(n31900), .C(n25840), .Y(n31889) );
  NAND3X1 U26297 ( .A(n31901), .B(n31902), .C(n31903), .Y(n31900) );
  NOR2X1 U26298 ( .A(n31904), .B(n31905), .Y(n31903) );
  OAI22X1 U26299 ( .A(n25035), .B(n30393), .C(n25219), .D(n30059), .Y(n31905)
         );
  OAI21X1 U26300 ( .A(n25027), .B(n30060), .C(n31906), .Y(n31904) );
  AOI22X1 U26301 ( .A(reg_A[40]), .B(n25629), .C(reg_A[41]), .D(n25124), .Y(
        n31906) );
  AOI22X1 U26302 ( .A(reg_A[34]), .B(n25235), .C(reg_A[37]), .D(n25635), .Y(
        n31902) );
  AOI22X1 U26303 ( .A(reg_A[36]), .B(n25325), .C(reg_A[49]), .D(n25125), .Y(
        n31901) );
  NAND3X1 U26304 ( .A(n31907), .B(n31908), .C(n31909), .Y(n31899) );
  NOR2X1 U26305 ( .A(n31910), .B(n31911), .Y(n31909) );
  OAI22X1 U26306 ( .A(n25040), .B(n30068), .C(n25041), .D(n30069), .Y(n31911)
         );
  OAI21X1 U26307 ( .A(n25042), .B(n29655), .C(n31912), .Y(n31910) );
  AOI22X1 U26308 ( .A(reg_A[32]), .B(n25246), .C(reg_A[33]), .D(n25247), .Y(
        n31912) );
  AOI22X1 U26309 ( .A(reg_A[43]), .B(n25253), .C(reg_A[42]), .D(n25628), .Y(
        n31908) );
  AOI22X1 U26310 ( .A(reg_A[45]), .B(n25072), .C(reg_A[44]), .D(n25123), .Y(
        n31907) );
  NOR2X1 U26311 ( .A(n31913), .B(n31914), .Y(n31834) );
  OAI21X1 U26312 ( .A(n25702), .B(n30043), .C(n31915), .Y(n31914) );
  OAI21X1 U26313 ( .A(n31916), .B(n31917), .C(n25932), .Y(n31915) );
  MUX2X1 U26314 ( .B(n31693), .A(n31513), .S(n30846), .Y(n31917) );
  OAI21X1 U26315 ( .A(reg_B[61]), .B(n31214), .C(n31918), .Y(n31513) );
  AOI21X1 U26316 ( .A(n31651), .B(n30296), .C(n31653), .Y(n31918) );
  INVX1 U26317 ( .A(n31919), .Y(n31653) );
  NAND3X1 U26318 ( .A(reg_B[61]), .B(n30395), .C(reg_B[59]), .Y(n31919) );
  NOR2X1 U26319 ( .A(n29973), .B(reg_B[59]), .Y(n31651) );
  NOR2X1 U26320 ( .A(n31920), .B(n31921), .Y(n31214) );
  OAI22X1 U26321 ( .A(reg_A[41]), .B(n30109), .C(reg_A[49]), .D(n29994), .Y(
        n31921) );
  OAI21X1 U26322 ( .A(reg_A[33]), .B(n31023), .C(n31024), .Y(n31920) );
  NAND2X1 U26323 ( .A(n30111), .B(n30395), .Y(n31024) );
  NOR2X1 U26324 ( .A(n30341), .B(n30853), .Y(n30111) );
  NOR2X1 U26325 ( .A(n30038), .B(n31922), .Y(n31916) );
  OR2X1 U26326 ( .A(n31690), .B(reg_B[59]), .Y(n31922) );
  MUX2X1 U26327 ( .B(n30040), .A(n31923), .S(reg_B[61]), .Y(n31690) );
  OAI21X1 U26328 ( .A(n27826), .B(n31630), .C(n31924), .Y(n31913) );
  INVX1 U26329 ( .A(n31925), .Y(n31924) );
  OAI22X1 U26330 ( .A(n31926), .B(n27821), .C(n31487), .D(n27825), .Y(n31925)
         );
  OAI21X1 U26331 ( .A(reg_B[2]), .B(n31388), .C(n31927), .Y(n31487) );
  AOI21X1 U26332 ( .A(n27570), .B(n30308), .C(n31631), .Y(n31927) );
  AND2X1 U26333 ( .A(n27828), .B(n30395), .Y(n31631) );
  NOR2X1 U26334 ( .A(n31928), .B(n31929), .Y(n31388) );
  OAI22X1 U26335 ( .A(reg_A[49]), .B(n26036), .C(reg_A[41]), .D(n25058), .Y(
        n31929) );
  OAI21X1 U26336 ( .A(reg_A[33]), .B(n25055), .C(n31072), .Y(n31928) );
  NAND2X1 U26337 ( .A(n26662), .B(n30395), .Y(n31072) );
  NAND3X1 U26338 ( .A(n31930), .B(n31931), .C(n31932), .Y(result[48]) );
  NOR2X1 U26339 ( .A(n31933), .B(n31934), .Y(n31932) );
  NAND2X1 U26340 ( .A(n31935), .B(n31936), .Y(n31934) );
  AOI21X1 U26341 ( .A(reg_A[41]), .B(n27860), .C(n31937), .Y(n31936) );
  OAI21X1 U26342 ( .A(n27839), .B(n31926), .C(n31938), .Y(n31937) );
  OAI21X1 U26343 ( .A(n27844), .B(n31884), .C(reg_A[48]), .Y(n31938) );
  OAI21X1 U26344 ( .A(n31366), .B(n31253), .C(n31939), .Y(n31884) );
  NAND3X1 U26345 ( .A(n26267), .B(n30853), .C(n30107), .Y(n31939) );
  NAND2X1 U26346 ( .A(n26186), .B(n31338), .Y(n31253) );
  OAI21X1 U26347 ( .A(reg_B[3]), .B(n31616), .C(n31940), .Y(n31926) );
  AOI22X1 U26348 ( .A(n26530), .B(n31941), .C(n25026), .D(n30232), .Y(n31940)
         );
  MUX2X1 U26349 ( .B(reg_A[38]), .A(reg_A[46]), .S(n26596), .Y(n30232) );
  INVX1 U26350 ( .A(n31942), .Y(n31941) );
  INVX1 U26351 ( .A(n31943), .Y(n31616) );
  OAI21X1 U26352 ( .A(reg_A[48]), .B(n27857), .C(n31944), .Y(n31943) );
  AOI22X1 U26353 ( .A(n27859), .B(n30744), .C(reg_B[2]), .D(n30536), .Y(n31944) );
  AOI22X1 U26354 ( .A(reg_A[33]), .B(n27861), .C(n27921), .D(n31945), .Y(
        n31935) );
  OAI21X1 U26355 ( .A(n27925), .B(n31630), .C(n31946), .Y(n31945) );
  AOI22X1 U26356 ( .A(n31947), .B(n26008), .C(n31888), .D(n25751), .Y(n31946)
         );
  INVX1 U26357 ( .A(n30046), .Y(n31630) );
  MUX2X1 U26358 ( .B(n30068), .A(n30059), .S(reg_B[1]), .Y(n30046) );
  NAND3X1 U26359 ( .A(n31948), .B(n31949), .C(n31950), .Y(n31933) );
  NOR2X1 U26360 ( .A(n31951), .B(n31952), .Y(n31950) );
  OAI21X1 U26361 ( .A(n30233), .B(n31953), .C(n31954), .Y(n31952) );
  NAND2X1 U26362 ( .A(n30342), .B(n31955), .Y(n31953) );
  INVX1 U26363 ( .A(n31956), .Y(n31951) );
  OAI21X1 U26364 ( .A(n31957), .B(n31958), .C(n25840), .Y(n31956) );
  NAND3X1 U26365 ( .A(n31959), .B(n31960), .C(n31961), .Y(n31958) );
  NOR2X1 U26366 ( .A(n31962), .B(n31963), .Y(n31961) );
  OAI22X1 U26367 ( .A(n25043), .B(n29655), .C(n25039), .D(n30393), .Y(n31963)
         );
  OAI22X1 U26368 ( .A(n25064), .B(n30058), .C(n25065), .D(n30170), .Y(n31962)
         );
  AOI22X1 U26369 ( .A(reg_A[40]), .B(n25124), .C(reg_A[37]), .D(n25222), .Y(
        n31960) );
  AOI22X1 U26370 ( .A(reg_A[38]), .B(n25637), .C(reg_A[34]), .D(n25234), .Y(
        n31959) );
  NAND3X1 U26371 ( .A(n31964), .B(n31965), .C(n31966), .Y(n31957) );
  NOR2X1 U26372 ( .A(n31967), .B(n31968), .Y(n31966) );
  OAI22X1 U26373 ( .A(n25033), .B(n30462), .C(n25040), .D(n30069), .Y(n31968)
         );
  OAI21X1 U26374 ( .A(n25041), .B(n30066), .C(n31969), .Y(n31967) );
  AOI22X1 U26375 ( .A(reg_A[32]), .B(n25247), .C(reg_A[47]), .D(n25135), .Y(
        n31969) );
  AOI22X1 U26376 ( .A(reg_A[41]), .B(n25628), .C(reg_A[44]), .D(n25069), .Y(
        n31965) );
  AOI22X1 U26377 ( .A(reg_A[43]), .B(n25123), .C(reg_A[39]), .D(n25629), .Y(
        n31964) );
  OAI21X1 U26378 ( .A(n31970), .B(n31971), .C(n25730), .Y(n31949) );
  NAND3X1 U26379 ( .A(n31972), .B(n31973), .C(n31974), .Y(n31971) );
  NOR2X1 U26380 ( .A(n31975), .B(n31976), .Y(n31974) );
  OAI22X1 U26381 ( .A(n25736), .B(n29655), .C(n25737), .D(n29989), .Y(n31976)
         );
  OAI22X1 U26382 ( .A(n25738), .B(n30015), .C(n25739), .D(n30007), .Y(n31975)
         );
  AOI22X1 U26383 ( .A(reg_A[56]), .B(n25615), .C(reg_A[59]), .D(n25616), .Y(
        n31973) );
  AOI22X1 U26384 ( .A(reg_A[58]), .B(n25607), .C(reg_A[62]), .D(n25608), .Y(
        n31972) );
  NAND3X1 U26385 ( .A(n31977), .B(n31978), .C(n31979), .Y(n31970) );
  NOR2X1 U26386 ( .A(n31980), .B(n31981), .Y(n31979) );
  OAI22X1 U26387 ( .A(n25745), .B(n30168), .C(n25746), .D(n30008), .Y(n31981)
         );
  OAI22X1 U26388 ( .A(n25747), .B(n30009), .C(n25748), .D(n30174), .Y(n31980)
         );
  AOI22X1 U26389 ( .A(reg_A[55]), .B(n25613), .C(reg_A[52]), .D(n25749), .Y(
        n31978) );
  AOI22X1 U26390 ( .A(reg_A[53]), .B(n25750), .C(reg_A[57]), .D(n25614), .Y(
        n31977) );
  OAI21X1 U26391 ( .A(n31982), .B(n31983), .C(n25310), .Y(n31948) );
  NAND3X1 U26392 ( .A(n31984), .B(n31985), .C(n31986), .Y(n31983) );
  NOR2X1 U26393 ( .A(n31987), .B(n31988), .Y(n31986) );
  OAI22X1 U26394 ( .A(n25043), .B(n29655), .C(n25039), .D(n29989), .Y(n31988)
         );
  OAI22X1 U26395 ( .A(n25064), .B(n30015), .C(n25065), .D(n30007), .Y(n31987)
         );
  AOI22X1 U26396 ( .A(reg_A[56]), .B(n25124), .C(reg_A[59]), .D(n25222), .Y(
        n31985) );
  AOI22X1 U26397 ( .A(reg_A[58]), .B(n25637), .C(reg_A[62]), .D(n25234), .Y(
        n31984) );
  NAND3X1 U26398 ( .A(n31989), .B(n31990), .C(n31991), .Y(n31982) );
  NOR2X1 U26399 ( .A(n31992), .B(n31993), .Y(n31991) );
  OAI22X1 U26400 ( .A(n25033), .B(n30168), .C(n25040), .D(n30008), .Y(n31993)
         );
  OAI22X1 U26401 ( .A(n25041), .B(n30009), .C(n25042), .D(n30174), .Y(n31992)
         );
  AOI22X1 U26402 ( .A(reg_A[55]), .B(n25628), .C(reg_A[52]), .D(n25068), .Y(
        n31990) );
  AOI22X1 U26403 ( .A(reg_A[53]), .B(n25123), .C(reg_A[57]), .D(n25629), .Y(
        n31989) );
  NOR2X1 U26404 ( .A(n31994), .B(n31995), .Y(n31931) );
  OAI21X1 U26405 ( .A(n31843), .B(n30198), .C(n31996), .Y(n31995) );
  OAI21X1 U26406 ( .A(n31997), .B(n31998), .C(n25382), .Y(n31996) );
  OAI22X1 U26407 ( .A(n31517), .B(n31628), .C(n31623), .D(n31999), .Y(n31998)
         );
  INVX1 U26408 ( .A(n32000), .Y(n31999) );
  AND2X1 U26409 ( .A(n25052), .B(n31039), .Y(n31623) );
  NAND2X1 U26410 ( .A(n25044), .B(n30341), .Y(n31039) );
  NAND2X1 U26411 ( .A(reg_B[53]), .B(n25029), .Y(n31628) );
  MUX2X1 U26412 ( .B(n32001), .A(n31726), .S(reg_B[54]), .Y(n31517) );
  MUX2X1 U26413 ( .B(n30043), .A(n30168), .S(n31338), .Y(n31726) );
  INVX1 U26414 ( .A(n31728), .Y(n32001) );
  MUX2X1 U26415 ( .B(reg_A[52]), .A(reg_A[53]), .S(reg_B[55]), .Y(n31728) );
  OAI21X1 U26416 ( .A(n31190), .B(n31516), .C(n32002), .Y(n31997) );
  AOI22X1 U26417 ( .A(n32003), .B(n31338), .C(n32004), .D(reg_A[49]), .Y(
        n32002) );
  INVX1 U26418 ( .A(n31719), .Y(n32004) );
  NAND2X1 U26419 ( .A(reg_B[55]), .B(n31194), .Y(n31719) );
  INVX1 U26420 ( .A(n31150), .Y(n31194) );
  INVX1 U26421 ( .A(reg_B[55]), .Y(n31338) );
  OAI22X1 U26422 ( .A(n30008), .B(n31190), .C(n29655), .D(n31150), .Y(n32003)
         );
  NAND2X1 U26423 ( .A(n31138), .B(n25029), .Y(n31150) );
  INVX1 U26424 ( .A(n31366), .Y(n31138) );
  NAND2X1 U26425 ( .A(n31369), .B(n31449), .Y(n31366) );
  INVX1 U26426 ( .A(reg_B[54]), .Y(n31449) );
  NAND2X1 U26427 ( .A(reg_B[55]), .B(reg_A[51]), .Y(n31516) );
  NAND2X1 U26428 ( .A(n31368), .B(n25029), .Y(n31190) );
  INVX1 U26429 ( .A(n31339), .Y(n31368) );
  NAND2X1 U26430 ( .A(reg_B[54]), .B(n31369), .Y(n31339) );
  INVX1 U26431 ( .A(reg_B[53]), .Y(n31369) );
  AND2X1 U26432 ( .A(n32005), .B(n32006), .Y(n31843) );
  AOI22X1 U26433 ( .A(n30024), .B(n31311), .C(n30141), .D(n31497), .Y(n32006)
         );
  OAI21X1 U26434 ( .A(n30744), .B(n30109), .C(n32007), .Y(n31311) );
  AOI22X1 U26435 ( .A(n30112), .B(reg_A[32]), .C(n30117), .D(reg_A[48]), .Y(
        n32007) );
  INVX1 U26436 ( .A(n31023), .Y(n30112) );
  AOI22X1 U26437 ( .A(n30201), .B(n31712), .C(n30342), .D(n32008), .Y(n32005)
         );
  OAI21X1 U26438 ( .A(n27919), .B(n30395), .C(n32009), .Y(n31994) );
  AOI22X1 U26439 ( .A(n26928), .B(n32010), .C(n32011), .D(n30341), .Y(n32009)
         );
  OAI21X1 U26440 ( .A(n30290), .B(n31898), .C(n32012), .Y(n32011) );
  AOI22X1 U26441 ( .A(n32013), .B(n30040), .C(n30120), .D(n32014), .Y(n32012)
         );
  OAI22X1 U26442 ( .A(n30021), .B(n30702), .C(n30256), .D(n30296), .Y(n32014)
         );
  MUX2X1 U26443 ( .B(reg_A[37]), .A(reg_A[45]), .S(n30853), .Y(n30296) );
  INVX1 U26444 ( .A(n31923), .Y(n30702) );
  MUX2X1 U26445 ( .B(n30160), .A(n30393), .S(reg_B[60]), .Y(n31923) );
  MUX2X1 U26446 ( .B(n30068), .A(n30059), .S(reg_B[60]), .Y(n30040) );
  NOR2X1 U26447 ( .A(n25024), .B(n29978), .Y(n32013) );
  OAI21X1 U26448 ( .A(reg_B[62]), .B(n31649), .C(n32015), .Y(n31898) );
  AOI22X1 U26449 ( .A(n32016), .B(n30342), .C(n30141), .D(n30243), .Y(n32015)
         );
  MUX2X1 U26450 ( .B(reg_A[38]), .A(reg_A[46]), .S(n30853), .Y(n30243) );
  MUX2X1 U26451 ( .B(reg_A[42]), .A(reg_A[34]), .S(reg_B[60]), .Y(n32016) );
  INVX1 U26452 ( .A(n32017), .Y(n31649) );
  OAI21X1 U26453 ( .A(reg_A[48]), .B(n29975), .C(n32018), .Y(n32017) );
  AOI22X1 U26454 ( .A(reg_B[61]), .B(n30513), .C(n30324), .D(n30744), .Y(
        n32018) );
  MUX2X1 U26455 ( .B(reg_A[36]), .A(reg_A[44]), .S(n30853), .Y(n30513) );
  OAI21X1 U26456 ( .A(n26944), .B(n30299), .C(n32019), .Y(n32010) );
  AOI22X1 U26457 ( .A(reg_A[54]), .B(n26010), .C(reg_A[55]), .D(n26002), .Y(
        n32019) );
  NOR2X1 U26458 ( .A(n25721), .B(n32020), .Y(n27919) );
  NOR2X1 U26459 ( .A(n32021), .B(n32022), .Y(n31930) );
  OAI22X1 U26460 ( .A(n25717), .B(n30008), .C(n25718), .D(n30009), .Y(n32022)
         );
  OAI21X1 U26461 ( .A(n25719), .B(n30174), .C(n32023), .Y(n32021) );
  AOI22X1 U26462 ( .A(n30261), .B(n32024), .C(reg_A[52]), .D(n25722), .Y(
        n32023) );
  NAND3X1 U26463 ( .A(n32025), .B(n32026), .C(n32027), .Y(result[47]) );
  NOR2X1 U26464 ( .A(n32028), .B(n32029), .Y(n32027) );
  NAND3X1 U26465 ( .A(n32030), .B(n32031), .C(n32032), .Y(n32029) );
  AOI21X1 U26466 ( .A(n32033), .B(n25935), .C(n32034), .Y(n32032) );
  OAI22X1 U26467 ( .A(n25941), .B(n32035), .C(n32036), .D(n32037), .Y(n32034)
         );
  OAI21X1 U26468 ( .A(n32038), .B(n32039), .C(n26480), .Y(n32031) );
  OAI22X1 U26469 ( .A(n32040), .B(n32041), .C(n32042), .D(n32043), .Y(n32039)
         );
  OAI22X1 U26470 ( .A(n32044), .B(n32045), .C(n32046), .D(n31023), .Y(n32038)
         );
  AOI22X1 U26471 ( .A(n25932), .B(n32047), .C(reg_A[46]), .D(n32048), .Y(
        n32030) );
  OAI21X1 U26472 ( .A(n32049), .B(n32050), .C(n32051), .Y(n32048) );
  NOR2X1 U26473 ( .A(n32052), .B(n32053), .Y(n32051) );
  OAI21X1 U26474 ( .A(n32054), .B(n29978), .C(n32055), .Y(n32047) );
  AOI22X1 U26475 ( .A(reg_B[61]), .B(n32056), .C(n30847), .D(n32057), .Y(
        n32055) );
  OAI22X1 U26476 ( .A(n30210), .B(n32058), .C(n32059), .D(n30320), .Y(n32056)
         );
  NAND3X1 U26477 ( .A(n32060), .B(n32061), .C(n32062), .Y(n32028) );
  NOR2X1 U26478 ( .A(n32063), .B(n32064), .Y(n32062) );
  OAI21X1 U26479 ( .A(n32065), .B(n32066), .C(n32067), .Y(n32064) );
  OAI21X1 U26480 ( .A(n32068), .B(n32069), .C(n25918), .Y(n32067) );
  NAND3X1 U26481 ( .A(n32070), .B(n32071), .C(n32072), .Y(n32069) );
  NOR2X1 U26482 ( .A(n32073), .B(n32074), .Y(n32072) );
  OAI22X1 U26483 ( .A(n25736), .B(n30068), .C(n25737), .D(n30394), .Y(n32074)
         );
  OAI22X1 U26484 ( .A(n25738), .B(n30393), .C(n25739), .D(n30395), .Y(n32073)
         );
  AOI22X1 U26485 ( .A(reg_A[39]), .B(n25615), .C(reg_A[36]), .D(n25616), .Y(
        n32071) );
  AOI22X1 U26486 ( .A(reg_A[37]), .B(n25607), .C(reg_A[33]), .D(n25608), .Y(
        n32070) );
  NAND3X1 U26487 ( .A(n32075), .B(n32076), .C(n32077), .Y(n32068) );
  NOR2X1 U26488 ( .A(n32078), .B(n32079), .Y(n32077) );
  OAI22X1 U26489 ( .A(n25061), .B(n30463), .C(n25746), .D(n30066), .Y(n32079)
         );
  OAI22X1 U26490 ( .A(n25747), .B(n30067), .C(n25748), .D(n30069), .Y(n32078)
         );
  AOI22X1 U26491 ( .A(reg_A[40]), .B(n25613), .C(reg_A[43]), .D(n25749), .Y(
        n32076) );
  AOI22X1 U26492 ( .A(reg_A[42]), .B(n25750), .C(reg_A[38]), .D(n25614), .Y(
        n32075) );
  AOI22X1 U26493 ( .A(n26267), .B(n32080), .C(n26186), .D(n32081), .Y(n32065)
         );
  INVX1 U26494 ( .A(n32082), .Y(n32063) );
  OAI21X1 U26495 ( .A(n32083), .B(n32084), .C(n25310), .Y(n32082) );
  NAND3X1 U26496 ( .A(n32085), .B(n32086), .C(n32087), .Y(n32084) );
  NOR2X1 U26497 ( .A(n32088), .B(n32089), .Y(n32087) );
  OAI22X1 U26498 ( .A(n25043), .B(n30068), .C(n25229), .D(n30015), .Y(n32089)
         );
  OAI22X1 U26499 ( .A(n25064), .B(n29984), .C(n25482), .D(n30016), .Y(n32088)
         );
  AOI22X1 U26500 ( .A(reg_A[55]), .B(n25124), .C(reg_A[58]), .D(n25222), .Y(
        n32086) );
  AOI22X1 U26501 ( .A(reg_A[57]), .B(n25637), .C(reg_A[61]), .D(n25234), .Y(
        n32085) );
  NAND3X1 U26502 ( .A(n32090), .B(n32091), .C(n32092), .Y(n32083) );
  NOR2X1 U26503 ( .A(n32093), .B(n32094), .Y(n32092) );
  OAI22X1 U26504 ( .A(n25033), .B(n30299), .C(n25040), .D(n30174), .Y(n32094)
         );
  OAI21X1 U26505 ( .A(n25041), .B(n30008), .C(n32095), .Y(n32093) );
  AOI22X1 U26506 ( .A(reg_A[63]), .B(n25247), .C(reg_A[48]), .D(n25135), .Y(
        n32095) );
  AOI22X1 U26507 ( .A(reg_A[54]), .B(n25628), .C(reg_A[51]), .D(n25069), .Y(
        n32091) );
  AOI22X1 U26508 ( .A(reg_A[52]), .B(n25123), .C(reg_A[56]), .D(n25629), .Y(
        n32090) );
  OAI21X1 U26509 ( .A(n32096), .B(n32097), .C(n25119), .Y(n32061) );
  NAND3X1 U26510 ( .A(n32098), .B(n32099), .C(n32100), .Y(n32097) );
  AOI21X1 U26511 ( .A(reg_A[47]), .B(n25125), .C(n32101), .Y(n32100) );
  OAI22X1 U26512 ( .A(n25039), .B(n30394), .C(n25231), .D(n30393), .Y(n32101)
         );
  AOI22X1 U26513 ( .A(reg_A[39]), .B(n25124), .C(reg_A[36]), .D(n25222), .Y(
        n32099) );
  AOI22X1 U26514 ( .A(reg_A[37]), .B(n25637), .C(reg_A[33]), .D(n25234), .Y(
        n32098) );
  NAND3X1 U26515 ( .A(n32102), .B(n32103), .C(n32104), .Y(n32096) );
  NOR2X1 U26516 ( .A(n32105), .B(n32106), .Y(n32104) );
  OAI22X1 U26517 ( .A(n25033), .B(n30463), .C(n25040), .D(n30066), .Y(n32106)
         );
  OAI22X1 U26518 ( .A(n25041), .B(n30067), .C(n25042), .D(n30069), .Y(n32105)
         );
  AOI22X1 U26519 ( .A(reg_A[40]), .B(n25628), .C(reg_A[43]), .D(n25069), .Y(
        n32103) );
  AOI22X1 U26520 ( .A(reg_A[42]), .B(n25123), .C(reg_A[38]), .D(n25629), .Y(
        n32102) );
  AOI21X1 U26521 ( .A(n32107), .B(reg_B[45]), .C(n31645), .Y(n32060) );
  NOR2X1 U26522 ( .A(n32108), .B(n25031), .Y(n32107) );
  AOI22X1 U26523 ( .A(n32109), .B(reg_A[42]), .C(n32110), .D(reg_A[43]), .Y(
        n32108) );
  NOR2X1 U26524 ( .A(n32111), .B(n32112), .Y(n32026) );
  OAI21X1 U26525 ( .A(n32113), .B(n30290), .C(n32114), .Y(n32112) );
  AOI22X1 U26526 ( .A(reg_A[43]), .B(n25948), .C(n32115), .D(n32116), .Y(
        n32114) );
  INVX1 U26527 ( .A(n32024), .Y(n32113) );
  OAI21X1 U26528 ( .A(n32117), .B(n30462), .C(n32118), .Y(n32111) );
  AOI21X1 U26529 ( .A(reg_A[47]), .B(n32119), .C(n32120), .Y(n32118) );
  AOI21X1 U26530 ( .A(n32121), .B(n32122), .C(n25697), .Y(n32120) );
  AOI22X1 U26531 ( .A(n32110), .B(n32123), .C(n30933), .D(n32024), .Y(n32122)
         );
  NAND2X1 U26532 ( .A(n32124), .B(n32125), .Y(n32024) );
  AOI22X1 U26533 ( .A(n30024), .B(n31373), .C(n30141), .D(n31578), .Y(n32125)
         );
  OAI22X1 U26534 ( .A(n30059), .B(n30109), .C(n29994), .D(n30068), .Y(n31373)
         );
  AOI22X1 U26535 ( .A(n30201), .B(n31847), .C(n30342), .D(n31955), .Y(n32124)
         );
  OAI21X1 U26536 ( .A(n30393), .B(n32126), .C(n32127), .Y(n32123) );
  AOI22X1 U26537 ( .A(n32128), .B(reg_A[43]), .C(n32129), .D(reg_A[39]), .Y(
        n32127) );
  AOI22X1 U26538 ( .A(n30862), .B(n32130), .C(n32131), .D(n32132), .Y(n32121)
         );
  INVX1 U26539 ( .A(n30095), .Y(n30862) );
  OAI21X1 U26540 ( .A(n32133), .B(n32134), .C(n32135), .Y(n32119) );
  INVX1 U26541 ( .A(n32136), .Y(n32133) );
  OAI21X1 U26542 ( .A(n32137), .B(n28105), .C(n32138), .Y(n32136) );
  NOR2X1 U26543 ( .A(n32139), .B(n32140), .Y(n32025) );
  OAI21X1 U26544 ( .A(n28066), .B(n30395), .C(n32141), .Y(n32140) );
  MUX2X1 U26545 ( .B(n32142), .A(n32143), .S(reg_B[46]), .Y(n32141) );
  NOR2X1 U26546 ( .A(n32144), .B(n25032), .Y(n32142) );
  AOI22X1 U26547 ( .A(n32145), .B(reg_B[45]), .C(n32146), .D(n32147), .Y(
        n32144) );
  NAND2X1 U26548 ( .A(n32148), .B(n32149), .Y(n32139) );
  OAI21X1 U26549 ( .A(n32150), .B(n32151), .C(n25999), .Y(n32149) );
  NAND2X1 U26550 ( .A(n32152), .B(n32153), .Y(n32151) );
  AOI22X1 U26551 ( .A(reg_A[40]), .B(n26002), .C(reg_A[43]), .D(n26003), .Y(
        n32153) );
  AOI22X1 U26552 ( .A(reg_A[42]), .B(n25751), .C(reg_A[47]), .D(n26004), .Y(
        n32152) );
  NAND2X1 U26553 ( .A(n32154), .B(n32155), .Y(n32150) );
  AOI22X1 U26554 ( .A(reg_A[46]), .B(n26007), .C(reg_A[44]), .D(n26008), .Y(
        n32155) );
  AOI22X1 U26555 ( .A(reg_A[45]), .B(n26009), .C(reg_A[41]), .D(n26010), .Y(
        n32154) );
  AOI22X1 U26556 ( .A(n32156), .B(n26262), .C(n32157), .D(n32158), .Y(n32148)
         );
  INVX1 U26557 ( .A(n32159), .Y(n32156) );
  NAND3X1 U26558 ( .A(n32160), .B(n32161), .C(n32162), .Y(result[46]) );
  NOR2X1 U26559 ( .A(n32163), .B(n32164), .Y(n32162) );
  NAND3X1 U26560 ( .A(n32165), .B(n32166), .C(n32167), .Y(n32164) );
  NOR2X1 U26561 ( .A(n32168), .B(n32169), .Y(n32167) );
  OAI21X1 U26562 ( .A(n28276), .B(n30067), .C(n32170), .Y(n32169) );
  OAI21X1 U26563 ( .A(n32171), .B(n32172), .C(n25119), .Y(n32170) );
  NAND3X1 U26564 ( .A(n32173), .B(n32174), .C(n32175), .Y(n32172) );
  AOI21X1 U26565 ( .A(reg_A[46]), .B(n25125), .C(n32176), .Y(n32175) );
  OAI22X1 U26566 ( .A(n25039), .B(n30170), .C(n25231), .D(n30394), .Y(n32176)
         );
  AOI22X1 U26567 ( .A(reg_A[37]), .B(n25629), .C(reg_A[38]), .D(n25124), .Y(
        n32174) );
  AOI22X1 U26568 ( .A(reg_A[35]), .B(n25222), .C(reg_A[36]), .D(n25637), .Y(
        n32173) );
  NAND3X1 U26569 ( .A(n32177), .B(n32178), .C(n32179), .Y(n32171) );
  AOI21X1 U26570 ( .A(reg_A[41]), .B(n25123), .C(n32180), .Y(n32179) );
  OAI22X1 U26571 ( .A(n26431), .B(n30462), .C(n25129), .D(n30059), .Y(n32180)
         );
  AOI22X1 U26572 ( .A(reg_A[45]), .B(n25135), .C(reg_A[43]), .D(n25136), .Y(
        n32178) );
  AOI22X1 U26573 ( .A(reg_A[44]), .B(n25252), .C(reg_A[40]), .D(n25253), .Y(
        n32177) );
  OAI22X1 U26574 ( .A(n32135), .B(n30069), .C(n30226), .D(n30462), .Y(n32168)
         );
  OAI21X1 U26575 ( .A(n32181), .B(n32182), .C(n26045), .Y(n32166) );
  NAND2X1 U26576 ( .A(n32183), .B(n32184), .Y(n32182) );
  AOI22X1 U26577 ( .A(reg_A[43]), .B(n25442), .C(reg_A[42]), .D(n27387), .Y(
        n32184) );
  AOI22X1 U26578 ( .A(reg_A[44]), .B(n28312), .C(reg_A[46]), .D(n25434), .Y(
        n32183) );
  NAND2X1 U26579 ( .A(n32185), .B(n32186), .Y(n32181) );
  AOI22X1 U26580 ( .A(reg_A[41]), .B(n30446), .C(reg_A[40]), .D(n25440), .Y(
        n32186) );
  INVX1 U26581 ( .A(n25449), .Y(n30446) );
  AOI22X1 U26582 ( .A(n25604), .B(n32187), .C(reg_A[45]), .D(n32188), .Y(
        n32185) );
  NAND3X1 U26583 ( .A(n32189), .B(n32190), .C(n32191), .Y(n32187) );
  NOR2X1 U26584 ( .A(n32192), .B(n32193), .Y(n32191) );
  OAI22X1 U26585 ( .A(n25737), .B(n30170), .C(n25738), .D(n30394), .Y(n32193)
         );
  OAI22X1 U26586 ( .A(n32194), .B(n30395), .C(n31398), .D(n30058), .Y(n32192)
         );
  AOI22X1 U26587 ( .A(reg_A[39]), .B(n25613), .C(reg_A[37]), .D(n25614), .Y(
        n32190) );
  AOI22X1 U26588 ( .A(reg_A[38]), .B(n25615), .C(reg_A[35]), .D(n25616), .Y(
        n32189) );
  AOI22X1 U26589 ( .A(n32157), .B(n32195), .C(n31076), .D(n32130), .Y(n32165)
         );
  NAND2X1 U26590 ( .A(n32196), .B(n32197), .Y(n32130) );
  AOI22X1 U26591 ( .A(n30141), .B(n31712), .C(n30024), .D(n31497), .Y(n32197)
         );
  INVX1 U26592 ( .A(n30256), .Y(n30141) );
  NAND2X1 U26593 ( .A(reg_B[62]), .B(n29973), .Y(n30256) );
  AOI22X1 U26594 ( .A(n30201), .B(n32008), .C(n30342), .D(n32198), .Y(n32196)
         );
  INVX1 U26595 ( .A(n30255), .Y(n30342) );
  NAND3X1 U26596 ( .A(n32199), .B(n32200), .C(n32201), .Y(n32163) );
  AOI21X1 U26597 ( .A(reg_A[41]), .B(n28282), .C(n32202), .Y(n32201) );
  OAI22X1 U26598 ( .A(n32203), .B(n30744), .C(n32204), .D(n30395), .Y(n32202)
         );
  AOI22X1 U26599 ( .A(n32205), .B(reg_B[46]), .C(reg_B[45]), .D(n32206), .Y(
        n32200) );
  AOI22X1 U26600 ( .A(n32207), .B(n26139), .C(reg_A[47]), .D(n28280), .Y(
        n32199) );
  NOR2X1 U26601 ( .A(n32208), .B(n32209), .Y(n32161) );
  NAND3X1 U26602 ( .A(n32210), .B(n32211), .C(n32212), .Y(n32209) );
  OAI21X1 U26603 ( .A(n32213), .B(n32214), .C(n25932), .Y(n32212) );
  OAI22X1 U26604 ( .A(n30255), .B(n32058), .C(n32059), .D(n30032), .Y(n32214)
         );
  OAI22X1 U26605 ( .A(n32054), .B(n30103), .C(n32215), .D(n30038), .Y(n32213)
         );
  INVX1 U26606 ( .A(n32057), .Y(n32215) );
  OAI21X1 U26607 ( .A(reg_B[61]), .B(n32216), .C(n32217), .Y(n32057) );
  INVX1 U26608 ( .A(n31497), .Y(n32054) );
  OAI22X1 U26609 ( .A(n30060), .B(n30109), .C(n29994), .D(n30069), .Y(n31497)
         );
  OAI21X1 U26610 ( .A(n32218), .B(n32219), .C(n32220), .Y(n32211) );
  INVX1 U26611 ( .A(n32221), .Y(n32218) );
  OAI21X1 U26612 ( .A(n30120), .B(n30261), .C(n32222), .Y(n32210) );
  INVX1 U26613 ( .A(n30233), .Y(n30120) );
  NAND2X1 U26614 ( .A(reg_B[63]), .B(n25932), .Y(n30233) );
  NAND3X1 U26615 ( .A(n32223), .B(n31954), .C(n32224), .Y(n32208) );
  AOI22X1 U26616 ( .A(n32225), .B(n26186), .C(n32226), .D(n32227), .Y(n32224)
         );
  NOR2X1 U26617 ( .A(n25032), .B(n32228), .Y(n32226) );
  AND2X1 U26618 ( .A(n32229), .B(n32132), .Y(n32225) );
  OAI21X1 U26619 ( .A(n30069), .B(n32049), .C(n32230), .Y(n32132) );
  MUX2X1 U26620 ( .B(n32231), .A(n32232), .S(reg_B[46]), .Y(n32230) );
  NOR2X1 U26621 ( .A(n30462), .B(n32233), .Y(n32231) );
  NAND3X1 U26622 ( .A(n32081), .B(n29315), .C(n32109), .Y(n32223) );
  NOR2X1 U26623 ( .A(n32234), .B(n32235), .Y(n32160) );
  NAND3X1 U26624 ( .A(n32236), .B(n32237), .C(n32238), .Y(n32235) );
  OAI21X1 U26625 ( .A(n28206), .B(n32239), .C(reg_A[43]), .Y(n32238) );
  OAI21X1 U26626 ( .A(n32138), .B(n32240), .C(n32241), .Y(n32239) );
  NAND3X1 U26627 ( .A(reg_B[47]), .B(n26186), .C(n32242), .Y(n32241) );
  OAI21X1 U26628 ( .A(n32243), .B(n32244), .C(n26480), .Y(n32237) );
  OAI22X1 U26629 ( .A(n32245), .B(n32043), .C(n32246), .D(n32045), .Y(n32244)
         );
  OAI22X1 U26630 ( .A(n30870), .B(n32041), .C(n30257), .D(n32247), .Y(n32243)
         );
  INVX1 U26631 ( .A(n32248), .Y(n30257) );
  INVX1 U26632 ( .A(n32249), .Y(n30870) );
  OAI21X1 U26633 ( .A(n32250), .B(n32251), .C(n26267), .Y(n32236) );
  OAI22X1 U26634 ( .A(n32252), .B(n32253), .C(reg_B[47]), .D(n32036), .Y(
        n32251) );
  MUX2X1 U26635 ( .B(n32254), .A(n32255), .S(reg_B[46]), .Y(n32036) );
  INVX1 U26636 ( .A(n32256), .Y(n32255) );
  NAND2X1 U26637 ( .A(n32257), .B(n32258), .Y(n32254) );
  AOI22X1 U26638 ( .A(n32259), .B(reg_B[44]), .C(n32147), .D(reg_A[38]), .Y(
        n32258) );
  NOR2X1 U26639 ( .A(n30394), .B(n32233), .Y(n32259) );
  AOI22X1 U26640 ( .A(n32260), .B(reg_A[42]), .C(n32261), .D(reg_A[46]), .Y(
        n32257) );
  NOR2X1 U26641 ( .A(n32262), .B(n32240), .Y(n32250) );
  NAND3X1 U26642 ( .A(n32263), .B(n32264), .C(n32265), .Y(n32234) );
  AOI22X1 U26643 ( .A(n32266), .B(n28253), .C(n32267), .D(n32268), .Y(n32265)
         );
  OAI21X1 U26644 ( .A(n32269), .B(n32270), .C(n25310), .Y(n32264) );
  NAND3X1 U26645 ( .A(n32271), .B(n32272), .C(n32273), .Y(n32270) );
  NOR2X1 U26646 ( .A(n32274), .B(n32275), .Y(n32273) );
  OAI22X1 U26647 ( .A(n25035), .B(n30015), .C(n25036), .D(n30254), .Y(n32275)
         );
  OAI21X1 U26648 ( .A(n25027), .B(n29990), .C(n32276), .Y(n32274) );
  AOI22X1 U26649 ( .A(reg_A[55]), .B(n25629), .C(reg_A[54]), .D(n25124), .Y(
        n32276) );
  AOI22X1 U26650 ( .A(reg_A[61]), .B(n25235), .C(reg_A[58]), .D(n25635), .Y(
        n32272) );
  AOI22X1 U26651 ( .A(reg_A[59]), .B(n25325), .C(reg_A[46]), .D(n25125), .Y(
        n32271) );
  NAND3X1 U26652 ( .A(n32277), .B(n32278), .C(n32279), .Y(n32269) );
  NOR2X1 U26653 ( .A(n32280), .B(n32281), .Y(n32279) );
  OAI22X1 U26654 ( .A(n25040), .B(n29655), .C(n25254), .D(n30174), .Y(n32281)
         );
  OAI21X1 U26655 ( .A(n25042), .B(n30068), .C(n32282), .Y(n32280) );
  AOI22X1 U26656 ( .A(reg_A[63]), .B(n25246), .C(reg_A[62]), .D(n25247), .Y(
        n32282) );
  AOI22X1 U26657 ( .A(reg_A[52]), .B(n25253), .C(reg_A[53]), .D(n25628), .Y(
        n32278) );
  AOI22X1 U26658 ( .A(reg_A[50]), .B(n25072), .C(reg_A[51]), .D(n25123), .Y(
        n32277) );
  OAI21X1 U26659 ( .A(n32053), .B(n28332), .C(reg_A[45]), .Y(n32263) );
  NOR2X1 U26660 ( .A(n32283), .B(n32253), .Y(n32053) );
  NAND3X1 U26661 ( .A(n32284), .B(n32285), .C(n32286), .Y(result[45]) );
  NOR2X1 U26662 ( .A(n32287), .B(n32288), .Y(n32286) );
  NAND3X1 U26663 ( .A(n32289), .B(n32290), .C(n32291), .Y(n32288) );
  AOI21X1 U26664 ( .A(reg_A[40]), .B(n32292), .C(n32293), .Y(n32291) );
  OAI21X1 U26665 ( .A(n32294), .B(n26147), .C(n32295), .Y(n32293) );
  OAI21X1 U26666 ( .A(n32296), .B(n32297), .C(n25932), .Y(n32295) );
  OAI22X1 U26667 ( .A(n32298), .B(n30210), .C(n32216), .D(n29978), .Y(n32297)
         );
  OAI22X1 U26668 ( .A(n31459), .B(n32058), .C(n30320), .D(n32217), .Y(n32296)
         );
  AOI21X1 U26669 ( .A(n32299), .B(n32300), .C(n32301), .Y(n32294) );
  OAI22X1 U26670 ( .A(n32256), .B(n32253), .C(n32252), .D(n32134), .Y(n32301)
         );
  INVX1 U26671 ( .A(n32080), .Y(n32252) );
  NAND2X1 U26672 ( .A(n32302), .B(n32303), .Y(n32080) );
  AOI22X1 U26673 ( .A(n32304), .B(reg_B[44]), .C(n32147), .D(reg_A[37]), .Y(
        n32303) );
  NOR2X1 U26674 ( .A(n30170), .B(n32233), .Y(n32304) );
  AOI22X1 U26675 ( .A(n32260), .B(reg_A[41]), .C(n32261), .D(reg_A[45]), .Y(
        n32302) );
  OAI21X1 U26676 ( .A(n32305), .B(n32306), .C(n26480), .Y(n32290) );
  OAI22X1 U26677 ( .A(n32307), .B(n32043), .C(n32308), .D(n32045), .Y(n32306)
         );
  OAI22X1 U26678 ( .A(n30889), .B(n32041), .C(n32309), .D(n32247), .Y(n32305)
         );
  INVX1 U26679 ( .A(n30285), .Y(n32309) );
  INVX1 U26680 ( .A(n32310), .Y(n30889) );
  AOI22X1 U26681 ( .A(reg_A[32]), .B(n28453), .C(n32311), .D(n32312), .Y(
        n32289) );
  OR2X1 U26682 ( .A(n32313), .B(n32314), .Y(n32287) );
  OAI21X1 U26683 ( .A(n32315), .B(n32316), .C(n32317), .Y(n32314) );
  AOI22X1 U26684 ( .A(reg_A[43]), .B(n32318), .C(n32115), .D(n32319), .Y(
        n32317) );
  AND2X1 U26685 ( .A(n32320), .B(n32321), .Y(n32115) );
  AOI22X1 U26686 ( .A(n26292), .B(n30463), .C(n26293), .D(n30066), .Y(n32321)
         );
  AOI22X1 U26687 ( .A(n26294), .B(n30744), .C(n26295), .D(n30067), .Y(n32320)
         );
  OAI21X1 U26688 ( .A(n32066), .B(n32322), .C(n28415), .Y(n32318) );
  NAND3X1 U26689 ( .A(n32323), .B(n31954), .C(n32324), .Y(n32313) );
  OAI21X1 U26690 ( .A(n32325), .B(n32326), .C(n25170), .Y(n32324) );
  OAI22X1 U26691 ( .A(n32327), .B(n30095), .C(n32328), .D(n30327), .Y(n32326)
         );
  INVX1 U26692 ( .A(n32329), .Y(n32327) );
  OAI22X1 U26693 ( .A(n32330), .B(n32331), .C(n32332), .D(n32333), .Y(n32325)
         );
  AOI22X1 U26694 ( .A(n32081), .B(n32334), .C(n32242), .D(reg_A[43]), .Y(
        n32332) );
  OAI21X1 U26695 ( .A(n32335), .B(n32336), .C(n25310), .Y(n32323) );
  NAND3X1 U26696 ( .A(n32337), .B(n32338), .C(n32339), .Y(n32336) );
  NOR2X1 U26697 ( .A(n32340), .B(n32341), .Y(n32339) );
  OAI22X1 U26698 ( .A(n25035), .B(n29984), .C(n25036), .D(n30043), .Y(n32341)
         );
  OAI21X1 U26699 ( .A(n25027), .B(n30254), .C(n32342), .Y(n32340) );
  AOI22X1 U26700 ( .A(reg_A[54]), .B(n25629), .C(reg_A[53]), .D(n25124), .Y(
        n32342) );
  AOI22X1 U26701 ( .A(reg_A[60]), .B(n25235), .C(reg_A[57]), .D(n25635), .Y(
        n32338) );
  AOI22X1 U26702 ( .A(reg_A[58]), .B(n25325), .C(reg_A[45]), .D(n25125), .Y(
        n32337) );
  NAND3X1 U26703 ( .A(n32343), .B(n32344), .C(n32345), .Y(n32335) );
  NOR2X1 U26704 ( .A(n32346), .B(n32347), .Y(n32345) );
  OAI22X1 U26705 ( .A(n25041), .B(n29655), .C(n25784), .D(n30069), .Y(n32347)
         );
  OAI21X1 U26706 ( .A(n25051), .B(n30007), .C(n32348), .Y(n32346) );
  AOI22X1 U26707 ( .A(reg_A[62]), .B(n25246), .C(reg_A[61]), .D(n25247), .Y(
        n32348) );
  AOI21X1 U26708 ( .A(reg_A[52]), .B(n25628), .C(n32349), .Y(n32344) );
  OAI22X1 U26709 ( .A(n25033), .B(n30009), .C(n25040), .D(n30068), .Y(n32349)
         );
  AOI22X1 U26710 ( .A(reg_A[49]), .B(n25072), .C(reg_A[50]), .D(n25123), .Y(
        n32343) );
  NOR2X1 U26711 ( .A(n32350), .B(n32351), .Y(n32285) );
  OAI21X1 U26712 ( .A(n32328), .B(n30290), .C(n32352), .Y(n32351) );
  AOI22X1 U26713 ( .A(reg_A[47]), .B(n25153), .C(reg_A[46]), .D(n28280), .Y(
        n32352) );
  INVX1 U26714 ( .A(n32222), .Y(n32328) );
  OAI21X1 U26715 ( .A(n32353), .B(n30293), .C(n32354), .Y(n32222) );
  AOI22X1 U26716 ( .A(n30024), .B(n31578), .C(n30201), .D(n31955), .Y(n32354)
         );
  OAI22X1 U26717 ( .A(n30057), .B(n30109), .C(n29994), .D(n30066), .Y(n31578)
         );
  OAI21X1 U26718 ( .A(n26854), .B(n32159), .C(n32355), .Y(n32350) );
  AOI22X1 U26719 ( .A(reg_A[42]), .B(n32356), .C(n32357), .D(n32358), .Y(
        n32355) );
  OAI21X1 U26720 ( .A(n32359), .B(n26452), .C(n32360), .Y(n32159) );
  AOI22X1 U26721 ( .A(n26293), .B(n30308), .C(n26295), .D(n30536), .Y(n32360)
         );
  INVX1 U26722 ( .A(n31704), .Y(n30536) );
  MUX2X1 U26723 ( .B(n30067), .A(n30058), .S(reg_B[1]), .Y(n31704) );
  INVX1 U26724 ( .A(n31947), .Y(n30308) );
  MUX2X1 U26725 ( .B(n30066), .A(n30057), .S(reg_B[1]), .Y(n31947) );
  INVX1 U26726 ( .A(n32361), .Y(n32359) );
  NOR2X1 U26727 ( .A(n32362), .B(n32363), .Y(n32284) );
  NAND2X1 U26728 ( .A(n32364), .B(n32365), .Y(n32363) );
  MUX2X1 U26729 ( .B(n32143), .A(n32205), .S(reg_B[46]), .Y(n32365) );
  OAI22X1 U26730 ( .A(n32366), .B(n32367), .C(n25342), .D(n32368), .Y(n32143)
         );
  MUX2X1 U26731 ( .B(n32081), .A(n32232), .S(reg_B[47]), .Y(n32368) );
  MUX2X1 U26732 ( .B(n30463), .A(n30066), .S(n32233), .Y(n32081) );
  OAI21X1 U26733 ( .A(n32369), .B(n32233), .C(n25188), .Y(n32367) );
  OAI22X1 U26734 ( .A(n32370), .B(n32228), .C(n32371), .D(n32372), .Y(n32366)
         );
  MUX2X1 U26735 ( .B(n30066), .A(n30067), .S(reg_B[47]), .Y(n32372) );
  AOI22X1 U26736 ( .A(n27676), .B(n32373), .C(reg_A[45]), .D(n28343), .Y(
        n32364) );
  OAI21X1 U26737 ( .A(n32374), .B(n27523), .C(n32375), .Y(n32362) );
  AOI22X1 U26738 ( .A(n32376), .B(n26262), .C(n32157), .D(n32377), .Y(n32375)
         );
  INVX1 U26739 ( .A(n32378), .Y(n32376) );
  NOR2X1 U26740 ( .A(n32379), .B(n32380), .Y(n32374) );
  NAND3X1 U26741 ( .A(n32381), .B(n32382), .C(n32383), .Y(n32380) );
  AOI21X1 U26742 ( .A(reg_A[45]), .B(n25434), .C(n32384), .Y(n32383) );
  OAI22X1 U26743 ( .A(n28353), .B(n30160), .C(n25205), .D(n30463), .Y(n32384)
         );
  AOI22X1 U26744 ( .A(n25097), .B(n32373), .C(reg_A[40]), .D(n28355), .Y(
        n32382) );
  NAND3X1 U26745 ( .A(n32385), .B(n32386), .C(n32387), .Y(n32373) );
  NOR2X1 U26746 ( .A(n32388), .B(n32389), .Y(n32387) );
  OAI21X1 U26747 ( .A(n25043), .B(n30066), .C(n32390), .Y(n32389) );
  AOI22X1 U26748 ( .A(reg_A[35]), .B(n25637), .C(reg_A[33]), .D(n25635), .Y(
        n32390) );
  OAI21X1 U26749 ( .A(n25027), .B(n30394), .C(n32391), .Y(n32388) );
  AOI22X1 U26750 ( .A(reg_A[36]), .B(n25629), .C(reg_A[37]), .D(n25124), .Y(
        n32391) );
  NOR2X1 U26751 ( .A(n32392), .B(n32393), .Y(n32386) );
  OAI22X1 U26752 ( .A(n25033), .B(n30059), .C(n25040), .D(n30160), .Y(n32393)
         );
  OAI22X1 U26753 ( .A(n25041), .B(n30462), .C(n25784), .D(n30067), .Y(n32392)
         );
  AOI21X1 U26754 ( .A(reg_A[40]), .B(n25123), .C(n32394), .Y(n32385) );
  OAI22X1 U26755 ( .A(n26431), .B(n30463), .C(n25129), .D(n30060), .Y(n32394)
         );
  AOI22X1 U26756 ( .A(reg_A[44]), .B(n25441), .C(reg_A[42]), .D(n27241), .Y(
        n32381) );
  NAND3X1 U26757 ( .A(n32395), .B(n32396), .C(n32397), .Y(n32379) );
  NOR2X1 U26758 ( .A(n32398), .B(n32399), .Y(n32397) );
  OAI22X1 U26759 ( .A(n28361), .B(n30395), .C(n28311), .D(n30059), .Y(n32399)
         );
  OAI22X1 U26760 ( .A(n28362), .B(n30393), .C(n28363), .D(n30394), .Y(n32398)
         );
  AOI22X1 U26761 ( .A(reg_A[33]), .B(n28364), .C(reg_A[36]), .D(n25500), .Y(
        n32396) );
  AOI22X1 U26762 ( .A(reg_A[37]), .B(n25501), .C(reg_A[38]), .D(n25502), .Y(
        n32395) );
  NAND2X1 U26763 ( .A(n32400), .B(n32401), .Y(result[44]) );
  NOR2X1 U26764 ( .A(n32402), .B(n32403), .Y(n32401) );
  NAND2X1 U26765 ( .A(n32404), .B(n32405), .Y(n32403) );
  NOR2X1 U26766 ( .A(n32406), .B(n32407), .Y(n32405) );
  OAI21X1 U26767 ( .A(n32408), .B(n27438), .C(n32409), .Y(n32407) );
  OAI21X1 U26768 ( .A(n32410), .B(n32411), .C(n26267), .Y(n32409) );
  OAI22X1 U26769 ( .A(n32412), .B(n32240), .C(n32413), .D(n32066), .Y(n32411)
         );
  OAI22X1 U26770 ( .A(n32262), .B(n32253), .C(n32256), .D(n32134), .Y(n32410)
         );
  NOR2X1 U26771 ( .A(n32414), .B(n32415), .Y(n32256) );
  OAI22X1 U26772 ( .A(n30744), .B(n32416), .C(n30067), .D(n32371), .Y(n32415)
         );
  OAI21X1 U26773 ( .A(n30058), .B(n32228), .C(n32417), .Y(n32414) );
  NOR2X1 U26774 ( .A(n32418), .B(n32419), .Y(n32408) );
  OAI22X1 U26775 ( .A(n29973), .B(n32058), .C(n32298), .D(n30038), .Y(n32419)
         );
  OAI22X1 U26776 ( .A(n32216), .B(n30103), .C(n29970), .D(n32217), .Y(n32418)
         );
  NAND2X1 U26777 ( .A(n32420), .B(reg_A[40]), .Y(n32217) );
  INVX1 U26778 ( .A(n31712), .Y(n32216) );
  OAI21X1 U26779 ( .A(n32138), .B(n32421), .C(n32422), .Y(n32406) );
  OAI21X1 U26780 ( .A(n32423), .B(n32424), .C(n26480), .Y(n32422) );
  OAI22X1 U26781 ( .A(n32425), .B(n32043), .C(n32426), .D(n32041), .Y(n32424)
         );
  INVX1 U26782 ( .A(n32427), .Y(n32425) );
  OAI22X1 U26783 ( .A(n32428), .B(n32045), .C(n30521), .D(n32247), .Y(n32423)
         );
  AOI21X1 U26784 ( .A(n32110), .B(reg_A[44]), .C(n32429), .Y(n32421) );
  OAI22X1 U26785 ( .A(n30463), .B(n32240), .C(n30462), .D(n32066), .Y(n32429)
         );
  INVX1 U26786 ( .A(n32220), .Y(n32138) );
  NAND2X1 U26787 ( .A(n32322), .B(n32283), .Y(n32220) );
  NOR2X1 U26788 ( .A(n32430), .B(n32431), .Y(n32404) );
  OAI22X1 U26789 ( .A(n32432), .B(n30462), .C(n32433), .D(n30463), .Y(n32431)
         );
  OAI21X1 U26790 ( .A(n32434), .B(n30395), .C(n32435), .Y(n32430) );
  OAI21X1 U26791 ( .A(n32436), .B(n32437), .C(n25188), .Y(n32435) );
  OAI22X1 U26792 ( .A(n32416), .B(n32438), .C(n32228), .D(n32439), .Y(n32437)
         );
  OAI21X1 U26793 ( .A(n32371), .B(n32440), .C(n32417), .Y(n32436) );
  INVX1 U26794 ( .A(n28494), .Y(n32434) );
  NAND3X1 U26795 ( .A(n32441), .B(n32442), .C(n32443), .Y(n32402) );
  NOR2X1 U26796 ( .A(n32444), .B(n32445), .Y(n32443) );
  OAI21X1 U26797 ( .A(n25198), .B(n32446), .C(n32447), .Y(n32445) );
  OAI21X1 U26798 ( .A(n32448), .B(n32449), .C(n25310), .Y(n32447) );
  NAND3X1 U26799 ( .A(n32450), .B(n32451), .C(n32452), .Y(n32449) );
  NOR2X1 U26800 ( .A(n32453), .B(n32454), .Y(n32452) );
  OAI22X1 U26801 ( .A(n25043), .B(n30067), .C(n25039), .D(n29990), .Y(n32454)
         );
  OAI21X1 U26802 ( .A(n25064), .B(n30254), .C(n32455), .Y(n32453) );
  AOI22X1 U26803 ( .A(reg_A[58]), .B(n25234), .C(reg_A[59]), .D(n25235), .Y(
        n32455) );
  AOI21X1 U26804 ( .A(reg_A[52]), .B(n25124), .C(n32456), .Y(n32451) );
  OAI22X1 U26805 ( .A(n25037), .B(n30299), .C(n25028), .D(n30174), .Y(n32456)
         );
  AOI22X1 U26806 ( .A(reg_A[55]), .B(n25222), .C(reg_A[54]), .D(n25637), .Y(
        n32450) );
  NAND3X1 U26807 ( .A(n32457), .B(n32458), .C(n32459), .Y(n32448) );
  NOR2X1 U26808 ( .A(n32460), .B(n32461), .Y(n32459) );
  OAI22X1 U26809 ( .A(n25042), .B(n30066), .C(n25331), .D(n30016), .Y(n32461)
         );
  OAI21X1 U26810 ( .A(n25038), .B(n30007), .C(n32462), .Y(n32460) );
  AOI22X1 U26811 ( .A(reg_A[61]), .B(n25246), .C(reg_A[60]), .D(n25247), .Y(
        n32462) );
  AOI21X1 U26812 ( .A(reg_A[50]), .B(n25253), .C(n32463), .Y(n32458) );
  OAI22X1 U26813 ( .A(n25040), .B(n30069), .C(n25254), .D(n30068), .Y(n32463)
         );
  AOI22X1 U26814 ( .A(reg_A[51]), .B(n25628), .C(reg_A[48]), .D(n25067), .Y(
        n32457) );
  AOI22X1 U26815 ( .A(n30212), .B(n32464), .C(n30847), .D(n32465), .Y(n32446)
         );
  OAI21X1 U26816 ( .A(n32466), .B(n32050), .C(n32467), .Y(n32444) );
  OAI21X1 U26817 ( .A(n32468), .B(n32469), .C(n25119), .Y(n32467) );
  OR2X1 U26818 ( .A(n32470), .B(n32471), .Y(n32469) );
  OAI21X1 U26819 ( .A(n25034), .B(n30058), .C(n32472), .Y(n32471) );
  AOI22X1 U26820 ( .A(reg_A[38]), .B(n25253), .C(reg_A[37]), .D(n25628), .Y(
        n32472) );
  OAI21X1 U26821 ( .A(n25036), .B(n30394), .C(n32473), .Y(n32470) );
  AOI22X1 U26822 ( .A(reg_A[35]), .B(n25629), .C(reg_A[33]), .D(n25222), .Y(
        n32473) );
  OR2X1 U26823 ( .A(n32474), .B(n32475), .Y(n32468) );
  OAI21X1 U26824 ( .A(n25043), .B(n30067), .C(n32476), .Y(n32475) );
  AOI22X1 U26825 ( .A(reg_A[43]), .B(n25135), .C(reg_A[42]), .D(n25252), .Y(
        n32476) );
  OAI21X1 U26826 ( .A(n25028), .B(n30059), .C(n32477), .Y(n32474) );
  AOI22X1 U26827 ( .A(reg_A[41]), .B(n25136), .C(reg_A[40]), .D(n25068), .Y(
        n32477) );
  NAND2X1 U26828 ( .A(reg_B[47]), .B(n26504), .Y(n32050) );
  AOI22X1 U26829 ( .A(n32267), .B(n32478), .C(reg_A[33]), .D(n28549), .Y(
        n32442) );
  AOI22X1 U26830 ( .A(reg_A[34]), .B(n28649), .C(n25170), .D(n32479), .Y(
        n32441) );
  OAI21X1 U26831 ( .A(n32480), .B(n32331), .C(n32481), .Y(n32479) );
  AOI22X1 U26832 ( .A(n32482), .B(n32483), .C(n30933), .D(n32329), .Y(n32481)
         );
  OAI21X1 U26833 ( .A(n32298), .B(n30293), .C(n32484), .Y(n32329) );
  AOI22X1 U26834 ( .A(n30201), .B(n32198), .C(n30024), .D(n31712), .Y(n32484)
         );
  OAI22X1 U26835 ( .A(n30058), .B(n30109), .C(n29994), .D(n30067), .Y(n31712)
         );
  INVX1 U26836 ( .A(n30021), .Y(n30201) );
  NAND2X1 U26837 ( .A(reg_B[61]), .B(n30293), .Y(n30021) );
  INVX1 U26838 ( .A(n32485), .Y(n32298) );
  INVX1 U26839 ( .A(n30327), .Y(n30933) );
  INVX1 U26840 ( .A(n32330), .Y(n32483) );
  AOI22X1 U26841 ( .A(reg_A[42]), .B(n32242), .C(n32334), .D(n32232), .Y(
        n32330) );
  MUX2X1 U26842 ( .B(n30067), .A(n30744), .S(reg_B[45]), .Y(n32232) );
  INVX1 U26843 ( .A(n32486), .Y(n32242) );
  NOR2X1 U26844 ( .A(n32487), .B(n32488), .Y(n32400) );
  NAND3X1 U26845 ( .A(n32489), .B(n32490), .C(n32491), .Y(n32488) );
  NOR2X1 U26846 ( .A(n32492), .B(n32493), .Y(n32491) );
  OAI22X1 U26847 ( .A(n32494), .B(n30744), .C(n32495), .D(n30067), .Y(n32493)
         );
  OAI22X1 U26848 ( .A(n32496), .B(n30160), .C(n25148), .D(n30066), .Y(n32492)
         );
  AOI22X1 U26849 ( .A(n32157), .B(n32497), .C(reg_A[37]), .D(n32498), .Y(
        n32489) );
  NAND3X1 U26850 ( .A(n32499), .B(n32500), .C(n32501), .Y(n32487) );
  NOR2X1 U26851 ( .A(n32502), .B(n32503), .Y(n32501) );
  OAI22X1 U26852 ( .A(n28569), .B(n30069), .C(n28570), .D(n30068), .Y(n32503)
         );
  OAI22X1 U26853 ( .A(n28571), .B(n30059), .C(n25178), .D(n30058), .Y(n32502)
         );
  AOI22X1 U26854 ( .A(reg_A[35]), .B(n28572), .C(n32504), .D(n26139), .Y(
        n32500) );
  AOI22X1 U26855 ( .A(n32505), .B(n28575), .C(reg_A[38]), .D(n28576), .Y(
        n32499) );
  INVX1 U26856 ( .A(n32506), .Y(n32505) );
  NAND2X1 U26857 ( .A(n32507), .B(n32508), .Y(result[43]) );
  NOR2X1 U26858 ( .A(n32509), .B(n32510), .Y(n32508) );
  NAND3X1 U26859 ( .A(n32511), .B(n32512), .C(n32513), .Y(n32510) );
  NOR2X1 U26860 ( .A(n32514), .B(n32515), .Y(n32513) );
  OAI21X1 U26861 ( .A(n32516), .B(n30210), .C(n32517), .Y(n32515) );
  OAI21X1 U26862 ( .A(n32518), .B(n32519), .C(n26267), .Y(n32517) );
  OAI22X1 U26863 ( .A(n32412), .B(n32066), .C(n32262), .D(n32134), .Y(n32519)
         );
  INVX1 U26864 ( .A(n32300), .Y(n32262) );
  OAI21X1 U26865 ( .A(n30160), .B(n32371), .C(n32520), .Y(n32300) );
  AOI22X1 U26866 ( .A(n32147), .B(reg_A[35]), .C(n32260), .D(reg_A[39]), .Y(
        n32520) );
  NOR2X1 U26867 ( .A(n32521), .B(n32240), .Y(n32518) );
  OAI21X1 U26868 ( .A(n32522), .B(n30395), .C(n32523), .Y(n32514) );
  OAI21X1 U26869 ( .A(n32524), .B(n32525), .C(n26480), .Y(n32523) );
  OAI22X1 U26870 ( .A(n32042), .B(n32041), .C(n32044), .D(n32043), .Y(n32525)
         );
  INVX1 U26871 ( .A(n32526), .Y(n32042) );
  OAI22X1 U26872 ( .A(n32527), .B(n32045), .C(n30677), .D(n31023), .Y(n32524)
         );
  NAND2X1 U26873 ( .A(reg_B[59]), .B(n30853), .Y(n31023) );
  AOI22X1 U26874 ( .A(n32109), .B(n32358), .C(reg_A[41]), .D(n32528), .Y(
        n32512) );
  OAI22X1 U26875 ( .A(n32413), .B(n26147), .C(n30462), .D(n32322), .Y(n32358)
         );
  AOI22X1 U26876 ( .A(reg_A[34]), .B(n28572), .C(reg_A[37]), .D(n28576), .Y(
        n32511) );
  NAND3X1 U26877 ( .A(n32529), .B(n32530), .C(n32531), .Y(n32509) );
  NOR2X1 U26878 ( .A(n32532), .B(n32533), .Y(n32531) );
  OAI21X1 U26879 ( .A(n32534), .B(n25697), .C(n32535), .Y(n32533) );
  OAI21X1 U26880 ( .A(n32536), .B(n32537), .C(n25310), .Y(n32535) );
  NAND3X1 U26881 ( .A(n32538), .B(n32539), .C(n32540), .Y(n32537) );
  NOR2X1 U26882 ( .A(n32541), .B(n32542), .Y(n32540) );
  OAI22X1 U26883 ( .A(n25043), .B(n30160), .C(n25039), .D(n30254), .Y(n32542)
         );
  OAI21X1 U26884 ( .A(n25064), .B(n30043), .C(n32543), .Y(n32541) );
  AOI22X1 U26885 ( .A(reg_A[57]), .B(n25234), .C(reg_A[58]), .D(n25235), .Y(
        n32543) );
  AOI21X1 U26886 ( .A(reg_A[51]), .B(n25124), .C(n32544), .Y(n32539) );
  OAI22X1 U26887 ( .A(n25037), .B(n30378), .C(n26703), .D(n29655), .Y(n32544)
         );
  AOI22X1 U26888 ( .A(reg_A[54]), .B(n25222), .C(reg_A[53]), .D(n25637), .Y(
        n32538) );
  NAND3X1 U26889 ( .A(n32545), .B(n32546), .C(n32547), .Y(n32536) );
  NOR2X1 U26890 ( .A(n32548), .B(n32549), .Y(n32547) );
  OAI21X1 U26891 ( .A(n25042), .B(n30067), .C(n32550), .Y(n32549) );
  AOI22X1 U26892 ( .A(reg_A[61]), .B(n25241), .C(reg_A[63]), .D(n25339), .Y(
        n32550) );
  OAI21X1 U26893 ( .A(n25038), .B(n30016), .C(n32551), .Y(n32548) );
  AOI22X1 U26894 ( .A(reg_A[60]), .B(n25246), .C(reg_A[59]), .D(n25247), .Y(
        n32551) );
  AOI21X1 U26895 ( .A(reg_A[49]), .B(n25253), .C(n32552), .Y(n32546) );
  OAI22X1 U26896 ( .A(n25040), .B(n30066), .C(n25041), .D(n30069), .Y(n32552)
         );
  AOI22X1 U26897 ( .A(reg_A[50]), .B(n25628), .C(reg_A[47]), .D(n25067), .Y(
        n32545) );
  AOI22X1 U26898 ( .A(n32131), .B(n32553), .C(n32482), .D(n32554), .Y(n32534)
         );
  INVX1 U26899 ( .A(n32333), .Y(n32482) );
  INVX1 U26900 ( .A(n32331), .Y(n32131) );
  NAND2X1 U26901 ( .A(reg_B[47]), .B(n25029), .Y(n32331) );
  OAI21X1 U26902 ( .A(n25087), .B(n32555), .C(n32556), .Y(n32532) );
  AOI22X1 U26903 ( .A(n32557), .B(n32312), .C(n32558), .D(n26504), .Y(n32556)
         );
  NOR2X1 U26904 ( .A(reg_B[47]), .B(n32480), .Y(n32558) );
  INVX1 U26905 ( .A(n32554), .Y(n32480) );
  OAI21X1 U26906 ( .A(n30463), .B(n32486), .C(n32466), .Y(n32554) );
  NAND2X1 U26907 ( .A(n32559), .B(reg_A[43]), .Y(n32466) );
  INVX1 U26908 ( .A(n32560), .Y(n32312) );
  OAI21X1 U26909 ( .A(n32146), .B(n32416), .C(n32561), .Y(n32560) );
  AOI21X1 U26910 ( .A(n32562), .B(n32233), .C(n32563), .Y(n32561) );
  INVX1 U26911 ( .A(n32145), .Y(n32562) );
  MUX2X1 U26912 ( .B(n32564), .A(n32565), .S(reg_B[47]), .Y(n32145) );
  INVX1 U26913 ( .A(n32566), .Y(n32565) );
  MUX2X1 U26914 ( .B(reg_A[43]), .A(reg_A[35]), .S(reg_B[44]), .Y(n32564) );
  NOR2X1 U26915 ( .A(reg_B[46]), .B(n25032), .Y(n32557) );
  NAND2X1 U26916 ( .A(n32567), .B(n32568), .Y(n32555) );
  AOI22X1 U26917 ( .A(n32569), .B(n30672), .C(reg_A[33]), .D(n28649), .Y(
        n32530) );
  NAND2X1 U26918 ( .A(n29973), .B(n30210), .Y(n30672) );
  AOI22X1 U26919 ( .A(reg_A[47]), .B(n28802), .C(n32570), .D(n32311), .Y(
        n32529) );
  INVX1 U26920 ( .A(n32571), .Y(n32311) );
  NOR2X1 U26921 ( .A(n32572), .B(n32573), .Y(n32507) );
  NAND3X1 U26922 ( .A(n32574), .B(n32575), .C(n32576), .Y(n32573) );
  NOR2X1 U26923 ( .A(n32577), .B(n32578), .Y(n32576) );
  OAI21X1 U26924 ( .A(n32240), .B(n32579), .C(n32490), .Y(n32578) );
  OAI22X1 U26925 ( .A(n28562), .B(n30058), .C(n32580), .D(n30524), .Y(n32577)
         );
  AOI22X1 U26926 ( .A(reg_A[43]), .B(n28661), .C(reg_A[42]), .D(n26626), .Y(
        n32575) );
  AOI22X1 U26927 ( .A(n32581), .B(n26756), .C(n32582), .D(n25119), .Y(n32574)
         );
  NAND3X1 U26928 ( .A(n32583), .B(n32584), .C(n32585), .Y(n32582) );
  NOR2X1 U26929 ( .A(n32586), .B(n32587), .Y(n32585) );
  OAI21X1 U26930 ( .A(n25056), .B(n30059), .C(n32588), .Y(n32587) );
  AOI22X1 U26931 ( .A(reg_A[37]), .B(n25253), .C(reg_A[36]), .D(n25628), .Y(
        n32588) );
  OAI21X1 U26932 ( .A(n25040), .B(n30463), .C(n32589), .Y(n32586) );
  AOI22X1 U26933 ( .A(reg_A[42]), .B(n25135), .C(reg_A[40]), .D(n25136), .Y(
        n32589) );
  AOI21X1 U26934 ( .A(reg_A[35]), .B(n25124), .C(n32590), .Y(n32584) );
  OAI22X1 U26935 ( .A(n25037), .B(n30394), .C(n26703), .D(n30060), .Y(n32590)
         );
  AOI22X1 U26936 ( .A(reg_A[33]), .B(n25637), .C(reg_A[43]), .D(n25125), .Y(
        n32583) );
  OAI21X1 U26937 ( .A(n32591), .B(n30038), .C(n32592), .Y(n32581) );
  AOI22X1 U26938 ( .A(n30846), .B(n32464), .C(n30212), .D(n32485), .Y(n32592)
         );
  INVX1 U26939 ( .A(n32353), .Y(n32464) );
  AOI22X1 U26940 ( .A(n31847), .B(n29973), .C(reg_A[39]), .D(n32420), .Y(
        n32353) );
  OAI22X1 U26941 ( .A(n30393), .B(n25045), .C(n29994), .D(n30160), .Y(n31847)
         );
  NAND3X1 U26942 ( .A(n32593), .B(n32594), .C(n32595), .Y(n32572) );
  NOR2X1 U26943 ( .A(n32596), .B(n32597), .Y(n32595) );
  OAI22X1 U26944 ( .A(n28570), .B(n30069), .C(n26854), .D(n32378), .Y(n32597)
         );
  OAI21X1 U26945 ( .A(reg_B[2]), .B(n32598), .C(n32599), .Y(n32378) );
  AOI22X1 U26946 ( .A(n26455), .B(n30395), .C(n26456), .D(n32600), .Y(n32599)
         );
  INVX1 U26947 ( .A(n32033), .Y(n32600) );
  INVX1 U26948 ( .A(n32035), .Y(n32598) );
  OAI21X1 U26949 ( .A(reg_B[4]), .B(n31888), .C(n32601), .Y(n32035) );
  AOI22X1 U26950 ( .A(n26462), .B(n30462), .C(n26463), .D(n30394), .Y(n32601)
         );
  MUX2X1 U26951 ( .B(n30160), .A(n30393), .S(reg_B[1]), .Y(n31888) );
  OAI21X1 U26952 ( .A(n28571), .B(n30060), .C(n32602), .Y(n32596) );
  AOI22X1 U26953 ( .A(reg_A[39]), .B(n25181), .C(reg_A[35]), .D(n28717), .Y(
        n32602) );
  AOI22X1 U26954 ( .A(reg_A[45]), .B(n25153), .C(reg_A[44]), .D(n28280), .Y(
        n32594) );
  AOI22X1 U26955 ( .A(reg_A[40]), .B(n32603), .C(n32604), .D(n26262), .Y(
        n32593) );
  NAND2X1 U26956 ( .A(n32605), .B(n32606), .Y(result[42]) );
  NOR2X1 U26957 ( .A(n32607), .B(n32608), .Y(n32606) );
  NAND3X1 U26958 ( .A(n32609), .B(n32610), .C(n32611), .Y(n32608) );
  NOR2X1 U26959 ( .A(n32612), .B(n32613), .Y(n32611) );
  OAI21X1 U26960 ( .A(n32516), .B(n30038), .C(n32614), .Y(n32613) );
  OAI21X1 U26961 ( .A(n32615), .B(n32616), .C(n26267), .Y(n32614) );
  OAI22X1 U26962 ( .A(n32521), .B(n32066), .C(n32413), .D(n32134), .Y(n32616)
         );
  INVX1 U26963 ( .A(n32617), .Y(n32413) );
  OAI21X1 U26964 ( .A(n30462), .B(n32371), .C(n32618), .Y(n32617) );
  AOI22X1 U26965 ( .A(n32147), .B(reg_A[34]), .C(n32260), .D(reg_A[38]), .Y(
        n32618) );
  NOR2X1 U26966 ( .A(n32619), .B(n32240), .Y(n32615) );
  INVX1 U26967 ( .A(n32620), .Y(n32516) );
  OAI21X1 U26968 ( .A(n30744), .B(n32621), .C(n32622), .Y(n32620) );
  NAND2X1 U26969 ( .A(n30298), .B(n25932), .Y(n32621) );
  OAI21X1 U26970 ( .A(n28592), .B(n30069), .C(n32623), .Y(n32612) );
  OAI21X1 U26971 ( .A(n32624), .B(n32625), .C(n26480), .Y(n32623) );
  OAI22X1 U26972 ( .A(n32245), .B(n32041), .C(n32246), .D(n32043), .Y(n32625)
         );
  OAI21X1 U26973 ( .A(n32626), .B(n32045), .C(n32627), .Y(n32624) );
  AOI22X1 U26974 ( .A(n32628), .B(n32248), .C(n30340), .D(n32249), .Y(n32627)
         );
  AOI22X1 U26975 ( .A(n32206), .B(n32233), .C(reg_A[40]), .D(n28772), .Y(
        n32610) );
  OAI22X1 U26976 ( .A(n32629), .B(n32630), .C(n25031), .D(n32631), .Y(n32206)
         );
  OAI21X1 U26977 ( .A(n32632), .B(n32253), .C(n25188), .Y(n32630) );
  OAI21X1 U26978 ( .A(n32566), .B(n32134), .C(n32633), .Y(n32629) );
  AOI22X1 U26979 ( .A(n32634), .B(n32635), .C(n32636), .D(reg_B[46]), .Y(
        n32633) );
  INVX1 U26980 ( .A(n32637), .Y(n32636) );
  OAI22X1 U26981 ( .A(reg_A[39]), .B(n32240), .C(reg_A[40]), .D(n32066), .Y(
        n32634) );
  MUX2X1 U26982 ( .B(n30462), .A(n30394), .S(reg_B[44]), .Y(n32566) );
  AOI22X1 U26983 ( .A(n32109), .B(n32638), .C(reg_A[33]), .D(n28572), .Y(
        n32609) );
  NAND3X1 U26984 ( .A(n32639), .B(n32640), .C(n32641), .Y(n32607) );
  NOR2X1 U26985 ( .A(n32642), .B(n32643), .Y(n32641) );
  OAI21X1 U26986 ( .A(n32644), .B(n25794), .C(n32645), .Y(n32643) );
  OAI21X1 U26987 ( .A(n32646), .B(n32647), .C(n25310), .Y(n32645) );
  NAND3X1 U26988 ( .A(n32648), .B(n32649), .C(n32650), .Y(n32647) );
  NOR2X1 U26989 ( .A(n32651), .B(n32652), .Y(n32650) );
  OAI21X1 U26990 ( .A(n25036), .B(n30378), .C(n32653), .Y(n32652) );
  AOI22X1 U26991 ( .A(reg_A[50]), .B(n25124), .C(reg_A[53]), .D(n25222), .Y(
        n32653) );
  OAI21X1 U26992 ( .A(n25037), .B(n30009), .C(n32654), .Y(n32651) );
  AOI22X1 U26993 ( .A(reg_A[46]), .B(n25072), .C(reg_A[47]), .D(n25123), .Y(
        n32654) );
  AOI21X1 U26994 ( .A(reg_A[54]), .B(n25635), .C(n32655), .Y(n32649) );
  OAI22X1 U26995 ( .A(n25065), .B(n29990), .C(n25475), .D(n30254), .Y(n32655)
         );
  AOI22X1 U26996 ( .A(reg_A[55]), .B(n25325), .C(reg_A[42]), .D(n25125), .Y(
        n32648) );
  NAND3X1 U26997 ( .A(n32656), .B(n32657), .C(n32658), .Y(n32646) );
  NOR2X1 U26998 ( .A(n32659), .B(n32660), .Y(n32658) );
  OAI21X1 U26999 ( .A(n26719), .B(n30007), .C(n32661), .Y(n32660) );
  AOI22X1 U27000 ( .A(reg_A[60]), .B(n25241), .C(reg_A[62]), .D(n25339), .Y(
        n32661) );
  OAI21X1 U27001 ( .A(n25038), .B(n29989), .C(n32662), .Y(n32659) );
  AOI22X1 U27002 ( .A(reg_A[59]), .B(n25246), .C(reg_A[58]), .D(n25247), .Y(
        n32662) );
  AOI21X1 U27003 ( .A(reg_A[44]), .B(n25252), .C(n32663), .Y(n32657) );
  OAI22X1 U27004 ( .A(n25041), .B(n30066), .C(n25042), .D(n30160), .Y(n32663)
         );
  AOI22X1 U27005 ( .A(reg_A[48]), .B(n25253), .C(reg_A[49]), .D(n25628), .Y(
        n32656) );
  AOI21X1 U27006 ( .A(n32227), .B(n32260), .C(n32664), .Y(n32644) );
  INVX1 U27007 ( .A(n32417), .Y(n32664) );
  NAND2X1 U27008 ( .A(n32665), .B(reg_B[45]), .Y(n32417) );
  AND2X1 U27009 ( .A(n32666), .B(n32667), .Y(n32227) );
  AOI22X1 U27010 ( .A(n32299), .B(n30058), .C(n32109), .D(n30057), .Y(n32667)
         );
  AOI22X1 U27011 ( .A(n32357), .B(n30393), .C(n32110), .D(n30060), .Y(n32666)
         );
  OAI21X1 U27012 ( .A(n32333), .B(n32668), .C(n32669), .Y(n32642) );
  AOI21X1 U27013 ( .A(n32670), .B(n32128), .C(n31645), .Y(n32669) );
  INVX1 U27014 ( .A(n32671), .Y(n32128) );
  NOR2X1 U27015 ( .A(n32672), .B(n25087), .Y(n32670) );
  NAND2X1 U27016 ( .A(n25170), .B(n32553), .Y(n32668) );
  OAI22X1 U27017 ( .A(n30744), .B(n32486), .C(n30462), .D(n32049), .Y(n32553)
         );
  NAND2X1 U27018 ( .A(reg_B[46]), .B(n32233), .Y(n32486) );
  NAND2X1 U27019 ( .A(n25029), .B(n32229), .Y(n32333) );
  AOI22X1 U27020 ( .A(n32266), .B(n28735), .C(n32267), .D(n32673), .Y(n32640)
         );
  INVX1 U27021 ( .A(n32316), .Y(n32267) );
  NAND2X1 U27022 ( .A(n32674), .B(n25382), .Y(n32316) );
  NOR2X1 U27023 ( .A(n32675), .B(n32676), .Y(n32266) );
  OAI22X1 U27024 ( .A(n32677), .B(n27454), .C(n31942), .D(n26599), .Y(n32676)
         );
  MUX2X1 U27025 ( .B(n30462), .A(n30394), .S(reg_B[1]), .Y(n31942) );
  OAI21X1 U27026 ( .A(reg_A[32]), .B(n28739), .C(n32678), .Y(n32675) );
  AOI22X1 U27027 ( .A(n28741), .B(n30059), .C(n28742), .D(n30744), .Y(n32678)
         );
  AOI22X1 U27028 ( .A(reg_A[47]), .B(n28726), .C(n32569), .D(n30223), .Y(
        n32639) );
  NOR2X1 U27029 ( .A(n32679), .B(n32680), .Y(n32605) );
  NAND3X1 U27030 ( .A(n32681), .B(n32682), .C(n32683), .Y(n32680) );
  NOR2X1 U27031 ( .A(n32684), .B(n32685), .Y(n32683) );
  OAI22X1 U27032 ( .A(n32559), .B(n32579), .C(n28562), .D(n30393), .Y(n32685)
         );
  INVX1 U27033 ( .A(n32049), .Y(n32559) );
  NAND2X1 U27034 ( .A(n32233), .B(n32334), .Y(n32049) );
  OAI21X1 U27035 ( .A(n32686), .B(n30524), .C(n32687), .Y(n32684) );
  OAI21X1 U27036 ( .A(n32688), .B(n32689), .C(n25119), .Y(n32687) );
  OR2X1 U27037 ( .A(n32690), .B(n32691), .Y(n32689) );
  OAI22X1 U27038 ( .A(n25043), .B(n30462), .C(n25467), .D(n30394), .Y(n32691)
         );
  OAI21X1 U27039 ( .A(n25037), .B(n30170), .C(n32692), .Y(n32690) );
  AOI22X1 U27040 ( .A(reg_A[38]), .B(n25073), .C(reg_A[37]), .D(n25123), .Y(
        n32692) );
  OR2X1 U27041 ( .A(n32693), .B(n32694), .Y(n32688) );
  OAI22X1 U27042 ( .A(n25030), .B(n30393), .C(n25033), .D(n30058), .Y(n32694)
         );
  OAI21X1 U27043 ( .A(n25040), .B(n30744), .C(n32695), .Y(n32693) );
  AOI22X1 U27044 ( .A(reg_A[41]), .B(n25135), .C(reg_A[39]), .D(n25136), .Y(
        n32695) );
  AOI22X1 U27045 ( .A(reg_A[32]), .B(n28700), .C(reg_A[42]), .D(n28661), .Y(
        n32682) );
  AOI22X1 U27046 ( .A(reg_A[41]), .B(n26626), .C(n32696), .D(n26756), .Y(
        n32681) );
  OAI21X1 U27047 ( .A(n32697), .B(n30210), .C(n32698), .Y(n32696) );
  AOI22X1 U27048 ( .A(n30846), .B(n32485), .C(n30212), .D(n32465), .Y(n32698)
         );
  OAI22X1 U27049 ( .A(n32059), .B(reg_B[61]), .C(n30060), .D(n32045), .Y(
        n32485) );
  INVX1 U27050 ( .A(n32008), .Y(n32059) );
  OAI22X1 U27051 ( .A(n30394), .B(n30109), .C(n29994), .D(n30462), .Y(n32008)
         );
  NAND3X1 U27052 ( .A(n32699), .B(n32700), .C(n32701), .Y(n32679) );
  NOR2X1 U27053 ( .A(n32702), .B(n32703), .Y(n32701) );
  OAI22X1 U27054 ( .A(n25178), .B(n30394), .C(n28679), .D(n30060), .Y(n32703)
         );
  OAI21X1 U27055 ( .A(n28714), .B(n30058), .C(n32704), .Y(n32702) );
  AOI22X1 U27056 ( .A(n32207), .B(n28575), .C(reg_A[39]), .D(n25180), .Y(
        n32704) );
  AOI22X1 U27057 ( .A(reg_A[37]), .B(n25149), .C(reg_A[45]), .D(n25152), .Y(
        n32700) );
  AOI22X1 U27058 ( .A(reg_A[44]), .B(n25153), .C(reg_A[43]), .D(n28280), .Y(
        n32699) );
  NAND3X1 U27059 ( .A(n32705), .B(n32706), .C(n32707), .Y(result[41]) );
  NOR2X1 U27060 ( .A(n32708), .B(n32709), .Y(n32707) );
  NAND3X1 U27061 ( .A(n32710), .B(n32711), .C(n32712), .Y(n32709) );
  NOR2X1 U27062 ( .A(n32713), .B(n32714), .Y(n32712) );
  OAI21X1 U27063 ( .A(n32715), .B(n25087), .C(n32490), .Y(n32714) );
  NOR2X1 U27064 ( .A(n31645), .B(n32205), .Y(n32490) );
  NOR2X1 U27065 ( .A(n32579), .B(n32233), .Y(n32205) );
  INVX1 U27066 ( .A(n31954), .Y(n31645) );
  NAND2X1 U27067 ( .A(n31689), .B(n25932), .Y(n31954) );
  INVX1 U27068 ( .A(n31693), .Y(n31689) );
  NAND2X1 U27069 ( .A(reg_B[59]), .B(reg_A[32]), .Y(n31693) );
  AOI21X1 U27070 ( .A(n32674), .B(n32716), .C(n32717), .Y(n32715) );
  OAI21X1 U27071 ( .A(n32315), .B(n32671), .C(n32718), .Y(n32717) );
  OAI21X1 U27072 ( .A(n32719), .B(n32720), .C(n25044), .Y(n32718) );
  OAI21X1 U27073 ( .A(n32721), .B(n29976), .C(n32722), .Y(n32720) );
  AOI22X1 U27074 ( .A(n30039), .B(n32723), .C(n32724), .D(n32725), .Y(n32722)
         );
  OAI21X1 U27075 ( .A(n32726), .B(n32045), .C(n32727), .Y(n32719) );
  AOI22X1 U27076 ( .A(n32628), .B(n30285), .C(n30340), .D(n32310), .Y(n32727)
         );
  INVX1 U27077 ( .A(n32137), .Y(n32674) );
  MUX2X1 U27078 ( .B(n32728), .A(n32579), .S(n32134), .Y(n32713) );
  NAND2X1 U27079 ( .A(reg_A[40]), .B(n26504), .Y(n32579) );
  INVX1 U27080 ( .A(n32638), .Y(n32728) );
  OAI21X1 U27081 ( .A(n32412), .B(n26147), .C(n32729), .Y(n32638) );
  OAI21X1 U27082 ( .A(n32730), .B(n32731), .C(reg_A[41]), .Y(n32729) );
  INVX1 U27083 ( .A(n32322), .Y(n32731) );
  NAND2X1 U27084 ( .A(n26504), .B(n32233), .Y(n32322) );
  NOR2X1 U27085 ( .A(reg_B[45]), .B(n26151), .Y(n32730) );
  INVX1 U27086 ( .A(n32732), .Y(n32412) );
  OAI21X1 U27087 ( .A(n30463), .B(n32371), .C(n32733), .Y(n32732) );
  AOI22X1 U27088 ( .A(n32147), .B(reg_A[33]), .C(n32260), .D(reg_A[37]), .Y(
        n32733) );
  OAI21X1 U27089 ( .A(n32734), .B(n32735), .C(n25119), .Y(n32711) );
  NAND2X1 U27090 ( .A(n32736), .B(n32737), .Y(n32735) );
  AOI22X1 U27091 ( .A(reg_A[37]), .B(n25073), .C(reg_A[36]), .D(n25123), .Y(
        n32737) );
  AOI22X1 U27092 ( .A(reg_A[33]), .B(n25124), .C(reg_A[41]), .D(n25125), .Y(
        n32736) );
  OR2X1 U27093 ( .A(n32738), .B(n32739), .Y(n32734) );
  OAI22X1 U27094 ( .A(n25030), .B(n30394), .C(n25033), .D(n30393), .Y(n32739)
         );
  OAI21X1 U27095 ( .A(n25040), .B(n30059), .C(n32740), .Y(n32738) );
  AOI22X1 U27096 ( .A(reg_A[40]), .B(n25135), .C(reg_A[38]), .D(n25136), .Y(
        n32740) );
  AOI22X1 U27097 ( .A(reg_A[32]), .B(n25137), .C(reg_A[39]), .D(n25138), .Y(
        n32710) );
  OR2X1 U27098 ( .A(n32741), .B(n28572), .Y(n25137) );
  NAND3X1 U27099 ( .A(n32742), .B(n32743), .C(n32744), .Y(n32708) );
  AOI21X1 U27100 ( .A(n30212), .B(n32745), .C(n32746), .Y(n32744) );
  OAI22X1 U27101 ( .A(n25145), .B(n30463), .C(n25148), .D(n30462), .Y(n32746)
         );
  AOI22X1 U27102 ( .A(reg_A[36]), .B(n25149), .C(n32604), .D(n25150), .Y(
        n32743) );
  AND2X1 U27103 ( .A(n32747), .B(n32748), .Y(n32604) );
  AOI22X1 U27104 ( .A(n26859), .B(n30058), .C(n26860), .D(n30057), .Y(n32748)
         );
  AOI22X1 U27105 ( .A(n26455), .B(n30395), .C(n32361), .D(n26452), .Y(n32747)
         );
  OAI21X1 U27106 ( .A(reg_A[32]), .B(n26861), .C(n32749), .Y(n32361) );
  AOI22X1 U27107 ( .A(n32750), .B(n26863), .C(n26462), .D(n30744), .Y(n32749)
         );
  INVX1 U27108 ( .A(n32677), .Y(n32750) );
  MUX2X1 U27109 ( .B(n30463), .A(n30170), .S(reg_B[1]), .Y(n32677) );
  AOI22X1 U27110 ( .A(reg_A[44]), .B(n25152), .C(reg_A[43]), .D(n25153), .Y(
        n32742) );
  NOR2X1 U27111 ( .A(n32751), .B(n32752), .Y(n32706) );
  OAI21X1 U27112 ( .A(n25162), .B(n30393), .C(n32753), .Y(n32752) );
  AOI22X1 U27113 ( .A(n32569), .B(n30103), .C(n32033), .D(n25166), .Y(n32753)
         );
  NAND2X1 U27114 ( .A(n26878), .B(n27067), .Y(n25162) );
  NAND2X1 U27115 ( .A(n32754), .B(n32755), .Y(n32751) );
  AOI22X1 U27116 ( .A(n32756), .B(n32109), .C(n26267), .D(n32757), .Y(n32755)
         );
  OAI22X1 U27117 ( .A(n32758), .B(n32240), .C(n32619), .D(n32066), .Y(n32757)
         );
  AND2X1 U27118 ( .A(n32759), .B(n25170), .Y(n32756) );
  AOI22X1 U27119 ( .A(reg_A[40]), .B(n32760), .C(n32761), .D(n26756), .Y(
        n32754) );
  OAI21X1 U27120 ( .A(n32762), .B(n30210), .C(n32763), .Y(n32761) );
  AOI22X1 U27121 ( .A(n30846), .B(n32465), .C(n29987), .D(n32764), .Y(n32763)
         );
  INVX1 U27122 ( .A(n32591), .Y(n32465) );
  AOI22X1 U27123 ( .A(n31955), .B(n29973), .C(reg_A[37]), .D(n32420), .Y(
        n32591) );
  OAI22X1 U27124 ( .A(n30170), .B(n30109), .C(n29994), .D(n30463), .Y(n31955)
         );
  OAI21X1 U27125 ( .A(n27438), .B(n32765), .C(n28870), .Y(n32760) );
  NOR2X1 U27126 ( .A(n32766), .B(n32767), .Y(n32705) );
  OAI21X1 U27127 ( .A(n25178), .B(n30170), .C(n32768), .Y(n32767) );
  AOI22X1 U27128 ( .A(reg_A[38]), .B(n25180), .C(reg_A[37]), .D(n25181), .Y(
        n32768) );
  OAI21X1 U27129 ( .A(n25184), .B(n30394), .C(n32769), .Y(n32766) );
  AND2X1 U27130 ( .A(n32770), .B(n32771), .Y(n32769) );
  OAI21X1 U27131 ( .A(n32772), .B(n32773), .C(n25203), .Y(n32771) );
  OAI22X1 U27132 ( .A(n25204), .B(n30463), .C(n25205), .D(n30066), .Y(n32773)
         );
  OAI21X1 U27133 ( .A(n25207), .B(n30069), .C(n32774), .Y(n32772) );
  AOI22X1 U27134 ( .A(n25097), .B(n32775), .C(reg_A[47]), .D(n25211), .Y(
        n32774) );
  NAND3X1 U27135 ( .A(n32776), .B(n32777), .C(n32778), .Y(n32775) );
  AND2X1 U27136 ( .A(n32779), .B(n32780), .Y(n32778) );
  NOR2X1 U27137 ( .A(n32781), .B(n32782), .Y(n32780) );
  OAI21X1 U27138 ( .A(n25036), .B(n30009), .C(n32783), .Y(n32782) );
  AOI22X1 U27139 ( .A(reg_A[49]), .B(n25124), .C(reg_A[52]), .D(n25222), .Y(
        n32783) );
  OAI21X1 U27140 ( .A(n25037), .B(n30008), .C(n32784), .Y(n32781) );
  AOI22X1 U27141 ( .A(reg_A[45]), .B(n25073), .C(reg_A[46]), .D(n25123), .Y(
        n32784) );
  NOR2X1 U27142 ( .A(n32785), .B(n32786), .Y(n32779) );
  OAI22X1 U27143 ( .A(n25043), .B(n30463), .C(n25039), .D(n30168), .Y(n32786)
         );
  OAI21X1 U27144 ( .A(n25064), .B(n30299), .C(n32787), .Y(n32785) );
  AOI22X1 U27145 ( .A(reg_A[55]), .B(n25234), .C(reg_A[56]), .D(n25235), .Y(
        n32787) );
  NOR2X1 U27146 ( .A(n32788), .B(n32789), .Y(n32777) );
  OAI21X1 U27147 ( .A(n25238), .B(n29989), .C(n32790), .Y(n32789) );
  AOI22X1 U27148 ( .A(reg_A[59]), .B(n25241), .C(reg_A[63]), .D(n25242), .Y(
        n32790) );
  OAI21X1 U27149 ( .A(n25038), .B(n30015), .C(n32791), .Y(n32788) );
  AOI22X1 U27150 ( .A(reg_A[58]), .B(n25246), .C(reg_A[57]), .D(n25247), .Y(
        n32791) );
  NOR2X1 U27151 ( .A(n32792), .B(n32793), .Y(n32776) );
  OAI21X1 U27152 ( .A(n25030), .B(n29655), .C(n32794), .Y(n32793) );
  AOI22X1 U27153 ( .A(reg_A[43]), .B(n25252), .C(reg_A[47]), .D(n25253), .Y(
        n32794) );
  OAI21X1 U27154 ( .A(n25041), .B(n30067), .C(n32795), .Y(n32792) );
  AOI22X1 U27155 ( .A(reg_A[62]), .B(n25257), .C(reg_A[42]), .D(n25135), .Y(
        n32795) );
  OAI21X1 U27156 ( .A(n32796), .B(n32797), .C(n25188), .Y(n32770) );
  OAI21X1 U27157 ( .A(n32066), .B(n32798), .C(n32799), .Y(n32797) );
  MUX2X1 U27158 ( .B(n32570), .A(n32665), .S(reg_B[46]), .Y(n32799) );
  INVX1 U27159 ( .A(n32800), .Y(n32570) );
  OAI21X1 U27160 ( .A(reg_B[45]), .B(n32369), .C(n32801), .Y(n32800) );
  AOI21X1 U27161 ( .A(n32260), .B(n32802), .C(n32563), .Y(n32801) );
  NOR2X1 U27162 ( .A(n32637), .B(n32233), .Y(n32563) );
  INVX1 U27163 ( .A(n32370), .Y(n32802) );
  MUX2X1 U27164 ( .B(n30057), .A(n30058), .S(reg_B[47]), .Y(n32370) );
  MUX2X1 U27165 ( .B(n32803), .A(n32804), .S(reg_B[47]), .Y(n32369) );
  OAI21X1 U27166 ( .A(reg_B[44]), .B(reg_A[40]), .C(n32637), .Y(n32804) );
  NAND2X1 U27167 ( .A(reg_B[44]), .B(n30395), .Y(n32637) );
  INVX1 U27168 ( .A(n32632), .Y(n32803) );
  MUX2X1 U27169 ( .B(n30463), .A(n30170), .S(reg_B[44]), .Y(n32632) );
  OAI22X1 U27170 ( .A(n32240), .B(n32805), .C(n32806), .D(n32807), .Y(n32796)
         );
  INVX1 U27171 ( .A(n32146), .Y(n32806) );
  MUX2X1 U27172 ( .B(n30059), .A(n30060), .S(reg_B[47]), .Y(n32146) );
  AOI21X1 U27173 ( .A(n30910), .B(n25613), .C(n32498), .Y(n25184) );
  NAND3X1 U27174 ( .A(n32808), .B(n32809), .C(n32810), .Y(result[40]) );
  NOR2X1 U27175 ( .A(n32811), .B(n32812), .Y(n32810) );
  NAND3X1 U27176 ( .A(n32813), .B(n32814), .C(n32815), .Y(n32812) );
  AOI21X1 U27177 ( .A(reg_A[33]), .B(n26673), .C(n32816), .Y(n32815) );
  OAI22X1 U27178 ( .A(n26675), .B(n30067), .C(n26676), .D(n30060), .Y(n32816)
         );
  INVX1 U27179 ( .A(n28942), .Y(n26676) );
  OAI21X1 U27180 ( .A(n28516), .B(n25133), .C(n32817), .Y(n28942) );
  INVX1 U27181 ( .A(n28943), .Y(n26675) );
  OAI21X1 U27182 ( .A(n26801), .B(n27152), .C(n32818), .Y(n28943) );
  OAI21X1 U27183 ( .A(n28516), .B(n25129), .C(n28562), .Y(n26673) );
  AOI22X1 U27184 ( .A(reg_A[34]), .B(n26678), .C(reg_A[35]), .D(n26679), .Y(
        n32814) );
  OAI21X1 U27185 ( .A(n28516), .B(n26703), .C(n28571), .Y(n26679) );
  OAI21X1 U27186 ( .A(n28516), .B(n25131), .C(n28714), .Y(n26678) );
  AOI22X1 U27187 ( .A(reg_A[36]), .B(n26680), .C(reg_A[37]), .D(n26681), .Y(
        n32813) );
  OAI21X1 U27188 ( .A(n28516), .B(n25254), .C(n28715), .Y(n26681) );
  OAI21X1 U27189 ( .A(n28516), .B(n26431), .C(n28679), .Y(n26680) );
  NAND2X1 U27190 ( .A(n32819), .B(n32820), .Y(n32811) );
  NOR2X1 U27191 ( .A(n32821), .B(n32822), .Y(n32820) );
  OAI21X1 U27192 ( .A(n32134), .B(n32823), .C(n32824), .Y(n32822) );
  OAI21X1 U27193 ( .A(n32825), .B(n26690), .C(reg_A[40]), .Y(n32824) );
  NAND3X1 U27194 ( .A(n32826), .B(n32827), .C(n32828), .Y(n26690) );
  AOI21X1 U27195 ( .A(n25125), .B(n25119), .C(n32829), .Y(n32828) );
  NAND2X1 U27196 ( .A(n25170), .B(n32759), .Y(n32823) );
  OAI21X1 U27197 ( .A(n32521), .B(n25415), .C(n32830), .Y(n32759) );
  NAND3X1 U27198 ( .A(n25589), .B(n32233), .C(reg_A[40]), .Y(n32830) );
  INVX1 U27199 ( .A(n32831), .Y(n32521) );
  OAI21X1 U27200 ( .A(n30744), .B(n32371), .C(n32832), .Y(n32831) );
  AOI22X1 U27201 ( .A(n32665), .B(n32233), .C(n32260), .D(reg_A[36]), .Y(
        n32832) );
  OAI21X1 U27202 ( .A(n32439), .B(n32833), .C(n32834), .Y(n32821) );
  OAI21X1 U27203 ( .A(n32835), .B(n32836), .C(n25310), .Y(n32834) );
  NAND2X1 U27204 ( .A(n32837), .B(n32838), .Y(n32836) );
  NOR2X1 U27205 ( .A(n32839), .B(n32840), .Y(n32838) );
  OAI21X1 U27206 ( .A(n25043), .B(n30744), .C(n32841), .Y(n32840) );
  AOI22X1 U27207 ( .A(reg_A[41]), .B(n25135), .C(reg_A[42]), .D(n25252), .Y(
        n32841) );
  OAI21X1 U27208 ( .A(n25028), .B(n30066), .C(n32842), .Y(n32839) );
  AOI22X1 U27209 ( .A(reg_A[43]), .B(n25136), .C(reg_A[44]), .D(n25066), .Y(
        n32842) );
  NOR2X1 U27210 ( .A(n32843), .B(n32844), .Y(n32837) );
  OAI21X1 U27211 ( .A(n25034), .B(n29655), .C(n32845), .Y(n32844) );
  AOI22X1 U27212 ( .A(reg_A[46]), .B(n25253), .C(reg_A[47]), .D(n25628), .Y(
        n32845) );
  OAI21X1 U27213 ( .A(n25036), .B(n30008), .C(n32846), .Y(n32843) );
  AOI22X1 U27214 ( .A(reg_A[49]), .B(n25629), .C(reg_A[51]), .D(n25222), .Y(
        n32846) );
  NAND2X1 U27215 ( .A(n32847), .B(n32848), .Y(n32835) );
  NOR2X1 U27216 ( .A(n32849), .B(n32850), .Y(n32848) );
  OAI21X1 U27217 ( .A(n25039), .B(n30299), .C(n32851), .Y(n32850) );
  AOI22X1 U27218 ( .A(reg_A[54]), .B(n25234), .C(reg_A[52]), .D(n25635), .Y(
        n32851) );
  OAI21X1 U27219 ( .A(n25065), .B(n30043), .C(n32852), .Y(n32849) );
  AOI22X1 U27220 ( .A(reg_A[57]), .B(n25246), .C(reg_A[56]), .D(n25247), .Y(
        n32852) );
  NOR2X1 U27221 ( .A(n32853), .B(n32854), .Y(n32847) );
  OAI21X1 U27222 ( .A(n25238), .B(n30015), .C(n32855), .Y(n32854) );
  AOI22X1 U27223 ( .A(reg_A[59]), .B(n25487), .C(reg_A[58]), .D(n25241), .Y(
        n32855) );
  OAI21X1 U27224 ( .A(n26719), .B(n29989), .C(n32856), .Y(n32853) );
  AOI22X1 U27225 ( .A(reg_A[62]), .B(n25242), .C(reg_A[63]), .D(n25338), .Y(
        n32856) );
  NAND2X1 U27226 ( .A(n32260), .B(n25188), .Y(n32833) );
  NAND2X1 U27227 ( .A(n32857), .B(n32858), .Y(n32439) );
  AOI22X1 U27228 ( .A(n32299), .B(n30394), .C(n32109), .D(n30393), .Y(n32858)
         );
  AOI22X1 U27229 ( .A(n32357), .B(n30170), .C(n32110), .D(n30058), .Y(n32857)
         );
  AOI21X1 U27230 ( .A(n26267), .B(n32859), .C(n32860), .Y(n32819) );
  OAI22X1 U27231 ( .A(n32283), .B(n32438), .C(n26729), .D(n32506), .Y(n32860)
         );
  NAND2X1 U27232 ( .A(n32861), .B(n32862), .Y(n32506) );
  AOI22X1 U27233 ( .A(n26601), .B(n30060), .C(n26602), .D(n30057), .Y(n32862)
         );
  AOI22X1 U27234 ( .A(n27012), .B(n30744), .C(n26597), .D(n30059), .Y(n32861)
         );
  NAND2X1 U27235 ( .A(n32863), .B(n32864), .Y(n32438) );
  AOI22X1 U27236 ( .A(n32299), .B(n30060), .C(n32109), .D(n30059), .Y(n32864)
         );
  AOI22X1 U27237 ( .A(n32357), .B(n30057), .C(n32110), .D(n30744), .Y(n32863)
         );
  OAI21X1 U27238 ( .A(n32865), .B(n32240), .C(n32866), .Y(n32859) );
  AOI22X1 U27239 ( .A(n32109), .B(n32867), .C(n32299), .D(n32868), .Y(n32866)
         );
  NOR2X1 U27240 ( .A(n32869), .B(n32870), .Y(n32809) );
  OAI21X1 U27241 ( .A(n32622), .B(n29970), .C(n32871), .Y(n32870) );
  AOI22X1 U27242 ( .A(n32504), .B(n28575), .C(reg_A[32]), .D(n28958), .Y(
        n32871) );
  NAND2X1 U27243 ( .A(n32872), .B(n25178), .Y(n28958) );
  INVX1 U27244 ( .A(n32745), .Y(n32622) );
  OAI21X1 U27245 ( .A(n27438), .B(n32873), .C(n32874), .Y(n32745) );
  OAI21X1 U27246 ( .A(n32875), .B(n32876), .C(n25699), .Y(n32874) );
  INVX1 U27247 ( .A(n32873), .Y(n32876) );
  AND2X1 U27248 ( .A(n29973), .B(n32198), .Y(n32875) );
  OAI22X1 U27249 ( .A(n30395), .B(n30109), .C(n29994), .D(n30744), .Y(n32198)
         );
  NAND2X1 U27250 ( .A(n32420), .B(reg_A[36]), .Y(n32873) );
  NAND2X1 U27251 ( .A(n32877), .B(n32878), .Y(n32869) );
  AOI22X1 U27252 ( .A(reg_A[45]), .B(n26746), .C(reg_A[46]), .D(n26747), .Y(
        n32878) );
  OAI22X1 U27253 ( .A(n25061), .B(n27152), .C(n25754), .D(n25726), .Y(n26747)
         );
  OAI22X1 U27254 ( .A(n26800), .B(n27152), .C(n26944), .D(n25726), .Y(n26746)
         );
  AOI22X1 U27255 ( .A(reg_A[47]), .B(n26748), .C(reg_A[39]), .D(n26749), .Y(
        n32877) );
  OAI21X1 U27256 ( .A(n28516), .B(n25784), .C(n32879), .Y(n26749) );
  INVX1 U27257 ( .A(n32880), .Y(n32879) );
  OAI22X1 U27258 ( .A(n26936), .B(n27152), .C(n25753), .D(n25726), .Y(n26748)
         );
  NOR2X1 U27259 ( .A(n32881), .B(n32882), .Y(n32808) );
  NAND3X1 U27260 ( .A(n32883), .B(n32884), .C(n32885), .Y(n32882) );
  NAND2X1 U27261 ( .A(n32886), .B(n26756), .Y(n32884) );
  OAI21X1 U27262 ( .A(n32887), .B(n30210), .C(n32888), .Y(n32886) );
  AOI22X1 U27263 ( .A(n30212), .B(n32764), .C(n29987), .D(n32889), .Y(n32888)
         );
  OAI21X1 U27264 ( .A(n32890), .B(n32891), .C(n25382), .Y(n32883) );
  OAI21X1 U27265 ( .A(n32892), .B(n32671), .C(n32893), .Y(n32891) );
  OAI21X1 U27266 ( .A(n32894), .B(n32895), .C(n25044), .Y(n32893) );
  OAI21X1 U27267 ( .A(n32428), .B(n32043), .C(n32896), .Y(n32895) );
  AOI22X1 U27268 ( .A(n32420), .B(n32497), .C(n32724), .D(n32427), .Y(n32896)
         );
  OAI21X1 U27269 ( .A(n32897), .B(n29976), .C(n32898), .Y(n32894) );
  AOI22X1 U27270 ( .A(n32628), .B(n31044), .C(n30340), .D(n31032), .Y(n32898)
         );
  INVX1 U27271 ( .A(n32247), .Y(n30340) );
  NAND2X1 U27272 ( .A(reg_B[59]), .B(n30325), .Y(n32247) );
  NOR2X1 U27273 ( .A(n30220), .B(n30341), .Y(n32628) );
  NAND2X1 U27274 ( .A(reg_B[45]), .B(n32568), .Y(n32671) );
  NOR2X1 U27275 ( .A(n32899), .B(n32137), .Y(n32890) );
  NAND2X1 U27276 ( .A(n32233), .B(n32568), .Y(n32137) );
  OAI21X1 U27277 ( .A(reg_B[44]), .B(n25415), .C(n26999), .Y(n32568) );
  OAI21X1 U27278 ( .A(n26781), .B(n30463), .C(n32900), .Y(n32881) );
  AOI22X1 U27279 ( .A(reg_A[43]), .B(n26739), .C(reg_A[42]), .D(n26783), .Y(
        n32900) );
  NAND3X1 U27280 ( .A(n32901), .B(n32902), .C(n32903), .Y(result[3]) );
  NOR2X1 U27281 ( .A(n32904), .B(n32905), .Y(n32903) );
  NAND2X1 U27282 ( .A(n32906), .B(n32907), .Y(n32905) );
  AOI21X1 U27283 ( .A(reg_A[15]), .B(n25363), .C(n32908), .Y(n32907) );
  OAI21X1 U27284 ( .A(n32909), .B(n25132), .C(n32910), .Y(n32908) );
  OAI21X1 U27285 ( .A(n32911), .B(n32912), .C(n25310), .Y(n32910) );
  NAND3X1 U27286 ( .A(n32913), .B(n32914), .C(n32915), .Y(n32912) );
  NOR2X1 U27287 ( .A(n32916), .B(n32917), .Y(n32915) );
  OAI22X1 U27288 ( .A(n25239), .B(n25316), .C(n29286), .D(n25318), .Y(n32917)
         );
  OAI22X1 U27289 ( .A(n32918), .B(n25320), .C(n25244), .D(n25322), .Y(n32916)
         );
  AOI22X1 U27290 ( .A(n25324), .B(reg_A[31]), .C(n25234), .D(reg_A[17]), .Y(
        n32914) );
  AOI22X1 U27291 ( .A(n25235), .B(reg_A[18]), .C(n25325), .D(reg_A[16]), .Y(
        n32913) );
  NAND3X1 U27292 ( .A(n32919), .B(n32920), .C(n32921), .Y(n32911) );
  NOR2X1 U27293 ( .A(n32922), .B(n32923), .Y(n32921) );
  OAI22X1 U27294 ( .A(n25331), .B(n25232), .C(n25243), .D(n25230), .Y(n32923)
         );
  OAI22X1 U27295 ( .A(n25334), .B(n25220), .C(n25336), .D(n30587), .Y(n32922)
         );
  AOI22X1 U27296 ( .A(n25242), .B(reg_A[25]), .C(n25338), .D(reg_A[26]), .Y(
        n32920) );
  AOI22X1 U27297 ( .A(reg_A[23]), .B(n25339), .C(reg_A[24]), .D(n25257), .Y(
        n32919) );
  AOI21X1 U27298 ( .A(reg_A[13]), .B(n25299), .C(n32924), .Y(n32906) );
  OAI22X1 U27299 ( .A(n25360), .B(n26677), .C(n27420), .D(n29265), .Y(n32924)
         );
  INVX1 U27300 ( .A(n25364), .Y(n27420) );
  NAND3X1 U27301 ( .A(n32925), .B(n32926), .C(n32927), .Y(n32904) );
  AOI21X1 U27302 ( .A(n32928), .B(n31822), .C(n32929), .Y(n32927) );
  OAI21X1 U27303 ( .A(n25177), .B(n32930), .C(n32931), .Y(n32929) );
  NAND2X1 U27304 ( .A(n29569), .B(n29565), .Y(n32930) );
  OAI21X1 U27305 ( .A(n25177), .B(n31833), .C(n32932), .Y(n31822) );
  NAND3X1 U27306 ( .A(n32933), .B(n32934), .C(reg_A[3]), .Y(n32932) );
  OAI21X1 U27307 ( .A(n25517), .B(n32935), .C(n31828), .Y(n32928) );
  OAI21X1 U27308 ( .A(n32936), .B(n32937), .C(reg_A[0]), .Y(n32926) );
  OAI21X1 U27309 ( .A(n25194), .B(n25794), .C(n32938), .Y(n32937) );
  AOI22X1 U27310 ( .A(n30621), .B(reg_B[7]), .C(n30910), .D(n32939), .Y(n32938) );
  INVX1 U27311 ( .A(n32940), .Y(n30621) );
  NAND3X1 U27312 ( .A(n30636), .B(n27943), .C(n32941), .Y(n32936) );
  OAI21X1 U27313 ( .A(n32942), .B(n32943), .C(n27358), .Y(n32941) );
  AOI21X1 U27314 ( .A(reg_A[2]), .B(n32944), .C(n32945), .Y(n32925) );
  AOI21X1 U27315 ( .A(n32946), .B(n25518), .C(n25130), .Y(n32945) );
  OAI21X1 U27316 ( .A(n32947), .B(n25517), .C(n32948), .Y(n32944) );
  NOR2X1 U27317 ( .A(n32949), .B(n25173), .Y(n32948) );
  NOR2X1 U27318 ( .A(n32950), .B(n25024), .Y(n25173) );
  INVX1 U27319 ( .A(n25566), .Y(n32949) );
  NOR2X1 U27320 ( .A(n32951), .B(n32952), .Y(n32902) );
  OAI21X1 U27321 ( .A(n27971), .B(n25147), .C(n32953), .Y(n32952) );
  AOI22X1 U27322 ( .A(reg_A[8]), .B(n29030), .C(reg_A[9]), .D(n29031), .Y(
        n32953) );
  OAI21X1 U27323 ( .A(n27512), .B(n27967), .C(n32954), .Y(n32951) );
  AOI22X1 U27324 ( .A(reg_A[14]), .B(n25300), .C(reg_A[12]), .D(n25301), .Y(
        n32954) );
  NOR2X1 U27325 ( .A(n32955), .B(n32956), .Y(n32901) );
  NAND2X1 U27326 ( .A(n32957), .B(n32958), .Y(n32956) );
  MUX2X1 U27327 ( .B(n32959), .A(n32960), .S(reg_B[7]), .Y(n32958) );
  NOR2X1 U27328 ( .A(n32961), .B(n26151), .Y(n32960) );
  NOR2X1 U27329 ( .A(n28213), .B(n31825), .Y(n32959) );
  AOI22X1 U27330 ( .A(reg_A[1]), .B(n30613), .C(reg_A[3]), .D(n30612), .Y(
        n31825) );
  MUX2X1 U27331 ( .B(n31820), .A(n32962), .S(reg_B[15]), .Y(n32957) );
  AND2X1 U27332 ( .A(n32963), .B(n26267), .Y(n32962) );
  NOR2X1 U27333 ( .A(n27354), .B(n32964), .Y(n31820) );
  INVX1 U27334 ( .A(n32965), .Y(n32964) );
  OAI21X1 U27335 ( .A(n25177), .B(n25197), .C(n32966), .Y(n32965) );
  NAND3X1 U27336 ( .A(n31796), .B(n29256), .C(reg_A[3]), .Y(n32966) );
  OAI21X1 U27337 ( .A(n32967), .B(n30547), .C(n32968), .Y(n32955) );
  AOI22X1 U27338 ( .A(reg_A[4]), .B(n25282), .C(n25382), .D(n32969), .Y(n32968) );
  NAND3X1 U27339 ( .A(n32970), .B(n32971), .C(n32972), .Y(n32969) );
  NOR2X1 U27340 ( .A(n32973), .B(n32974), .Y(n32972) );
  OAI21X1 U27341 ( .A(n32975), .B(n32976), .C(n32977), .Y(n32974) );
  OAI21X1 U27342 ( .A(n32978), .B(n32979), .C(n25044), .Y(n32977) );
  NAND2X1 U27343 ( .A(n32980), .B(n32981), .Y(n32979) );
  AOI22X1 U27344 ( .A(n30644), .B(n32982), .C(n26772), .D(n32983), .Y(n32981)
         );
  AOI22X1 U27345 ( .A(n32984), .B(reg_A[4]), .C(n32985), .D(reg_A[3]), .Y(
        n32980) );
  NAND2X1 U27346 ( .A(n32986), .B(n32987), .Y(n32978) );
  AOI22X1 U27347 ( .A(n32988), .B(n25258), .C(n29307), .D(n26761), .Y(n32987)
         );
  NOR2X1 U27348 ( .A(n26775), .B(n26677), .Y(n29307) );
  INVX1 U27349 ( .A(n30620), .Y(n32988) );
  AOI22X1 U27350 ( .A(n25101), .B(n28036), .C(reg_B[27]), .D(n32989), .Y(
        n32986) );
  NAND2X1 U27351 ( .A(n32990), .B(n32991), .Y(n28036) );
  AOI22X1 U27352 ( .A(n25156), .B(reg_A[7]), .C(n25142), .D(reg_A[8]), .Y(
        n32991) );
  AOI22X1 U27353 ( .A(n25258), .B(reg_A[9]), .C(reg_A[10]), .D(n26761), .Y(
        n32990) );
  INVX1 U27354 ( .A(n28024), .Y(n32975) );
  OAI21X1 U27355 ( .A(n25194), .B(n25147), .C(n32992), .Y(n28024) );
  AOI22X1 U27356 ( .A(reg_A[9]), .B(n26733), .C(n25172), .D(reg_A[8]), .Y(
        n32992) );
  OAI21X1 U27357 ( .A(n32993), .B(n25132), .C(n32994), .Y(n32973) );
  NAND3X1 U27358 ( .A(reg_B[12]), .B(n32995), .C(n25604), .Y(n32994) );
  INVX1 U27359 ( .A(n32996), .Y(n32995) );
  AOI22X1 U27360 ( .A(n32997), .B(n27986), .C(n28038), .D(n25116), .Y(n32993)
         );
  AOI22X1 U27361 ( .A(reg_A[5]), .B(n32998), .C(reg_A[4]), .D(n32999), .Y(
        n32971) );
  AOI22X1 U27362 ( .A(reg_A[6]), .B(n33000), .C(reg_A[3]), .D(n28040), .Y(
        n32970) );
  NAND3X1 U27363 ( .A(n33001), .B(n33002), .C(n33003), .Y(result[39]) );
  NOR2X1 U27364 ( .A(n33004), .B(n33005), .Y(n33003) );
  NAND2X1 U27365 ( .A(n33006), .B(n33007), .Y(n33005) );
  NOR2X1 U27366 ( .A(n33008), .B(n33009), .Y(n33007) );
  OAI21X1 U27367 ( .A(n25198), .B(n33010), .C(n33011), .Y(n33009) );
  OAI21X1 U27368 ( .A(n33012), .B(n33013), .C(n25382), .Y(n33011) );
  INVX1 U27369 ( .A(n33014), .Y(n33013) );
  AOI22X1 U27370 ( .A(n33015), .B(n33016), .C(n33017), .D(n33018), .Y(n33014)
         );
  OAI21X1 U27371 ( .A(n33019), .B(n33020), .C(n33021), .Y(n33012) );
  OAI21X1 U27372 ( .A(n33022), .B(n33023), .C(n25044), .Y(n33021) );
  OAI22X1 U27373 ( .A(n32580), .B(n32045), .C(n32044), .D(n32041), .Y(n33023)
         );
  INVX1 U27374 ( .A(n33024), .Y(n32044) );
  INVX1 U27375 ( .A(n33025), .Y(n32580) );
  OAI21X1 U27376 ( .A(n32527), .B(n32043), .C(n33026), .Y(n33022) );
  AOI22X1 U27377 ( .A(reg_B[59]), .B(n31236), .C(n30298), .D(n33027), .Y(
        n33026) );
  OAI21X1 U27378 ( .A(n32040), .B(n30220), .C(n33028), .Y(n31236) );
  AOI22X1 U27379 ( .A(reg_B[60]), .B(n29981), .C(n30325), .D(n32526), .Y(
        n33028) );
  INVX1 U27380 ( .A(n32046), .Y(n29981) );
  NAND2X1 U27381 ( .A(reg_A[63]), .B(n30107), .Y(n32046) );
  INVX1 U27382 ( .A(n33029), .Y(n32040) );
  NAND2X1 U27383 ( .A(n32110), .B(reg_A[47]), .Y(n33020) );
  AOI21X1 U27384 ( .A(n29987), .B(n33030), .C(n33031), .Y(n33010) );
  OAI22X1 U27385 ( .A(n32762), .B(n30320), .C(n32697), .D(n29970), .Y(n33031)
         );
  INVX1 U27386 ( .A(n32764), .Y(n32697) );
  OAI22X1 U27387 ( .A(n29976), .B(n30059), .C(n30393), .D(n32045), .Y(n32764)
         );
  INVX1 U27388 ( .A(n32889), .Y(n32762) );
  OAI21X1 U27389 ( .A(n27354), .B(n33032), .C(n33033), .Y(n33008) );
  OAI21X1 U27390 ( .A(n33034), .B(n33035), .C(reg_A[39]), .Y(n33033) );
  OAI21X1 U27391 ( .A(n28105), .B(n33036), .C(n33037), .Y(n33035) );
  AOI21X1 U27392 ( .A(n32299), .B(n33038), .C(n33039), .Y(n33032) );
  OAI22X1 U27393 ( .A(n32758), .B(n32253), .C(n32619), .D(n32134), .Y(n33039)
         );
  INVX1 U27394 ( .A(n32867), .Y(n32619) );
  OAI21X1 U27395 ( .A(n30059), .B(n32371), .C(n32798), .Y(n32867) );
  NAND2X1 U27396 ( .A(n32260), .B(reg_A[35]), .Y(n32798) );
  INVX1 U27397 ( .A(n32868), .Y(n32758) );
  AOI21X1 U27398 ( .A(n32357), .B(n33040), .C(n33041), .Y(n33006) );
  OAI21X1 U27399 ( .A(n27108), .B(n30394), .C(n33042), .Y(n33041) );
  OAI21X1 U27400 ( .A(n33043), .B(n33044), .C(n25999), .Y(n33042) );
  OAI22X1 U27401 ( .A(n25754), .B(n30170), .C(n31144), .D(n30057), .Y(n33044)
         );
  OAI22X1 U27402 ( .A(n30090), .B(n30058), .C(n27925), .D(n30060), .Y(n33043)
         );
  NAND3X1 U27403 ( .A(n33045), .B(n33046), .C(n33047), .Y(n33004) );
  NOR2X1 U27404 ( .A(n33048), .B(n33049), .Y(n33047) );
  OAI21X1 U27405 ( .A(n28516), .B(n33050), .C(n33051), .Y(n33049) );
  OAI21X1 U27406 ( .A(n33052), .B(n33053), .C(n27067), .Y(n33051) );
  OAI21X1 U27407 ( .A(n25060), .B(n30059), .C(n33054), .Y(n33053) );
  AOI22X1 U27408 ( .A(reg_A[35]), .B(n25749), .C(reg_A[34]), .D(n25750), .Y(
        n33054) );
  NAND2X1 U27409 ( .A(n33055), .B(n33056), .Y(n33052) );
  AOI22X1 U27410 ( .A(reg_A[38]), .B(n26803), .C(reg_A[36]), .D(n26804), .Y(
        n33056) );
  AOI22X1 U27411 ( .A(reg_A[37]), .B(n26927), .C(reg_A[33]), .D(n26878), .Y(
        n33055) );
  NOR2X1 U27412 ( .A(n33057), .B(n33058), .Y(n33050) );
  OAI21X1 U27413 ( .A(n25043), .B(n30059), .C(n33059), .Y(n33058) );
  AOI22X1 U27414 ( .A(reg_A[35]), .B(n25073), .C(reg_A[34]), .D(n25123), .Y(
        n33059) );
  NAND2X1 U27415 ( .A(n33060), .B(n33061), .Y(n33057) );
  AOI22X1 U27416 ( .A(reg_A[38]), .B(n25135), .C(reg_A[36]), .D(n25136), .Y(
        n33061) );
  AOI22X1 U27417 ( .A(reg_A[37]), .B(n25252), .C(reg_A[33]), .D(n25253), .Y(
        n33060) );
  INVX1 U27418 ( .A(n25119), .Y(n28516) );
  OAI21X1 U27419 ( .A(n33062), .B(n33063), .C(n33064), .Y(n33048) );
  NAND3X1 U27420 ( .A(n26186), .B(n33065), .C(reg_B[39]), .Y(n33064) );
  AOI22X1 U27421 ( .A(n33066), .B(reg_A[37]), .C(reg_B[37]), .D(n33067), .Y(
        n33062) );
  OAI21X1 U27422 ( .A(n28055), .B(n33068), .C(reg_A[32]), .Y(n33046) );
  OAI21X1 U27423 ( .A(n29973), .B(n31514), .C(n33069), .Y(n33068) );
  NAND3X1 U27424 ( .A(reg_B[45]), .B(n25188), .C(n32357), .Y(n33069) );
  AOI22X1 U27425 ( .A(n32033), .B(n27110), .C(n26504), .D(n33070), .Y(n33045)
         );
  OAI21X1 U27426 ( .A(n33071), .B(n33072), .C(n33073), .Y(n33070) );
  AOI22X1 U27427 ( .A(n33074), .B(n33075), .C(n33076), .D(n33077), .Y(n33073)
         );
  INVX1 U27428 ( .A(n33078), .Y(n33077) );
  NOR2X1 U27429 ( .A(n30393), .B(n33079), .Y(n33074) );
  MUX2X1 U27430 ( .B(n30059), .A(n30060), .S(reg_B[4]), .Y(n32033) );
  NOR2X1 U27431 ( .A(n33080), .B(n33081), .Y(n33002) );
  OAI21X1 U27432 ( .A(n27938), .B(n30463), .C(n33082), .Y(n33081) );
  AOI22X1 U27433 ( .A(reg_A[40]), .B(n27940), .C(reg_A[47]), .D(n25302), .Y(
        n33082) );
  NAND2X1 U27434 ( .A(n33083), .B(n33084), .Y(n33080) );
  INVX1 U27435 ( .A(n33085), .Y(n33084) );
  OAI21X1 U27436 ( .A(n25945), .B(n33086), .C(n33087), .Y(n33085) );
  OAI21X1 U27437 ( .A(n33088), .B(n33089), .C(n25310), .Y(n33087) );
  NAND3X1 U27438 ( .A(n33090), .B(n33091), .C(n33092), .Y(n33089) );
  NOR2X1 U27439 ( .A(n33093), .B(n33094), .Y(n33092) );
  OAI22X1 U27440 ( .A(n25036), .B(n30174), .C(n25473), .D(n30008), .Y(n33094)
         );
  OAI22X1 U27441 ( .A(n25037), .B(n29655), .C(n25320), .D(n30007), .Y(n33093)
         );
  AOI22X1 U27442 ( .A(reg_A[53]), .B(n25234), .C(reg_A[54]), .D(n25235), .Y(
        n33091) );
  AOI22X1 U27443 ( .A(reg_A[51]), .B(n25635), .C(reg_A[52]), .D(n25325), .Y(
        n33090) );
  NAND3X1 U27444 ( .A(n33095), .B(n33096), .C(n33097), .Y(n33088) );
  NOR2X1 U27445 ( .A(n33098), .B(n33099), .Y(n33097) );
  OAI22X1 U27446 ( .A(n25331), .B(n29990), .C(n25243), .D(n30219), .Y(n33099)
         );
  OAI22X1 U27447 ( .A(n25334), .B(n30043), .C(n25336), .D(n30254), .Y(n33098)
         );
  AOI22X1 U27448 ( .A(reg_A[61]), .B(n25242), .C(reg_A[62]), .D(n25338), .Y(
        n33096) );
  AOI22X1 U27449 ( .A(reg_A[59]), .B(n25339), .C(reg_A[60]), .D(n25257), .Y(
        n33095) );
  AOI22X1 U27450 ( .A(n27132), .B(reg_A[35]), .C(n33100), .D(n30847), .Y(
        n33083) );
  NOR2X1 U27451 ( .A(n33101), .B(n33102), .Y(n33001) );
  NAND2X1 U27452 ( .A(n33103), .B(n32885), .Y(n33102) );
  AOI22X1 U27453 ( .A(reg_A[45]), .B(n29031), .C(reg_A[46]), .D(n25293), .Y(
        n33103) );
  OAI21X1 U27454 ( .A(n25297), .B(n30067), .C(n33104), .Y(n33101) );
  AOI22X1 U27455 ( .A(reg_A[42]), .B(n29051), .C(reg_A[43]), .D(n29029), .Y(
        n33104) );
  NAND3X1 U27456 ( .A(n33105), .B(n33106), .C(n33107), .Y(result[38]) );
  NOR2X1 U27457 ( .A(n33108), .B(n33109), .Y(n33107) );
  NAND3X1 U27458 ( .A(n32885), .B(n33110), .C(n33111), .Y(n33109) );
  AOI21X1 U27459 ( .A(reg_A[33]), .B(n29130), .C(n33112), .Y(n33111) );
  OAI22X1 U27460 ( .A(n29129), .B(n30394), .C(n26781), .D(n30059), .Y(n33112)
         );
  INVX1 U27461 ( .A(n29248), .Y(n29130) );
  OAI21X1 U27462 ( .A(n33113), .B(n33114), .C(n25382), .Y(n33110) );
  OAI21X1 U27463 ( .A(n33115), .B(n33116), .C(n33117), .Y(n33114) );
  AOI22X1 U27464 ( .A(n33018), .B(n32673), .C(n32129), .D(n32268), .Y(n33117)
         );
  INVX1 U27465 ( .A(n32672), .Y(n32268) );
  OAI21X1 U27466 ( .A(n30060), .B(n33036), .C(n33118), .Y(n33113) );
  INVX1 U27467 ( .A(n33119), .Y(n33118) );
  OAI21X1 U27468 ( .A(n33120), .B(n30059), .C(n33121), .Y(n33119) );
  OAI21X1 U27469 ( .A(n33122), .B(n33123), .C(n25044), .Y(n33121) );
  OAI22X1 U27470 ( .A(n32686), .B(n32045), .C(n32246), .D(n32041), .Y(n33123)
         );
  INVX1 U27471 ( .A(n33124), .Y(n32246) );
  INVX1 U27472 ( .A(n33125), .Y(n32686) );
  OAI21X1 U27473 ( .A(n32626), .B(n32043), .C(n33126), .Y(n33122) );
  AOI22X1 U27474 ( .A(reg_B[59]), .B(n31265), .C(n30298), .D(n33127), .Y(
        n33126) );
  OAI21X1 U27475 ( .A(n32245), .B(n29975), .C(n33128), .Y(n31265) );
  AOI22X1 U27476 ( .A(n30326), .B(n32249), .C(n30324), .D(n32248), .Y(n33128)
         );
  INVX1 U27477 ( .A(n33129), .Y(n32245) );
  INVX1 U27478 ( .A(n32195), .Y(n32626) );
  INVX1 U27479 ( .A(n33130), .Y(n33036) );
  NAND3X1 U27480 ( .A(n33131), .B(n33132), .C(n33133), .Y(n33108) );
  AOI22X1 U27481 ( .A(reg_A[37]), .B(n29291), .C(reg_A[35]), .D(n29155), .Y(
        n33133) );
  OAI21X1 U27482 ( .A(n33134), .B(n33135), .C(n25310), .Y(n33132) );
  NAND3X1 U27483 ( .A(n33136), .B(n33137), .C(n33138), .Y(n33135) );
  NOR2X1 U27484 ( .A(n33139), .B(n33140), .Y(n33138) );
  OAI21X1 U27485 ( .A(n25043), .B(n30060), .C(n33141), .Y(n33140) );
  AOI22X1 U27486 ( .A(reg_A[50]), .B(n25635), .C(reg_A[51]), .D(n25325), .Y(
        n33141) );
  OAI21X1 U27487 ( .A(n25065), .B(n30299), .C(n33142), .Y(n33139) );
  AOI22X1 U27488 ( .A(reg_A[48]), .B(n25637), .C(reg_A[52]), .D(n25234), .Y(
        n33142) );
  NOR2X1 U27489 ( .A(n33143), .B(n33144), .Y(n33137) );
  OAI22X1 U27490 ( .A(n25028), .B(n30160), .C(n26431), .D(n30462), .Y(n33144)
         );
  OAI22X1 U27491 ( .A(n25030), .B(n30066), .C(n25131), .D(n30067), .Y(n33143)
         );
  AOI21X1 U27492 ( .A(reg_A[49]), .B(n25222), .C(n33145), .Y(n33136) );
  OAI22X1 U27493 ( .A(n25034), .B(n30069), .C(n25223), .D(n30068), .Y(n33145)
         );
  NAND3X1 U27494 ( .A(n33146), .B(n33147), .C(n33148), .Y(n33134) );
  NOR2X1 U27495 ( .A(n33149), .B(n33150), .Y(n33148) );
  OAI21X1 U27496 ( .A(n25040), .B(n30744), .C(n33151), .Y(n33150) );
  AOI22X1 U27497 ( .A(reg_A[39]), .B(n25135), .C(reg_A[41]), .D(n25136), .Y(
        n33151) );
  OAI21X1 U27498 ( .A(n25057), .B(n30016), .C(n33152), .Y(n33149) );
  AOI22X1 U27499 ( .A(reg_A[59]), .B(n25257), .C(reg_A[63]), .D(n25857), .Y(
        n33152) );
  NOR2X1 U27500 ( .A(n33153), .B(n33154), .Y(n33147) );
  OAI22X1 U27501 ( .A(n25331), .B(n30254), .C(n25243), .D(n29990), .Y(n33154)
         );
  OAI22X1 U27502 ( .A(n25334), .B(n30168), .C(n25336), .D(n30043), .Y(n33153)
         );
  AOI21X1 U27503 ( .A(reg_A[58]), .B(n25339), .C(n33155), .Y(n33146) );
  OAI22X1 U27504 ( .A(n25491), .B(n29989), .C(n25492), .D(n30015), .Y(n33155)
         );
  AOI22X1 U27505 ( .A(n29987), .B(n33100), .C(n25730), .D(n33156), .Y(n33131)
         );
  NAND3X1 U27506 ( .A(n33157), .B(n33158), .C(n33159), .Y(n33156) );
  NOR2X1 U27507 ( .A(n33160), .B(n33161), .Y(n33159) );
  OAI22X1 U27508 ( .A(n26936), .B(n30066), .C(n25745), .D(n30067), .Y(n33161)
         );
  OAI22X1 U27509 ( .A(n25746), .B(n30744), .C(n25747), .D(n30463), .Y(n33160)
         );
  AOI22X1 U27510 ( .A(reg_A[42]), .B(n25749), .C(reg_A[43]), .D(n25750), .Y(
        n33158) );
  AOI22X1 U27511 ( .A(reg_A[47]), .B(n25614), .C(reg_A[46]), .D(n25615), .Y(
        n33157) );
  OAI22X1 U27512 ( .A(n27438), .B(n33162), .C(n33163), .D(n26610), .Y(n33100)
         );
  INVX1 U27513 ( .A(n33164), .Y(n33162) );
  NOR2X1 U27514 ( .A(n33165), .B(n33166), .Y(n33106) );
  OAI21X1 U27515 ( .A(n33167), .B(n30058), .C(n33168), .Y(n33166) );
  INVX1 U27516 ( .A(n33169), .Y(n33168) );
  OAI22X1 U27517 ( .A(n33170), .B(n27354), .C(n33171), .D(n25198), .Y(n33169)
         );
  AOI22X1 U27518 ( .A(reg_B[63]), .B(n33172), .C(n32889), .D(n30846), .Y(
        n33171) );
  OAI21X1 U27519 ( .A(n30394), .B(n32045), .C(n33173), .Y(n32889) );
  AOI22X1 U27520 ( .A(n33174), .B(reg_B[47]), .C(n32868), .D(n32110), .Y(
        n33170) );
  OAI21X1 U27521 ( .A(n30060), .B(n32371), .C(n32805), .Y(n32868) );
  NAND2X1 U27522 ( .A(n32260), .B(reg_A[34]), .Y(n32805) );
  NOR2X1 U27523 ( .A(n33175), .B(n29220), .Y(n33167) );
  OAI21X1 U27524 ( .A(n33176), .B(n33177), .C(n33178), .Y(n33165) );
  AOI21X1 U27525 ( .A(n33179), .B(n33075), .C(n33180), .Y(n33178) );
  NOR2X1 U27526 ( .A(n33078), .B(n25031), .Y(n33179) );
  NAND2X1 U27527 ( .A(n33181), .B(n29315), .Y(n33177) );
  NOR2X1 U27528 ( .A(n33182), .B(n33183), .Y(n33105) );
  OAI21X1 U27529 ( .A(n33184), .B(n32066), .C(n33185), .Y(n33183) );
  OAI21X1 U27530 ( .A(n29127), .B(n33186), .C(reg_A[32]), .Y(n33185) );
  OAI22X1 U27531 ( .A(n27438), .B(n30255), .C(n32233), .D(n32571), .Y(n33186)
         );
  NAND2X1 U27532 ( .A(reg_B[61]), .B(reg_B[62]), .Y(n30255) );
  INVX1 U27533 ( .A(n33040), .Y(n33184) );
  OAI22X1 U27534 ( .A(n25794), .B(n33187), .C(n33188), .D(n26147), .Y(n33040)
         );
  OAI21X1 U27535 ( .A(n29207), .B(n30060), .C(n33189), .Y(n33182) );
  AOI22X1 U27536 ( .A(n32207), .B(n29209), .C(n33190), .D(n33065), .Y(n33189)
         );
  MUX2X1 U27537 ( .B(n33191), .A(n33078), .S(n33071), .Y(n33065) );
  MUX2X1 U27538 ( .B(reg_A[38]), .A(reg_A[34]), .S(reg_B[37]), .Y(n33078) );
  AND2X1 U27539 ( .A(n33192), .B(n33193), .Y(n32207) );
  AOI22X1 U27540 ( .A(n26601), .B(n30058), .C(n26602), .D(n30393), .Y(n33193)
         );
  AOI22X1 U27541 ( .A(n27012), .B(n30060), .C(n26597), .D(n30057), .Y(n33192)
         );
  INVX1 U27542 ( .A(n29325), .Y(n29207) );
  NAND2X1 U27543 ( .A(n33194), .B(n33195), .Y(n29325) );
  NAND3X1 U27544 ( .A(n33196), .B(n33197), .C(n33198), .Y(result[37]) );
  NOR2X1 U27545 ( .A(n33199), .B(n33200), .Y(n33198) );
  NAND3X1 U27546 ( .A(n33201), .B(n32885), .C(n33202), .Y(n33200) );
  AOI21X1 U27547 ( .A(n30261), .B(n33203), .C(n33204), .Y(n33202) );
  OAI21X1 U27548 ( .A(n33205), .B(n27152), .C(n33206), .Y(n33204) );
  OAI21X1 U27549 ( .A(n33207), .B(n33208), .C(n27358), .Y(n33206) );
  OAI21X1 U27550 ( .A(n29339), .B(n30057), .C(n33209), .Y(n33208) );
  AOI22X1 U27551 ( .A(reg_A[33]), .B(n25650), .C(reg_A[36]), .D(n29341), .Y(
        n33209) );
  NAND2X1 U27552 ( .A(n33210), .B(n33211), .Y(n33207) );
  AOI22X1 U27553 ( .A(n33212), .B(n29345), .C(reg_A[34]), .D(n29346), .Y(
        n33211) );
  INVX1 U27554 ( .A(n33086), .Y(n33212) );
  NAND2X1 U27555 ( .A(n33213), .B(n33214), .Y(n33086) );
  AOI22X1 U27556 ( .A(n26292), .B(n30170), .C(n26293), .D(n30057), .Y(n33214)
         );
  AOI22X1 U27557 ( .A(n26294), .B(n30395), .C(n26295), .D(n30058), .Y(n33213)
         );
  AOI22X1 U27558 ( .A(reg_A[35]), .B(n29349), .C(reg_A[32]), .D(n29350), .Y(
        n33210) );
  AND2X1 U27559 ( .A(n33215), .B(n33216), .Y(n33205) );
  NOR2X1 U27560 ( .A(n33217), .B(n33218), .Y(n33216) );
  OAI21X1 U27561 ( .A(n26801), .B(n30463), .C(n33219), .Y(n33218) );
  AOI22X1 U27562 ( .A(reg_A[43]), .B(n26878), .C(reg_A[44]), .D(n25613), .Y(
        n33219) );
  OAI21X1 U27563 ( .A(n25062), .B(n30059), .C(n33220), .Y(n33217) );
  AOI22X1 U27564 ( .A(reg_A[38]), .B(n26803), .C(reg_A[40]), .D(n26804), .Y(
        n33220) );
  NOR2X1 U27565 ( .A(n33221), .B(n33222), .Y(n33215) );
  OAI22X1 U27566 ( .A(n25736), .B(n30057), .C(n31398), .D(n30068), .Y(n33222)
         );
  OAI21X1 U27567 ( .A(n27252), .B(n30066), .C(n33223), .Y(n33221) );
  AOI22X1 U27568 ( .A(reg_A[42]), .B(n25750), .C(reg_A[46]), .D(n25614), .Y(
        n33223) );
  INVX1 U27569 ( .A(n31363), .Y(n30261) );
  AOI21X1 U27570 ( .A(n25188), .B(n32665), .C(n32569), .Y(n32885) );
  NOR2X1 U27571 ( .A(n32058), .B(n25024), .Y(n32569) );
  NAND2X1 U27572 ( .A(reg_A[32]), .B(n29994), .Y(n32058) );
  NOR2X1 U27573 ( .A(n32635), .B(n30395), .Y(n32665) );
  AOI22X1 U27574 ( .A(reg_A[38]), .B(n27402), .C(reg_A[39]), .D(n29361), .Y(
        n33201) );
  NAND2X1 U27575 ( .A(n33224), .B(n33225), .Y(n33199) );
  AOI21X1 U27576 ( .A(reg_B[39]), .B(n33226), .C(n33227), .Y(n33225) );
  OAI21X1 U27577 ( .A(n33228), .B(n30394), .C(n33229), .Y(n33227) );
  OAI21X1 U27578 ( .A(n33230), .B(n33231), .C(n25382), .Y(n33229) );
  OAI22X1 U27579 ( .A(n33232), .B(n33116), .C(n32315), .D(n33019), .Y(n33231)
         );
  INVX1 U27580 ( .A(n33233), .Y(n33230) );
  AOI22X1 U27581 ( .A(n33234), .B(n33235), .C(n32716), .D(n33018), .Y(n33233)
         );
  AOI21X1 U27582 ( .A(n32357), .B(n33236), .C(n33237), .Y(n33228) );
  OAI21X1 U27583 ( .A(n29976), .B(n31514), .C(n30636), .Y(n33237) );
  NAND2X1 U27584 ( .A(n30847), .B(n25932), .Y(n31514) );
  INVX1 U27585 ( .A(n32283), .Y(n33236) );
  NAND2X1 U27586 ( .A(n32261), .B(n25188), .Y(n32283) );
  AOI21X1 U27587 ( .A(n32157), .B(n33238), .C(n33239), .Y(n33224) );
  OAI21X1 U27588 ( .A(n33240), .B(n30057), .C(n33241), .Y(n33239) );
  OAI21X1 U27589 ( .A(n33242), .B(n33243), .C(n25310), .Y(n33241) );
  NAND3X1 U27590 ( .A(n33244), .B(n33245), .C(n33246), .Y(n33243) );
  NOR2X1 U27591 ( .A(n33247), .B(n33248), .Y(n33246) );
  OAI21X1 U27592 ( .A(n25043), .B(n30057), .C(n33249), .Y(n33248) );
  AOI22X1 U27593 ( .A(reg_A[49]), .B(n25635), .C(reg_A[50]), .D(n25325), .Y(
        n33249) );
  OAI21X1 U27594 ( .A(n25065), .B(n30378), .C(n33250), .Y(n33247) );
  AOI22X1 U27595 ( .A(reg_A[47]), .B(n25637), .C(reg_A[51]), .D(n25234), .Y(
        n33250) );
  NOR2X1 U27596 ( .A(n33251), .B(n33252), .Y(n33245) );
  OAI22X1 U27597 ( .A(n25028), .B(n30462), .C(n26431), .D(n30463), .Y(n33252)
         );
  OAI22X1 U27598 ( .A(n25030), .B(n30067), .C(n25131), .D(n30160), .Y(n33251)
         );
  AOI21X1 U27599 ( .A(reg_A[48]), .B(n25222), .C(n33253), .Y(n33244) );
  OAI22X1 U27600 ( .A(n25034), .B(n30066), .C(n25037), .D(n30069), .Y(n33253)
         );
  NAND3X1 U27601 ( .A(n33254), .B(n33255), .C(n33256), .Y(n33242) );
  NOR2X1 U27602 ( .A(n33257), .B(n33258), .Y(n33256) );
  OAI21X1 U27603 ( .A(n25238), .B(n29990), .C(n33259), .Y(n33258) );
  AOI22X1 U27604 ( .A(reg_A[59]), .B(n25242), .C(reg_A[60]), .D(n25338), .Y(
        n33259) );
  NAND2X1 U27605 ( .A(n33260), .B(n33261), .Y(n33257) );
  AOI22X1 U27606 ( .A(reg_A[54]), .B(n25246), .C(reg_A[53]), .D(n25247), .Y(
        n33261) );
  AOI22X1 U27607 ( .A(reg_A[56]), .B(n25487), .C(reg_A[55]), .D(n25241), .Y(
        n33260) );
  NOR2X1 U27608 ( .A(n33262), .B(n33263), .Y(n33255) );
  OAI22X1 U27609 ( .A(n25316), .B(n30007), .C(n25320), .D(n29989), .Y(n33263)
         );
  OAI22X1 U27610 ( .A(n25322), .B(n30016), .C(n26719), .D(n30219), .Y(n33262)
         );
  AOI21X1 U27611 ( .A(reg_A[39]), .B(n25252), .C(n33264), .Y(n33254) );
  OAI22X1 U27612 ( .A(n25041), .B(n30744), .C(n25042), .D(n30060), .Y(n33264)
         );
  INVX1 U27613 ( .A(n29393), .Y(n33240) );
  NOR2X1 U27614 ( .A(n33265), .B(n33266), .Y(n33197) );
  NAND3X1 U27615 ( .A(n33267), .B(n33268), .C(n33269), .Y(n33266) );
  OAI21X1 U27616 ( .A(n33175), .B(n29394), .C(reg_A[35]), .Y(n33269) );
  INVX1 U27617 ( .A(n33270), .Y(n33175) );
  NAND3X1 U27618 ( .A(n26504), .B(n33176), .C(n33066), .Y(n33270) );
  INVX1 U27619 ( .A(n33271), .Y(n33066) );
  NAND3X1 U27620 ( .A(n32109), .B(n25188), .C(n33272), .Y(n33268) );
  OAI21X1 U27621 ( .A(n30236), .B(n31076), .C(n33172), .Y(n33267) );
  MUX2X1 U27622 ( .B(n32887), .A(n33273), .S(reg_B[62]), .Y(n33172) );
  INVX1 U27623 ( .A(n33030), .Y(n32887) );
  OAI21X1 U27624 ( .A(n30170), .B(n32045), .C(n33274), .Y(n33030) );
  INVX1 U27625 ( .A(n30290), .Y(n30236) );
  NAND2X1 U27626 ( .A(n25932), .B(n30028), .Y(n30290) );
  OAI21X1 U27627 ( .A(n33072), .B(n33275), .C(n33276), .Y(n33265) );
  AOI21X1 U27628 ( .A(n33277), .B(n33174), .C(n33180), .Y(n33276) );
  INVX1 U27629 ( .A(n33278), .Y(n33180) );
  NAND3X1 U27630 ( .A(reg_A[32]), .B(n26504), .C(n33279), .Y(n33278) );
  NOR2X1 U27631 ( .A(n33079), .B(n33071), .Y(n33279) );
  OAI22X1 U27632 ( .A(reg_B[46]), .B(n32865), .C(n30393), .D(n32807), .Y(
        n33174) );
  INVX1 U27633 ( .A(n33038), .Y(n32865) );
  OAI22X1 U27634 ( .A(n30057), .B(n32371), .C(n30170), .D(n32416), .Y(n33038)
         );
  NOR2X1 U27635 ( .A(reg_B[47]), .B(n27354), .Y(n33277) );
  NAND2X1 U27636 ( .A(n26504), .B(n33071), .Y(n33275) );
  INVX1 U27637 ( .A(n33280), .Y(n33072) );
  MUX2X1 U27638 ( .B(n33281), .A(n33191), .S(reg_B[39]), .Y(n33280) );
  NOR2X1 U27639 ( .A(n33282), .B(n33283), .Y(n33196) );
  NAND2X1 U27640 ( .A(n33284), .B(n33285), .Y(n33283) );
  OAI21X1 U27641 ( .A(n33286), .B(n33287), .C(n26480), .Y(n33285) );
  OAI22X1 U27642 ( .A(n32721), .B(n32045), .C(n32308), .D(n32041), .Y(n33287)
         );
  INVX1 U27643 ( .A(n32723), .Y(n32308) );
  INVX1 U27644 ( .A(n33288), .Y(n32721) );
  OAI22X1 U27645 ( .A(n32726), .B(n32043), .C(n31402), .D(n30341), .Y(n33286)
         );
  INVX1 U27646 ( .A(n33289), .Y(n31402) );
  OAI21X1 U27647 ( .A(n32307), .B(n29975), .C(n33290), .Y(n33289) );
  AOI22X1 U27648 ( .A(n30326), .B(n32310), .C(n30324), .D(n30285), .Y(n33290)
         );
  INVX1 U27649 ( .A(n32725), .Y(n32307) );
  INVX1 U27650 ( .A(n32377), .Y(n32726) );
  AOI22X1 U27651 ( .A(n33190), .B(n33181), .C(reg_A[32]), .D(n33291), .Y(
        n33284) );
  OAI21X1 U27652 ( .A(n27438), .B(n31459), .C(n33292), .Y(n33291) );
  AOI21X1 U27653 ( .A(n33293), .B(reg_B[45]), .C(n29368), .Y(n33292) );
  INVX1 U27654 ( .A(n30649), .Y(n29368) );
  NOR2X1 U27655 ( .A(n32110), .B(n25032), .Y(n33293) );
  NAND2X1 U27656 ( .A(reg_B[61]), .B(n29970), .Y(n31459) );
  OAI22X1 U27657 ( .A(n30393), .B(n33271), .C(reg_B[38]), .D(n33281), .Y(
        n33181) );
  MUX2X1 U27658 ( .B(reg_A[37]), .A(reg_A[33]), .S(reg_B[37]), .Y(n33281) );
  OAI21X1 U27659 ( .A(n29397), .B(n30170), .C(n33294), .Y(n33282) );
  AOI22X1 U27660 ( .A(reg_A[36]), .B(n33295), .C(n33296), .D(n33297), .Y(
        n33294) );
  INVX1 U27661 ( .A(n32037), .Y(n33296) );
  OAI21X1 U27662 ( .A(n27438), .B(n32765), .C(n29366), .Y(n33295) );
  NAND2X1 U27663 ( .A(n33298), .B(n33299), .Y(result[36]) );
  NOR2X1 U27664 ( .A(n33300), .B(n33301), .Y(n33299) );
  NAND2X1 U27665 ( .A(n33302), .B(n33303), .Y(n33301) );
  NOR2X1 U27666 ( .A(n33304), .B(n33305), .Y(n33303) );
  OAI22X1 U27667 ( .A(n33306), .B(n30394), .C(n33307), .D(n30393), .Y(n33305)
         );
  INVX1 U27668 ( .A(n31793), .Y(n33306) );
  OAI21X1 U27669 ( .A(n27438), .B(n33308), .C(n33309), .Y(n33304) );
  OAI21X1 U27670 ( .A(n33310), .B(n33311), .C(reg_A[32]), .Y(n33309) );
  OAI21X1 U27671 ( .A(n25031), .B(n33079), .C(n31797), .Y(n33311) );
  OAI22X1 U27672 ( .A(n32261), .B(n25794), .C(n30298), .D(n27438), .Y(n33310)
         );
  AOI21X1 U27673 ( .A(reg_A[38]), .B(n25364), .C(n33312), .Y(n33302) );
  OAI21X1 U27674 ( .A(n33313), .B(n30170), .C(n33314), .Y(n33312) );
  OAI21X1 U27675 ( .A(n33315), .B(n33316), .C(n25310), .Y(n33314) );
  NAND3X1 U27676 ( .A(n33317), .B(n33318), .C(n33319), .Y(n33316) );
  NOR2X1 U27677 ( .A(n33320), .B(n33321), .Y(n33319) );
  OAI22X1 U27678 ( .A(n25316), .B(n30016), .C(n25318), .D(n30007), .Y(n33321)
         );
  OAI22X1 U27679 ( .A(n25320), .B(n30015), .C(n25322), .D(n29989), .Y(n33320)
         );
  AOI22X1 U27680 ( .A(reg_A[50]), .B(n25234), .C(reg_A[51]), .D(n25235), .Y(
        n33318) );
  AOI22X1 U27681 ( .A(reg_A[48]), .B(n25635), .C(reg_A[49]), .D(n25325), .Y(
        n33317) );
  NAND3X1 U27682 ( .A(n33322), .B(n33323), .C(n33324), .Y(n33315) );
  NOR2X1 U27683 ( .A(n33325), .B(n33326), .Y(n33324) );
  OAI22X1 U27684 ( .A(n25051), .B(n30168), .C(n25243), .D(n30043), .Y(n33326)
         );
  OAI22X1 U27685 ( .A(n25334), .B(n30378), .C(n25336), .D(n30299), .Y(n33325)
         );
  AOI22X1 U27686 ( .A(reg_A[58]), .B(n25242), .C(reg_A[59]), .D(n25338), .Y(
        n33323) );
  AOI22X1 U27687 ( .A(reg_A[56]), .B(n25339), .C(reg_A[57]), .D(n25257), .Y(
        n33322) );
  INVX1 U27688 ( .A(n31770), .Y(n33313) );
  NAND3X1 U27689 ( .A(n33327), .B(n33328), .C(n33329), .Y(n33300) );
  AOI21X1 U27690 ( .A(n25372), .B(n33330), .C(n33331), .Y(n33329) );
  OAI21X1 U27691 ( .A(n33332), .B(n26996), .C(n33333), .Y(n33331) );
  OAI21X1 U27692 ( .A(n33334), .B(n33335), .C(n25382), .Y(n33333) );
  OAI22X1 U27693 ( .A(n33336), .B(n33116), .C(n33337), .D(n33338), .Y(n33335)
         );
  OAI22X1 U27694 ( .A(n32899), .B(n33339), .C(n32892), .D(n33019), .Y(n33334)
         );
  INVX1 U27695 ( .A(n33340), .Y(n32899) );
  NOR2X1 U27696 ( .A(n33341), .B(n33342), .Y(n33332) );
  OAI22X1 U27697 ( .A(n32428), .B(n32041), .C(n33343), .D(n32043), .Y(n33342)
         );
  INVX1 U27698 ( .A(n32497), .Y(n33343) );
  INVX1 U27699 ( .A(n33344), .Y(n32428) );
  OAI22X1 U27700 ( .A(n32897), .B(n32045), .C(n31478), .D(n30341), .Y(n33341)
         );
  AOI21X1 U27701 ( .A(n32427), .B(n30325), .C(n33345), .Y(n31478) );
  OAI22X1 U27702 ( .A(n30220), .B(n32426), .C(n30136), .D(n30521), .Y(n33345)
         );
  INVX1 U27703 ( .A(n31044), .Y(n30521) );
  INVX1 U27704 ( .A(n31032), .Y(n32426) );
  INVX1 U27705 ( .A(n33346), .Y(n32897) );
  OAI21X1 U27706 ( .A(n33347), .B(n30095), .C(n33348), .Y(n33330) );
  AOI22X1 U27707 ( .A(n33349), .B(n33016), .C(n33350), .D(reg_A[36]), .Y(
        n33348) );
  INVX1 U27708 ( .A(n33116), .Y(n33016) );
  NOR2X1 U27709 ( .A(n30394), .B(n32066), .Y(n33349) );
  NAND2X1 U27710 ( .A(reg_B[63]), .B(n25044), .Y(n30095) );
  AOI22X1 U27711 ( .A(n33351), .B(reg_B[47]), .C(n33352), .D(n33297), .Y(
        n33328) );
  OAI22X1 U27712 ( .A(reg_B[46]), .B(n33188), .C(n30394), .D(n32807), .Y(
        n33297) );
  AOI21X1 U27713 ( .A(reg_A[32]), .B(n32260), .C(n33272), .Y(n33188) );
  INVX1 U27714 ( .A(n33187), .Y(n33272) );
  NAND2X1 U27715 ( .A(n32261), .B(reg_A[36]), .Y(n33187) );
  INVX1 U27716 ( .A(n33353), .Y(n33352) );
  NOR2X1 U27717 ( .A(n27354), .B(n33354), .Y(n33351) );
  AOI22X1 U27718 ( .A(n32504), .B(n29209), .C(reg_A[36]), .D(n33355), .Y(
        n33327) );
  NAND3X1 U27719 ( .A(n33037), .B(n33356), .C(n31790), .Y(n33355) );
  NOR2X1 U27720 ( .A(n25283), .B(n33357), .Y(n31790) );
  OAI21X1 U27721 ( .A(n29339), .B(n31658), .C(n33358), .Y(n33357) );
  NAND3X1 U27722 ( .A(n26504), .B(n33079), .C(n33075), .Y(n33037) );
  AND2X1 U27723 ( .A(n33359), .B(n33360), .Y(n32504) );
  AOI22X1 U27724 ( .A(n26601), .B(n30394), .C(n26602), .D(n30170), .Y(n33360)
         );
  AOI22X1 U27725 ( .A(n27012), .B(n30058), .C(n26597), .D(n30393), .Y(n33359)
         );
  NOR2X1 U27726 ( .A(n33361), .B(n33362), .Y(n33298) );
  NAND3X1 U27727 ( .A(n33363), .B(n33364), .C(n33365), .Y(n33362) );
  NOR2X1 U27728 ( .A(n33366), .B(n33367), .Y(n33365) );
  OAI22X1 U27729 ( .A(n33347), .B(n31363), .C(n33368), .D(n30198), .Y(n33367)
         );
  INVX1 U27730 ( .A(n33203), .Y(n33368) );
  OAI22X1 U27731 ( .A(reg_B[62]), .B(n33163), .C(n30394), .D(n33369), .Y(
        n33203) );
  AOI21X1 U27732 ( .A(reg_A[32]), .B(n32420), .C(n33164), .Y(n33163) );
  MUX2X1 U27733 ( .B(n33370), .A(n33371), .S(reg_B[39]), .Y(n33366) );
  NAND3X1 U27734 ( .A(n29315), .B(n33079), .C(n33067), .Y(n33371) );
  INVX1 U27735 ( .A(n33372), .Y(n33067) );
  INVX1 U27736 ( .A(n33226), .Y(n33370) );
  OAI21X1 U27737 ( .A(n33271), .B(n33373), .C(n33374), .Y(n33226) );
  NAND3X1 U27738 ( .A(n33375), .B(n33071), .C(n26186), .Y(n33374) );
  INVX1 U27739 ( .A(n33191), .Y(n33375) );
  MUX2X1 U27740 ( .B(reg_A[36]), .A(reg_A[32]), .S(reg_B[37]), .Y(n33191) );
  OAI21X1 U27741 ( .A(n26504), .B(n26186), .C(reg_A[34]), .Y(n33373) );
  AOI22X1 U27742 ( .A(reg_A[42]), .B(n29031), .C(reg_A[43]), .D(n25293), .Y(
        n33364) );
  AOI22X1 U27743 ( .A(reg_A[37]), .B(n25282), .C(n32157), .D(n33376), .Y(
        n33363) );
  INVX1 U27744 ( .A(n30524), .Y(n32157) );
  NAND2X1 U27745 ( .A(n30298), .B(n26480), .Y(n30524) );
  NAND3X1 U27746 ( .A(n33377), .B(n33378), .C(n33379), .Y(n33361) );
  AOI21X1 U27747 ( .A(reg_A[41]), .B(n29030), .C(n33380), .Y(n33379) );
  OAI22X1 U27748 ( .A(n27511), .B(n30744), .C(n27512), .D(n30067), .Y(n33380)
         );
  AOI22X1 U27749 ( .A(reg_A[39]), .B(n27622), .C(reg_A[46]), .D(n25299), .Y(
        n33378) );
  AOI22X1 U27750 ( .A(reg_A[47]), .B(n25300), .C(reg_A[45]), .D(n25301), .Y(
        n33377) );
  NAND3X1 U27751 ( .A(n33381), .B(n33382), .C(n33383), .Y(result[35]) );
  NOR2X1 U27752 ( .A(n33384), .B(n33385), .Y(n33383) );
  NAND3X1 U27753 ( .A(n33386), .B(n33387), .C(n33388), .Y(n33385) );
  AOI21X1 U27754 ( .A(n25310), .B(n33389), .C(n33390), .Y(n33388) );
  OAI22X1 U27755 ( .A(n25250), .B(n25583), .C(n29656), .D(n30395), .Y(n33390)
         );
  INVX1 U27756 ( .A(n25340), .Y(n29656) );
  NAND2X1 U27757 ( .A(n30636), .B(n33391), .Y(n25340) );
  OAI21X1 U27758 ( .A(n32943), .B(n33392), .C(n27358), .Y(n33391) );
  OR2X1 U27759 ( .A(n32942), .B(n33393), .Y(n33392) );
  NOR2X1 U27760 ( .A(n33394), .B(n33395), .Y(n32942) );
  NAND3X1 U27761 ( .A(n33396), .B(n33397), .C(n33398), .Y(n33389) );
  NOR2X1 U27762 ( .A(n33399), .B(n33400), .Y(n33398) );
  NAND3X1 U27763 ( .A(n33401), .B(n33402), .C(n33403), .Y(n33400) );
  AOI21X1 U27764 ( .A(reg_A[38]), .B(n25136), .C(n33404), .Y(n33403) );
  OAI22X1 U27765 ( .A(n25042), .B(n30058), .C(n25499), .D(n30007), .Y(n33404)
         );
  AOI22X1 U27766 ( .A(reg_A[60]), .B(n25857), .C(reg_A[59]), .D(n25647), .Y(
        n33402) );
  AOI22X1 U27767 ( .A(reg_A[62]), .B(n25648), .C(reg_A[61]), .D(n26432), .Y(
        n33401) );
  NAND3X1 U27768 ( .A(n33405), .B(n33406), .C(n33407), .Y(n33399) );
  NOR2X1 U27769 ( .A(n33408), .B(n33409), .Y(n33407) );
  OAI22X1 U27770 ( .A(n25051), .B(n30299), .C(n25243), .D(n30168), .Y(n33409)
         );
  OAI22X1 U27771 ( .A(n25334), .B(n30009), .C(n25336), .D(n30378), .Y(n33408)
         );
  AOI22X1 U27772 ( .A(reg_A[57]), .B(n25242), .C(reg_A[58]), .D(n25338), .Y(
        n33406) );
  AOI22X1 U27773 ( .A(reg_A[55]), .B(n25339), .C(reg_A[56]), .D(n25257), .Y(
        n33405) );
  NOR2X1 U27774 ( .A(n33410), .B(n33411), .Y(n33397) );
  OAI21X1 U27775 ( .A(n25034), .B(n30160), .C(n33412), .Y(n33411) );
  AOI22X1 U27776 ( .A(reg_A[40]), .B(n25123), .C(reg_A[44]), .D(n25629), .Y(
        n33412) );
  NAND2X1 U27777 ( .A(n33413), .B(n33414), .Y(n33410) );
  AOI22X1 U27778 ( .A(reg_A[37]), .B(n25252), .C(reg_A[41]), .D(n25253), .Y(
        n33414) );
  AOI22X1 U27779 ( .A(reg_A[42]), .B(n25628), .C(reg_A[39]), .D(n25068), .Y(
        n33413) );
  NOR2X1 U27780 ( .A(n33415), .B(n33416), .Y(n33396) );
  OAI21X1 U27781 ( .A(n25043), .B(n30393), .C(n33417), .Y(n33416) );
  AOI22X1 U27782 ( .A(reg_A[47]), .B(n25635), .C(reg_A[48]), .D(n25325), .Y(
        n33417) );
  NAND2X1 U27783 ( .A(n33418), .B(n33419), .Y(n33415) );
  AOI22X1 U27784 ( .A(reg_A[46]), .B(n25222), .C(reg_A[45]), .D(n25637), .Y(
        n33419) );
  AOI22X1 U27785 ( .A(reg_A[49]), .B(n25234), .C(reg_A[50]), .D(n25235), .Y(
        n33418) );
  OAI21X1 U27786 ( .A(n33420), .B(n33421), .C(n25372), .Y(n33387) );
  OAI21X1 U27787 ( .A(n33347), .B(n30327), .C(n33422), .Y(n33421) );
  AOI22X1 U27788 ( .A(reg_A[34]), .B(n33423), .C(reg_A[32]), .D(n33424), .Y(
        n33422) );
  OAI21X1 U27789 ( .A(n25403), .B(n30210), .C(n33425), .Y(n33424) );
  AOI22X1 U27790 ( .A(n33426), .B(n25589), .C(n32357), .D(n25604), .Y(n33425)
         );
  OAI21X1 U27791 ( .A(n25403), .B(n32765), .C(n33427), .Y(n33423) );
  NAND2X1 U27792 ( .A(n25044), .B(n30028), .Y(n30327) );
  INVX1 U27793 ( .A(n33428), .Y(n33347) );
  OAI21X1 U27794 ( .A(n25415), .B(n33429), .C(n33430), .Y(n33420) );
  AOI21X1 U27795 ( .A(n33431), .B(n33235), .C(n33432), .Y(n33430) );
  INVX1 U27796 ( .A(n33433), .Y(n33432) );
  NOR2X1 U27797 ( .A(reg_B[39]), .B(n33372), .Y(n33431) );
  NAND2X1 U27798 ( .A(n33434), .B(n32229), .Y(n33429) );
  OAI21X1 U27799 ( .A(n33435), .B(n33436), .C(n25730), .Y(n33386) );
  OR2X1 U27800 ( .A(n33437), .B(n33438), .Y(n33436) );
  OAI21X1 U27801 ( .A(n25060), .B(n30393), .C(n33439), .Y(n33438) );
  AOI22X1 U27802 ( .A(reg_A[45]), .B(n25607), .C(reg_A[47]), .D(n25609), .Y(
        n33439) );
  OAI21X1 U27803 ( .A(n29558), .B(n30069), .C(n33440), .Y(n33437) );
  AOI22X1 U27804 ( .A(reg_A[44]), .B(n25614), .C(reg_A[43]), .D(n25615), .Y(
        n33440) );
  NAND3X1 U27805 ( .A(n33441), .B(n33442), .C(n33443), .Y(n33435) );
  AOI21X1 U27806 ( .A(reg_A[40]), .B(n25750), .C(n33444), .Y(n33443) );
  OAI22X1 U27807 ( .A(n26801), .B(n30059), .C(n26936), .D(n30462), .Y(n33444)
         );
  AOI22X1 U27808 ( .A(reg_A[36]), .B(n26803), .C(reg_A[38]), .D(n26804), .Y(
        n33442) );
  AOI22X1 U27809 ( .A(reg_A[37]), .B(n26927), .C(reg_A[41]), .D(n26878), .Y(
        n33441) );
  OR2X1 U27810 ( .A(n33445), .B(n33446), .Y(n33384) );
  OAI21X1 U27811 ( .A(n33354), .B(n33353), .C(n33447), .Y(n33446) );
  OAI21X1 U27812 ( .A(n33448), .B(n33449), .C(n25382), .Y(n33447) );
  OAI21X1 U27813 ( .A(n33450), .B(n30393), .C(n33451), .Y(n33449) );
  AOI22X1 U27814 ( .A(reg_A[36]), .B(n33452), .C(reg_A[38]), .D(n33453), .Y(
        n33451) );
  NAND3X1 U27815 ( .A(n33454), .B(n33455), .C(n33456), .Y(n33448) );
  AOI22X1 U27816 ( .A(n33018), .B(n33015), .C(reg_A[37]), .D(n33457), .Y(
        n33456) );
  NAND2X1 U27817 ( .A(n33458), .B(n33459), .Y(n33015) );
  AOI22X1 U27818 ( .A(n32299), .B(reg_A[41]), .C(n32109), .D(reg_A[40]), .Y(
        n33459) );
  AOI22X1 U27819 ( .A(n32357), .B(reg_A[42]), .C(n32110), .D(reg_A[39]), .Y(
        n33458) );
  INVX1 U27820 ( .A(n33339), .Y(n33018) );
  NAND3X1 U27821 ( .A(n25604), .B(n32567), .C(reg_B[44]), .Y(n33455) );
  INVX1 U27822 ( .A(n33460), .Y(n32567) );
  MUX2X1 U27823 ( .B(n33017), .A(n33461), .S(reg_B[45]), .Y(n33460) );
  NOR2X1 U27824 ( .A(n30068), .B(n32134), .Y(n33461) );
  NAND2X1 U27825 ( .A(n33462), .B(n33463), .Y(n33017) );
  AOI22X1 U27826 ( .A(n32299), .B(reg_A[45]), .C(n32109), .D(reg_A[44]), .Y(
        n33463) );
  AOI22X1 U27827 ( .A(n32357), .B(reg_A[46]), .C(n32110), .D(reg_A[43]), .Y(
        n33462) );
  NAND3X1 U27828 ( .A(n33075), .B(reg_A[39]), .C(n33464), .Y(n33454) );
  INVX1 U27829 ( .A(n33434), .Y(n33354) );
  OAI21X1 U27830 ( .A(n30170), .B(n32807), .C(n33465), .Y(n33434) );
  NAND3X1 U27831 ( .A(reg_A[35]), .B(n32334), .C(n32261), .Y(n33465) );
  OAI21X1 U27832 ( .A(n33466), .B(n32037), .C(n33467), .Y(n33445) );
  AOI22X1 U27833 ( .A(n33468), .B(n33190), .C(n33469), .D(reg_B[39]), .Y(
        n33467) );
  AND2X1 U27834 ( .A(n33470), .B(n26186), .Y(n33469) );
  NOR2X1 U27835 ( .A(reg_B[37]), .B(n33372), .Y(n33468) );
  MUX2X1 U27836 ( .B(reg_A[35]), .A(reg_A[33]), .S(reg_B[38]), .Y(n33372) );
  NAND2X1 U27837 ( .A(reg_B[47]), .B(n26267), .Y(n32037) );
  NOR2X1 U27838 ( .A(n33471), .B(n33472), .Y(n33382) );
  OAI22X1 U27839 ( .A(n32818), .B(n30059), .C(n33473), .D(n31363), .Y(n33472)
         );
  NAND2X1 U27840 ( .A(reg_B[63]), .B(n25699), .Y(n31363) );
  OAI21X1 U27841 ( .A(n25279), .B(n33474), .C(n33475), .Y(n33471) );
  AOI22X1 U27842 ( .A(n26480), .B(n33476), .C(n31076), .D(n33428), .Y(n33475)
         );
  OAI21X1 U27843 ( .A(n30170), .B(n33369), .C(n33477), .Y(n33428) );
  NAND3X1 U27844 ( .A(n30117), .B(n30024), .C(reg_A[35]), .Y(n33477) );
  INVX1 U27845 ( .A(n30198), .Y(n31076) );
  NAND3X1 U27846 ( .A(n33478), .B(n33479), .C(n33480), .Y(n33476) );
  NOR2X1 U27847 ( .A(n33481), .B(n33482), .Y(n33480) );
  OAI22X1 U27848 ( .A(n32527), .B(n32041), .C(n33483), .D(n32045), .Y(n33482)
         );
  INVX1 U27849 ( .A(n33027), .Y(n33483) );
  NAND2X1 U27850 ( .A(n33484), .B(n33485), .Y(n33027) );
  AOI22X1 U27851 ( .A(reg_A[39]), .B(n30846), .C(n30212), .D(reg_A[40]), .Y(
        n33485) );
  AOI22X1 U27852 ( .A(reg_A[41]), .B(n29987), .C(n30847), .D(reg_A[42]), .Y(
        n33484) );
  INVX1 U27853 ( .A(n32158), .Y(n32527) );
  NAND2X1 U27854 ( .A(n33486), .B(n33487), .Y(n32158) );
  AOI22X1 U27855 ( .A(reg_A[47]), .B(n30846), .C(n30212), .D(reg_A[48]), .Y(
        n33487) );
  AOI22X1 U27856 ( .A(reg_A[49]), .B(n29987), .C(n30847), .D(reg_A[50]), .Y(
        n33486) );
  OAI22X1 U27857 ( .A(n30210), .B(n33173), .C(n30038), .D(n33274), .Y(n33481)
         );
  NAND2X1 U27858 ( .A(reg_A[38]), .B(n30298), .Y(n33173) );
  AOI22X1 U27859 ( .A(reg_B[59]), .B(n31625), .C(n30039), .D(n33025), .Y(
        n33479) );
  NAND2X1 U27860 ( .A(n33488), .B(n33489), .Y(n33025) );
  AOI22X1 U27861 ( .A(reg_A[43]), .B(n30846), .C(n30212), .D(reg_A[44]), .Y(
        n33489) );
  AOI22X1 U27862 ( .A(reg_A[45]), .B(n29987), .C(n30847), .D(reg_A[46]), .Y(
        n33488) );
  OAI21X1 U27863 ( .A(n30677), .B(n30853), .C(n33490), .Y(n31625) );
  AOI22X1 U27864 ( .A(n30325), .B(n33024), .C(n30326), .D(n32526), .Y(n33490)
         );
  NAND2X1 U27865 ( .A(n33491), .B(n33492), .Y(n32526) );
  AOI22X1 U27866 ( .A(reg_A[55]), .B(n30846), .C(n30212), .D(reg_A[56]), .Y(
        n33492) );
  AOI22X1 U27867 ( .A(reg_A[57]), .B(n29987), .C(n30847), .D(reg_A[58]), .Y(
        n33491) );
  NAND2X1 U27868 ( .A(n33493), .B(n33494), .Y(n33024) );
  AOI22X1 U27869 ( .A(reg_A[51]), .B(n30846), .C(n30212), .D(reg_A[52]), .Y(
        n33494) );
  AOI22X1 U27870 ( .A(reg_A[53]), .B(n29987), .C(n30847), .D(reg_A[54]), .Y(
        n33493) );
  AOI22X1 U27871 ( .A(n33029), .B(n29973), .C(n29991), .D(reg_A[63]), .Y(
        n30677) );
  INVX1 U27872 ( .A(n30032), .Y(n29991) );
  NAND2X1 U27873 ( .A(n30846), .B(reg_B[61]), .Y(n30032) );
  NAND2X1 U27874 ( .A(n33495), .B(n33496), .Y(n33029) );
  AOI22X1 U27875 ( .A(reg_A[59]), .B(n30846), .C(n30212), .D(reg_A[60]), .Y(
        n33496) );
  AOI22X1 U27876 ( .A(reg_A[61]), .B(n29987), .C(n30847), .D(reg_A[62]), .Y(
        n33495) );
  AOI22X1 U27877 ( .A(n33497), .B(reg_A[36]), .C(n33498), .D(reg_A[35]), .Y(
        n33478) );
  AOI21X1 U27878 ( .A(reg_A[35]), .B(n25284), .C(n33499), .Y(n33474) );
  OAI22X1 U27879 ( .A(n25286), .B(n30170), .C(n25288), .D(n30394), .Y(n33499)
         );
  INVX1 U27880 ( .A(n29568), .Y(n25288) );
  INVX1 U27881 ( .A(n29569), .Y(n25286) );
  NOR2X1 U27882 ( .A(n33500), .B(n33501), .Y(n33381) );
  OAI22X1 U27883 ( .A(n25717), .B(n30057), .C(n25718), .D(n30060), .Y(n33501)
         );
  OAI22X1 U27884 ( .A(n25719), .B(n30058), .C(n25795), .D(n30393), .Y(n33500)
         );
  NAND3X1 U27885 ( .A(n33502), .B(n33503), .C(n33504), .Y(result[34]) );
  NOR2X1 U27886 ( .A(n33505), .B(n33506), .Y(n33504) );
  OAI21X1 U27887 ( .A(n33507), .B(n30931), .C(n33508), .Y(n33506) );
  INVX1 U27888 ( .A(n33509), .Y(n33508) );
  NOR2X1 U27889 ( .A(n33510), .B(n33511), .Y(n33507) );
  NAND3X1 U27890 ( .A(n33512), .B(n33513), .C(n33514), .Y(n33511) );
  AOI21X1 U27891 ( .A(reg_A[34]), .B(n25434), .C(n33515), .Y(n33514) );
  OAI22X1 U27892 ( .A(n28353), .B(n30058), .C(n25205), .D(n30060), .Y(n33515)
         );
  AOI22X1 U27893 ( .A(n25097), .B(n33516), .C(reg_A[39]), .D(n28355), .Y(
        n33513) );
  NAND2X1 U27894 ( .A(n33517), .B(n33518), .Y(n33516) );
  NOR2X1 U27895 ( .A(n33519), .B(n33520), .Y(n33518) );
  NAND3X1 U27896 ( .A(n33521), .B(n33522), .C(n33523), .Y(n33520) );
  AOI21X1 U27897 ( .A(reg_A[49]), .B(n25235), .C(n33524), .Y(n33523) );
  OAI22X1 U27898 ( .A(n25334), .B(n30008), .C(n25336), .D(n30009), .Y(n33524)
         );
  AOI22X1 U27899 ( .A(reg_A[53]), .B(n25487), .C(reg_A[52]), .D(n25241), .Y(
        n33522) );
  AOI22X1 U27900 ( .A(reg_A[54]), .B(n25339), .C(reg_A[55]), .D(n25257), .Y(
        n33521) );
  NAND3X1 U27901 ( .A(n33525), .B(n33526), .C(n33527), .Y(n33519) );
  NOR2X1 U27902 ( .A(n33528), .B(n33529), .Y(n33527) );
  OAI22X1 U27903 ( .A(n25316), .B(n30015), .C(n25318), .D(n29989), .Y(n33529)
         );
  INVX1 U27904 ( .A(reg_A[60]), .Y(n30015) );
  OAI22X1 U27905 ( .A(n25498), .B(n30007), .C(n25499), .D(n30016), .Y(n33528)
         );
  AOI22X1 U27906 ( .A(reg_A[59]), .B(n25857), .C(reg_A[58]), .D(n25647), .Y(
        n33526) );
  AOI22X1 U27907 ( .A(reg_A[56]), .B(n25242), .C(reg_A[57]), .D(n25338), .Y(
        n33525) );
  NOR2X1 U27908 ( .A(n33530), .B(n33531), .Y(n33517) );
  NAND3X1 U27909 ( .A(n33532), .B(n33533), .C(n33534), .Y(n33531) );
  AOI21X1 U27910 ( .A(reg_A[34]), .B(n25125), .C(n33535), .Y(n33534) );
  OAI22X1 U27911 ( .A(n25040), .B(n30058), .C(n25042), .D(n30393), .Y(n33535)
         );
  AOI22X1 U27912 ( .A(reg_A[37]), .B(n25136), .C(reg_A[40]), .D(n25253), .Y(
        n33533) );
  AOI22X1 U27913 ( .A(reg_A[38]), .B(n25073), .C(reg_A[39]), .D(n25123), .Y(
        n33532) );
  NAND3X1 U27914 ( .A(n33536), .B(n33537), .C(n33538), .Y(n33530) );
  NOR2X1 U27915 ( .A(n33539), .B(n33540), .Y(n33538) );
  OAI22X1 U27916 ( .A(n25064), .B(n30069), .C(n25473), .D(n30066), .Y(n33540)
         );
  OAI22X1 U27917 ( .A(n25039), .B(n30068), .C(n25475), .D(n29655), .Y(n33539)
         );
  AOI22X1 U27918 ( .A(reg_A[43]), .B(n25629), .C(reg_A[44]), .D(n25637), .Y(
        n33537) );
  AOI22X1 U27919 ( .A(reg_A[41]), .B(n25628), .C(reg_A[42]), .D(n25124), .Y(
        n33536) );
  AOI22X1 U27920 ( .A(reg_A[35]), .B(n25441), .C(reg_A[37]), .D(n27241), .Y(
        n33512) );
  NAND3X1 U27921 ( .A(n33541), .B(n33542), .C(n33543), .Y(n33510) );
  NOR2X1 U27922 ( .A(n33544), .B(n33545), .Y(n33543) );
  OAI22X1 U27923 ( .A(n30444), .B(n30462), .C(n26229), .D(n30160), .Y(n33545)
         );
  INVX1 U27924 ( .A(reg_A[43]), .Y(n30160) );
  INVX1 U27925 ( .A(reg_A[42]), .Y(n30462) );
  OAI22X1 U27926 ( .A(n25451), .B(n30069), .C(n25453), .D(n30068), .Y(n33544)
         );
  AOI22X1 U27927 ( .A(reg_A[41]), .B(n25502), .C(reg_A[45]), .D(n25503), .Y(
        n33542) );
  AOI22X1 U27928 ( .A(reg_A[44]), .B(n25439), .C(reg_A[40]), .D(n25440), .Y(
        n33541) );
  OAI21X1 U27929 ( .A(n33473), .B(n30198), .C(n33546), .Y(n33505) );
  OAI21X1 U27930 ( .A(n33547), .B(n33548), .C(n25382), .Y(n33546) );
  NAND2X1 U27931 ( .A(n33549), .B(n33550), .Y(n33548) );
  AOI22X1 U27932 ( .A(reg_A[36]), .B(n33457), .C(reg_A[35]), .D(n33452), .Y(
        n33550) );
  AOI22X1 U27933 ( .A(reg_A[37]), .B(n33453), .C(reg_A[34]), .D(n33551), .Y(
        n33549) );
  OR2X1 U27934 ( .A(n33552), .B(n33553), .Y(n33547) );
  OAI21X1 U27935 ( .A(n33115), .B(n33339), .C(n33554), .Y(n33553) );
  OAI21X1 U27936 ( .A(n33555), .B(n33556), .C(n25044), .Y(n33554) );
  NAND2X1 U27937 ( .A(n33557), .B(n33558), .Y(n33556) );
  AOI22X1 U27938 ( .A(n30039), .B(n33125), .C(n33164), .D(n29987), .Y(n33558)
         );
  NAND2X1 U27939 ( .A(n33559), .B(n33560), .Y(n33125) );
  AOI22X1 U27940 ( .A(reg_A[42]), .B(n30846), .C(n30212), .D(reg_A[43]), .Y(
        n33560) );
  AOI22X1 U27941 ( .A(reg_A[44]), .B(n29987), .C(n30847), .D(reg_A[45]), .Y(
        n33559) );
  AOI22X1 U27942 ( .A(n33497), .B(reg_A[35]), .C(n33498), .D(reg_A[34]), .Y(
        n33557) );
  NAND2X1 U27943 ( .A(n33561), .B(n33562), .Y(n33555) );
  AOI22X1 U27944 ( .A(n33563), .B(n30847), .C(n32420), .D(n33127), .Y(n33562)
         );
  NAND2X1 U27945 ( .A(n33564), .B(n33565), .Y(n33127) );
  AOI22X1 U27946 ( .A(reg_A[38]), .B(n30846), .C(n30212), .D(reg_A[39]), .Y(
        n33565) );
  AOI22X1 U27947 ( .A(reg_A[40]), .B(n29987), .C(n30847), .D(reg_A[41]), .Y(
        n33564) );
  INVX1 U27948 ( .A(n33274), .Y(n33563) );
  NAND2X1 U27949 ( .A(reg_A[37]), .B(n30298), .Y(n33274) );
  AOI22X1 U27950 ( .A(n32724), .B(n32195), .C(reg_B[59]), .D(n31727), .Y(
        n33561) );
  NAND2X1 U27951 ( .A(n33566), .B(n33567), .Y(n31727) );
  AOI22X1 U27952 ( .A(n30323), .B(n32248), .C(n30324), .D(n32249), .Y(n33567)
         );
  NAND2X1 U27953 ( .A(n33568), .B(n33569), .Y(n32249) );
  AOI22X1 U27954 ( .A(reg_A[58]), .B(n30846), .C(n30212), .D(reg_A[59]), .Y(
        n33569) );
  AOI22X1 U27955 ( .A(reg_A[60]), .B(n29987), .C(n30847), .D(reg_A[61]), .Y(
        n33568) );
  OAI22X1 U27956 ( .A(n30007), .B(n30320), .C(n29970), .D(n30016), .Y(n32248)
         );
  AOI22X1 U27957 ( .A(n30325), .B(n33124), .C(n30326), .D(n33129), .Y(n33566)
         );
  NAND2X1 U27958 ( .A(n33570), .B(n33571), .Y(n33129) );
  AOI22X1 U27959 ( .A(reg_A[54]), .B(n30846), .C(n30212), .D(reg_A[55]), .Y(
        n33571) );
  AOI22X1 U27960 ( .A(reg_A[56]), .B(n29987), .C(n30847), .D(reg_A[57]), .Y(
        n33570) );
  NAND2X1 U27961 ( .A(n33572), .B(n33573), .Y(n33124) );
  AOI22X1 U27962 ( .A(reg_A[50]), .B(n30846), .C(n30212), .D(reg_A[51]), .Y(
        n33573) );
  AOI22X1 U27963 ( .A(reg_A[52]), .B(n29987), .C(n30847), .D(reg_A[53]), .Y(
        n33572) );
  NAND2X1 U27964 ( .A(n33574), .B(n33575), .Y(n32195) );
  AOI22X1 U27965 ( .A(reg_A[46]), .B(n30846), .C(n30212), .D(reg_A[47]), .Y(
        n33575) );
  AOI22X1 U27966 ( .A(n29987), .B(reg_A[48]), .C(n30847), .D(reg_A[49]), .Y(
        n33574) );
  AND2X1 U27967 ( .A(n33576), .B(n33577), .Y(n33115) );
  AOI22X1 U27968 ( .A(n32299), .B(reg_A[40]), .C(n32109), .D(reg_A[39]), .Y(
        n33577) );
  AOI22X1 U27969 ( .A(n32357), .B(reg_A[41]), .C(n32110), .D(reg_A[38]), .Y(
        n33576) );
  OAI21X1 U27970 ( .A(n32672), .B(n32126), .C(n33578), .Y(n33552) );
  AOI22X1 U27971 ( .A(n33464), .B(n33579), .C(n32129), .D(n32673), .Y(n33578)
         );
  NAND3X1 U27972 ( .A(n32221), .B(n32631), .C(n33580), .Y(n32673) );
  INVX1 U27973 ( .A(n33581), .Y(n33580) );
  OAI21X1 U27974 ( .A(n32240), .B(n30066), .C(n32440), .Y(n33581) );
  NAND2X1 U27975 ( .A(n32109), .B(reg_A[43]), .Y(n32440) );
  NAND2X1 U27976 ( .A(n32110), .B(reg_A[42]), .Y(n32631) );
  NAND2X1 U27977 ( .A(n32299), .B(reg_A[44]), .Y(n32221) );
  INVX1 U27978 ( .A(n33582), .Y(n33579) );
  AOI22X1 U27979 ( .A(reg_A[38]), .B(n33075), .C(reg_A[39]), .D(n33076), .Y(
        n33582) );
  AOI21X1 U27980 ( .A(reg_A[47]), .B(n32109), .C(n32219), .Y(n32672) );
  NOR2X1 U27981 ( .A(n32134), .B(n30069), .Y(n32219) );
  NAND2X1 U27982 ( .A(n25699), .B(n30028), .Y(n30198) );
  INVX1 U27983 ( .A(n33583), .Y(n33473) );
  OAI21X1 U27984 ( .A(n30395), .B(n33369), .C(n33584), .Y(n33583) );
  NAND3X1 U27985 ( .A(n30117), .B(n30024), .C(reg_A[34]), .Y(n33584) );
  NAND2X1 U27986 ( .A(n30298), .B(reg_B[62]), .Y(n33369) );
  AOI21X1 U27987 ( .A(n33190), .B(n33470), .C(n33585), .Y(n33503) );
  OAI21X1 U27988 ( .A(n33466), .B(n33353), .C(n33586), .Y(n33585) );
  OAI21X1 U27989 ( .A(n33587), .B(n33588), .C(reg_A[32]), .Y(n33586) );
  OAI21X1 U27990 ( .A(n27438), .B(n30293), .C(n25528), .Y(n33588) );
  AND2X1 U27991 ( .A(n29513), .B(n33589), .Y(n25528) );
  OAI21X1 U27992 ( .A(n32943), .B(n33590), .C(n27358), .Y(n33589) );
  NAND2X1 U27993 ( .A(n33591), .B(n33592), .Y(n33590) );
  OAI21X1 U27994 ( .A(n25031), .B(n33071), .C(n32571), .Y(n33587) );
  NAND2X1 U27995 ( .A(reg_B[46]), .B(n25188), .Y(n32571) );
  NAND2X1 U27996 ( .A(n26267), .B(n32229), .Y(n33353) );
  INVX1 U27997 ( .A(n33593), .Y(n33466) );
  OAI21X1 U27998 ( .A(n30395), .B(n32807), .C(n33594), .Y(n33593) );
  NAND3X1 U27999 ( .A(reg_A[34]), .B(n32334), .C(n32261), .Y(n33594) );
  NAND2X1 U28000 ( .A(n32261), .B(reg_B[46]), .Y(n32807) );
  OAI21X1 U28001 ( .A(n30395), .B(n33271), .C(n33595), .Y(n33470) );
  NAND3X1 U28002 ( .A(n33079), .B(n33071), .C(reg_A[34]), .Y(n33595) );
  NAND2X1 U28003 ( .A(reg_B[38]), .B(n33079), .Y(n33271) );
  INVX1 U28004 ( .A(n33063), .Y(n33190) );
  NAND2X1 U28005 ( .A(n26186), .B(n33176), .Y(n33063) );
  AOI22X1 U28006 ( .A(reg_A[34]), .B(n33596), .C(reg_A[33]), .D(n33597), .Y(
        n33502) );
  OAI21X1 U28007 ( .A(n25198), .B(n32765), .C(n33598), .Y(n33597) );
  INVX1 U28008 ( .A(n33599), .Y(n33598) );
  OAI21X1 U28009 ( .A(n33600), .B(n33427), .C(n25566), .Y(n33599) );
  INVX1 U28010 ( .A(n33452), .Y(n33427) );
  OAI21X1 U28011 ( .A(n33450), .B(n25517), .C(n33601), .Y(n33596) );
  NOR2X1 U28012 ( .A(n33602), .B(n32825), .Y(n33601) );
  INVX1 U28013 ( .A(n33356), .Y(n32825) );
  NAND2X1 U28014 ( .A(n33498), .B(n25932), .Y(n33356) );
  NAND3X1 U28015 ( .A(n33603), .B(n33604), .C(n33605), .Y(result[33]) );
  NOR2X1 U28016 ( .A(n33606), .B(n33607), .Y(n33605) );
  OAI22X1 U28017 ( .A(n29765), .B(n30058), .C(n29766), .D(n30393), .Y(n33607)
         );
  NAND3X1 U28018 ( .A(n33608), .B(n33609), .C(n33610), .Y(n33606) );
  OAI21X1 U28019 ( .A(n29773), .B(n33611), .C(reg_A[33]), .Y(n33610) );
  OAI22X1 U28020 ( .A(n25198), .B(n33612), .C(n33450), .D(n33600), .Y(n33611)
         );
  OAI21X1 U28021 ( .A(n29566), .B(n31658), .C(n33358), .Y(n29773) );
  OAI21X1 U28022 ( .A(n33613), .B(n33614), .C(reg_A[32]), .Y(n33609) );
  NAND2X1 U28023 ( .A(n33615), .B(n25693), .Y(n33614) );
  INVX1 U28024 ( .A(n33616), .Y(n25693) );
  OAI21X1 U28025 ( .A(n33617), .B(n31658), .C(n29366), .Y(n33616) );
  AOI21X1 U28026 ( .A(n25044), .B(n25043), .C(n33618), .Y(n33617) );
  AOI22X1 U28027 ( .A(n25188), .B(n32134), .C(n26504), .D(n33619), .Y(n33615)
         );
  OAI21X1 U28028 ( .A(n30846), .B(n27438), .C(n33620), .Y(n33613) );
  AOI22X1 U28029 ( .A(n25170), .B(n33452), .C(n33497), .D(n25699), .Y(n33620)
         );
  NAND2X1 U28030 ( .A(reg_A[39]), .B(n29779), .Y(n33608) );
  AOI21X1 U28031 ( .A(n25203), .B(n33621), .C(n33622), .Y(n33604) );
  OAI22X1 U28032 ( .A(n25652), .B(n30060), .C(n29782), .D(n30057), .Y(n33622)
         );
  NAND3X1 U28033 ( .A(n33623), .B(n33624), .C(n33625), .Y(n33621) );
  NOR2X1 U28034 ( .A(n33626), .B(n33627), .Y(n33625) );
  OAI22X1 U28035 ( .A(n25598), .B(n30393), .C(n25599), .D(n30058), .Y(n33627)
         );
  OAI21X1 U28036 ( .A(n25600), .B(n30060), .C(n33628), .Y(n33626) );
  OAI21X1 U28037 ( .A(n33629), .B(n33630), .C(n25604), .Y(n33628) );
  NAND2X1 U28038 ( .A(n33631), .B(n33632), .Y(n33630) );
  AOI22X1 U28039 ( .A(reg_A[43]), .B(n25607), .C(reg_A[47]), .D(n25608), .Y(
        n33632) );
  AOI22X1 U28040 ( .A(reg_A[45]), .B(n25609), .C(reg_A[46]), .D(n25610), .Y(
        n33631) );
  NAND2X1 U28041 ( .A(n33633), .B(n33634), .Y(n33629) );
  AOI22X1 U28042 ( .A(reg_A[40]), .B(n25613), .C(reg_A[42]), .D(n25614), .Y(
        n33634) );
  AOI22X1 U28043 ( .A(reg_A[41]), .B(n25615), .C(reg_A[44]), .D(n25616), .Y(
        n33633) );
  AOI21X1 U28044 ( .A(reg_A[34]), .B(n25617), .C(n33635), .Y(n33624) );
  OAI21X1 U28045 ( .A(n25619), .B(n30170), .C(n33636), .Y(n33635) );
  OAI21X1 U28046 ( .A(n33637), .B(n33638), .C(n25044), .Y(n33636) );
  NAND2X1 U28047 ( .A(n33639), .B(n33640), .Y(n33638) );
  NOR2X1 U28048 ( .A(n33641), .B(n33642), .Y(n33640) );
  OAI21X1 U28049 ( .A(n25034), .B(n30463), .C(n33643), .Y(n33642) );
  AOI22X1 U28050 ( .A(reg_A[40]), .B(n25628), .C(reg_A[42]), .D(n25629), .Y(
        n33643) );
  OAI21X1 U28051 ( .A(n25498), .B(n30016), .C(n33644), .Y(n33641) );
  AOI22X1 U28052 ( .A(reg_A[63]), .B(n25631), .C(reg_A[61]), .D(n25324), .Y(
        n33644) );
  INVX1 U28053 ( .A(reg_A[62]), .Y(n30016) );
  NOR2X1 U28054 ( .A(n33645), .B(n33646), .Y(n33639) );
  OAI21X1 U28055 ( .A(n25039), .B(n30069), .C(n33647), .Y(n33646) );
  AOI22X1 U28056 ( .A(reg_A[48]), .B(n25235), .C(reg_A[45]), .D(n25635), .Y(
        n33647) );
  INVX1 U28057 ( .A(reg_A[46]), .Y(n30069) );
  OAI21X1 U28058 ( .A(n25035), .B(n30068), .C(n33648), .Y(n33645) );
  AOI22X1 U28059 ( .A(reg_A[44]), .B(n25222), .C(reg_A[43]), .D(n25637), .Y(
        n33648) );
  NAND2X1 U28060 ( .A(n33649), .B(n33650), .Y(n33637) );
  NOR2X1 U28061 ( .A(n33651), .B(n33652), .Y(n33650) );
  OAI21X1 U28062 ( .A(n25050), .B(n30254), .C(n33653), .Y(n33652) );
  AOI22X1 U28063 ( .A(reg_A[51]), .B(n25241), .C(reg_A[55]), .D(n25242), .Y(
        n33653) );
  OAI21X1 U28064 ( .A(n25038), .B(n30378), .C(n33654), .Y(n33651) );
  AOI22X1 U28065 ( .A(reg_A[50]), .B(n25246), .C(reg_A[49]), .D(n25247), .Y(
        n33654) );
  NOR2X1 U28066 ( .A(n33655), .B(n33656), .Y(n33649) );
  OAI21X1 U28067 ( .A(n25059), .B(n29984), .C(n33657), .Y(n33656) );
  AOI22X1 U28068 ( .A(reg_A[57]), .B(n25647), .C(reg_A[60]), .D(n25648), .Y(
        n33657) );
  OAI21X1 U28069 ( .A(n25054), .B(n30219), .C(n33658), .Y(n33655) );
  AOI22X1 U28070 ( .A(reg_A[53]), .B(n25339), .C(reg_A[54]), .D(n25257), .Y(
        n33658) );
  AOI22X1 U28071 ( .A(reg_A[37]), .B(n25650), .C(reg_A[39]), .D(n25651), .Y(
        n33623) );
  AOI21X1 U28072 ( .A(n25382), .B(n33659), .C(n33509), .Y(n33603) );
  OAI22X1 U28073 ( .A(n25517), .B(n33433), .C(n25250), .D(n25583), .Y(n33509)
         );
  OAI21X1 U28074 ( .A(n33660), .B(n33661), .C(reg_A[32]), .Y(n33433) );
  OAI21X1 U28075 ( .A(n30298), .B(n25403), .C(n33662), .Y(n33661) );
  NOR2X1 U28076 ( .A(n32261), .B(n25415), .Y(n33660) );
  NAND3X1 U28077 ( .A(n33663), .B(n33664), .C(n33665), .Y(n33659) );
  NOR2X1 U28078 ( .A(n33666), .B(n33667), .Y(n33665) );
  OAI21X1 U28079 ( .A(n33232), .B(n33339), .C(n33668), .Y(n33667) );
  OAI21X1 U28080 ( .A(n33669), .B(n33670), .C(n25044), .Y(n33668) );
  NAND2X1 U28081 ( .A(n33671), .B(n33672), .Y(n33670) );
  AOI22X1 U28082 ( .A(reg_B[59]), .B(n31896), .C(n30039), .D(n33288), .Y(
        n33672) );
  NAND2X1 U28083 ( .A(n33673), .B(n33674), .Y(n33288) );
  AOI22X1 U28084 ( .A(reg_A[41]), .B(n30846), .C(n30212), .D(reg_A[42]), .Y(
        n33674) );
  AOI22X1 U28085 ( .A(reg_A[43]), .B(n29987), .C(n30847), .D(reg_A[44]), .Y(
        n33673) );
  NAND2X1 U28086 ( .A(n33675), .B(n33676), .Y(n31896) );
  AOI22X1 U28087 ( .A(n30323), .B(n30285), .C(n30324), .D(n32310), .Y(n33676)
         );
  NAND2X1 U28088 ( .A(n33677), .B(n33678), .Y(n32310) );
  AOI22X1 U28089 ( .A(reg_A[57]), .B(n30846), .C(n30212), .D(reg_A[58]), .Y(
        n33678) );
  AOI22X1 U28090 ( .A(reg_A[59]), .B(n29987), .C(n30847), .D(reg_A[60]), .Y(
        n33677) );
  OAI21X1 U28091 ( .A(n30038), .B(n30007), .C(n33679), .Y(n30285) );
  AOI22X1 U28092 ( .A(reg_A[61]), .B(n30846), .C(n30212), .D(reg_A[62]), .Y(
        n33679) );
  INVX1 U28093 ( .A(reg_A[63]), .Y(n30007) );
  AOI22X1 U28094 ( .A(n30325), .B(n32723), .C(n30326), .D(n32725), .Y(n33675)
         );
  NAND2X1 U28095 ( .A(n33680), .B(n33681), .Y(n32725) );
  AOI22X1 U28096 ( .A(reg_A[53]), .B(n30846), .C(n30212), .D(reg_A[54]), .Y(
        n33681) );
  AOI22X1 U28097 ( .A(reg_A[55]), .B(n29987), .C(n30847), .D(reg_A[56]), .Y(
        n33680) );
  NAND2X1 U28098 ( .A(n33682), .B(n33683), .Y(n32723) );
  AOI22X1 U28099 ( .A(reg_A[49]), .B(n30846), .C(n30212), .D(reg_A[50]), .Y(
        n33683) );
  AOI22X1 U28100 ( .A(reg_A[51]), .B(n29987), .C(n30847), .D(reg_A[52]), .Y(
        n33682) );
  AOI22X1 U28101 ( .A(n33497), .B(reg_A[34]), .C(n33498), .D(reg_A[33]), .Y(
        n33671) );
  INVX1 U28102 ( .A(n33612), .Y(n33498) );
  INVX1 U28103 ( .A(n32765), .Y(n33497) );
  NAND2X1 U28104 ( .A(n33684), .B(n33685), .Y(n33669) );
  AOI22X1 U28105 ( .A(n33686), .B(reg_A[35]), .C(n33164), .D(n30847), .Y(
        n33685) );
  NOR2X1 U28106 ( .A(n30058), .B(n29976), .Y(n33164) );
  NOR2X1 U28107 ( .A(n30038), .B(n29976), .Y(n33686) );
  AOI22X1 U28108 ( .A(n32420), .B(n33238), .C(n32724), .D(n32377), .Y(n33684)
         );
  NAND2X1 U28109 ( .A(n33687), .B(n33688), .Y(n32377) );
  AOI22X1 U28110 ( .A(reg_A[45]), .B(n30846), .C(n30212), .D(reg_A[46]), .Y(
        n33688) );
  AOI22X1 U28111 ( .A(reg_A[47]), .B(n29987), .C(n30847), .D(reg_A[48]), .Y(
        n33687) );
  NAND2X1 U28112 ( .A(n33689), .B(n33690), .Y(n33238) );
  AOI22X1 U28113 ( .A(reg_A[37]), .B(n30846), .C(n30212), .D(reg_A[38]), .Y(
        n33690) );
  AOI22X1 U28114 ( .A(reg_A[39]), .B(n29987), .C(n30847), .D(reg_A[40]), .Y(
        n33689) );
  AND2X1 U28115 ( .A(n33691), .B(n33692), .Y(n33232) );
  AOI22X1 U28116 ( .A(n32299), .B(reg_A[39]), .C(n32109), .D(reg_A[38]), .Y(
        n33692) );
  AOI22X1 U28117 ( .A(n32357), .B(reg_A[40]), .C(n32110), .D(reg_A[37]), .Y(
        n33691) );
  OAI21X1 U28118 ( .A(n32315), .B(n32126), .C(n33693), .Y(n33666) );
  AOI22X1 U28119 ( .A(n32129), .B(n32716), .C(n33464), .D(n33234), .Y(n33693)
         );
  OAI21X1 U28120 ( .A(n30057), .B(n33619), .C(n33694), .Y(n33234) );
  AOI22X1 U28121 ( .A(n33695), .B(reg_A[39]), .C(n33076), .D(reg_A[38]), .Y(
        n33694) );
  INVX1 U28122 ( .A(n33662), .Y(n33464) );
  NAND2X1 U28123 ( .A(n33696), .B(n33697), .Y(n32716) );
  AOI22X1 U28124 ( .A(n32299), .B(reg_A[43]), .C(n32109), .D(reg_A[42]), .Y(
        n33697) );
  AOI22X1 U28125 ( .A(n32357), .B(reg_A[44]), .C(n32110), .D(reg_A[41]), .Y(
        n33696) );
  INVX1 U28126 ( .A(n33698), .Y(n32315) );
  OAI21X1 U28127 ( .A(n30066), .B(n32134), .C(n33699), .Y(n33698) );
  AOI22X1 U28128 ( .A(n32299), .B(reg_A[47]), .C(n32109), .D(reg_A[46]), .Y(
        n33699) );
  AOI22X1 U28129 ( .A(reg_A[35]), .B(n33457), .C(reg_A[34]), .D(n33452), .Y(
        n33664) );
  AOI22X1 U28130 ( .A(reg_A[36]), .B(n33453), .C(reg_A[33]), .D(n33551), .Y(
        n33663) );
  NAND3X1 U28131 ( .A(n33700), .B(n33701), .C(n33702), .Y(result[32]) );
  NOR2X1 U28132 ( .A(n33703), .B(n33704), .Y(n33702) );
  OAI22X1 U28133 ( .A(n25717), .B(n30394), .C(n25718), .D(n30393), .Y(n33704)
         );
  OAI21X1 U28134 ( .A(n25719), .B(n30170), .C(n33705), .Y(n33703) );
  AOI22X1 U28135 ( .A(n25721), .B(reg_A[16]), .C(reg_A[36]), .D(n25722), .Y(
        n33705) );
  AOI21X1 U28136 ( .A(n26928), .B(n33706), .C(n33707), .Y(n33701) );
  OAI21X1 U28137 ( .A(n33708), .B(n30395), .C(n33709), .Y(n33707) );
  OAI21X1 U28138 ( .A(n33710), .B(n33711), .C(n25730), .Y(n33709) );
  NAND3X1 U28139 ( .A(n33712), .B(n33713), .C(n33714), .Y(n33711) );
  NOR2X1 U28140 ( .A(n33715), .B(n33716), .Y(n33714) );
  OAI22X1 U28141 ( .A(n25736), .B(n30395), .C(n25737), .D(n30066), .Y(n33716)
         );
  OAI22X1 U28142 ( .A(n25738), .B(n30067), .C(n25739), .D(n30068), .Y(n33715)
         );
  AOI22X1 U28143 ( .A(reg_A[40]), .B(n25615), .C(reg_A[43]), .D(n25616), .Y(
        n33713) );
  AOI22X1 U28144 ( .A(reg_A[42]), .B(n25607), .C(reg_A[46]), .D(n25608), .Y(
        n33712) );
  NAND3X1 U28145 ( .A(n33717), .B(n33718), .C(n33719), .Y(n33710) );
  NOR2X1 U28146 ( .A(n33720), .B(n33721), .Y(n33719) );
  OAI22X1 U28147 ( .A(n25061), .B(n30060), .C(n25746), .D(n30394), .Y(n33721)
         );
  OAI22X1 U28148 ( .A(n25747), .B(n30393), .C(n25748), .D(n30170), .Y(n33720)
         );
  AOI22X1 U28149 ( .A(reg_A[39]), .B(n25613), .C(reg_A[36]), .D(n25749), .Y(
        n33718) );
  AOI22X1 U28150 ( .A(reg_A[37]), .B(n25750), .C(reg_A[41]), .D(n25614), .Y(
        n33717) );
  NOR2X1 U28151 ( .A(n29881), .B(n33722), .Y(n33708) );
  OAI22X1 U28152 ( .A(n33450), .B(n25697), .C(n26610), .D(n33612), .Y(n33722)
         );
  NAND3X1 U28153 ( .A(n25795), .B(n25032), .C(n25789), .Y(n29881) );
  AOI21X1 U28154 ( .A(n26801), .B(n30910), .C(n33723), .Y(n25789) );
  OAI21X1 U28155 ( .A(n33724), .B(n33394), .C(n33358), .Y(n33723) );
  OAI21X1 U28156 ( .A(n26944), .B(n30057), .C(n33725), .Y(n33706) );
  AOI22X1 U28157 ( .A(reg_A[38]), .B(n26010), .C(reg_A[39]), .D(n26002), .Y(
        n33725) );
  INVX1 U28158 ( .A(reg_A[37]), .Y(n30057) );
  AOI22X1 U28159 ( .A(n25310), .B(n33726), .C(n25382), .D(n33727), .Y(n33700)
         );
  NAND3X1 U28160 ( .A(n33728), .B(n33729), .C(n33730), .Y(n33727) );
  NOR2X1 U28161 ( .A(n33731), .B(n33732), .Y(n33730) );
  OAI22X1 U28162 ( .A(n33336), .B(n33339), .C(n32892), .D(n32126), .Y(n33732)
         );
  NAND3X1 U28163 ( .A(reg_B[45]), .B(n25604), .C(reg_B[44]), .Y(n32126) );
  INVX1 U28164 ( .A(n32478), .Y(n32892) );
  NAND2X1 U28165 ( .A(n33733), .B(n33734), .Y(n32478) );
  AOI22X1 U28166 ( .A(n32299), .B(reg_A[46]), .C(n32109), .D(reg_A[45]), .Y(
        n33734) );
  AOI22X1 U28167 ( .A(n32357), .B(reg_A[47]), .C(n32110), .D(reg_A[44]), .Y(
        n33733) );
  NAND2X1 U28168 ( .A(n32260), .B(n25604), .Y(n33339) );
  INVX1 U28169 ( .A(n32416), .Y(n32260) );
  NAND2X1 U28170 ( .A(reg_B[45]), .B(n32635), .Y(n32416) );
  AND2X1 U28171 ( .A(n33735), .B(n33736), .Y(n33336) );
  AOI22X1 U28172 ( .A(n32299), .B(reg_A[38]), .C(n32109), .D(reg_A[37]), .Y(
        n33736) );
  AOI22X1 U28173 ( .A(n32357), .B(reg_A[39]), .C(n32110), .D(reg_A[36]), .Y(
        n33735) );
  OAI21X1 U28174 ( .A(n33337), .B(n33662), .C(n33737), .Y(n33731) );
  AOI22X1 U28175 ( .A(n32129), .B(n33340), .C(reg_A[34]), .D(n33457), .Y(
        n33737) );
  OAI22X1 U28176 ( .A(n32066), .B(n33116), .C(n33338), .D(n33738), .Y(n33457)
         );
  NAND2X1 U28177 ( .A(n33739), .B(n33740), .Y(n33340) );
  AOI22X1 U28178 ( .A(n32299), .B(reg_A[42]), .C(n32109), .D(reg_A[41]), .Y(
        n33740) );
  INVX1 U28179 ( .A(n32253), .Y(n32109) );
  INVX1 U28180 ( .A(n32066), .Y(n32299) );
  NAND2X1 U28181 ( .A(reg_B[46]), .B(n32229), .Y(n32066) );
  AOI22X1 U28182 ( .A(n32357), .B(reg_A[43]), .C(n32110), .D(reg_A[40]), .Y(
        n33739) );
  INVX1 U28183 ( .A(n32134), .Y(n32110) );
  INVX1 U28184 ( .A(n32240), .Y(n32357) );
  INVX1 U28185 ( .A(n33019), .Y(n32129) );
  NAND2X1 U28186 ( .A(n32147), .B(n25604), .Y(n33019) );
  INVX1 U28187 ( .A(n32228), .Y(n32147) );
  NAND2X1 U28188 ( .A(reg_B[44]), .B(n32233), .Y(n32228) );
  NAND2X1 U28189 ( .A(reg_B[37]), .B(n25589), .Y(n33662) );
  AND2X1 U28190 ( .A(n33741), .B(n33742), .Y(n33337) );
  AOI22X1 U28191 ( .A(n33695), .B(reg_A[38]), .C(n33426), .D(reg_A[39]), .Y(
        n33742) );
  INVX1 U28192 ( .A(n33743), .Y(n33426) );
  INVX1 U28193 ( .A(n33738), .Y(n33695) );
  NAND2X1 U28194 ( .A(reg_B[38]), .B(n33176), .Y(n33738) );
  AOI22X1 U28195 ( .A(n33076), .B(reg_A[37]), .C(n33075), .D(reg_A[36]), .Y(
        n33741) );
  INVX1 U28196 ( .A(n33619), .Y(n33075) );
  AOI22X1 U28197 ( .A(reg_A[33]), .B(n33452), .C(reg_A[35]), .D(n33453), .Y(
        n33729) );
  OAI22X1 U28198 ( .A(n32240), .B(n33116), .C(n33338), .D(n33743), .Y(n33453)
         );
  NAND2X1 U28199 ( .A(reg_B[39]), .B(reg_B[38]), .Y(n33743) );
  NAND2X1 U28200 ( .A(reg_B[46]), .B(reg_B[47]), .Y(n32240) );
  OAI21X1 U28201 ( .A(n32253), .B(n33116), .C(n33120), .Y(n33452) );
  NAND2X1 U28202 ( .A(n33235), .B(n33076), .Y(n33120) );
  NOR2X1 U28203 ( .A(n33176), .B(reg_B[38]), .Y(n33076) );
  INVX1 U28204 ( .A(n33338), .Y(n33235) );
  NAND2X1 U28205 ( .A(reg_B[47]), .B(n32334), .Y(n32253) );
  AOI22X1 U28206 ( .A(n25097), .B(n33744), .C(reg_A[32]), .D(n33551), .Y(
        n33728) );
  INVX1 U28207 ( .A(n33450), .Y(n33551) );
  NOR2X1 U28208 ( .A(n33350), .B(n33130), .Y(n33450) );
  NOR2X1 U28209 ( .A(n33338), .B(n33619), .Y(n33130) );
  NAND2X1 U28210 ( .A(n33176), .B(n33071), .Y(n33619) );
  INVX1 U28211 ( .A(reg_B[38]), .Y(n33071) );
  INVX1 U28212 ( .A(reg_B[39]), .Y(n33176) );
  NAND2X1 U28213 ( .A(n25029), .B(n33079), .Y(n33338) );
  INVX1 U28214 ( .A(reg_B[37]), .Y(n33079) );
  NOR2X1 U28215 ( .A(n33116), .B(n32134), .Y(n33350) );
  NAND2X1 U28216 ( .A(n32334), .B(n32229), .Y(n32134) );
  INVX1 U28217 ( .A(reg_B[47]), .Y(n32229) );
  INVX1 U28218 ( .A(reg_B[46]), .Y(n32334) );
  NAND2X1 U28219 ( .A(n32261), .B(n25604), .Y(n33116) );
  INVX1 U28220 ( .A(n32371), .Y(n32261) );
  NAND2X1 U28221 ( .A(n32635), .B(n32233), .Y(n32371) );
  INVX1 U28222 ( .A(reg_B[45]), .Y(n32233) );
  INVX1 U28223 ( .A(reg_B[44]), .Y(n32635) );
  NAND3X1 U28224 ( .A(n33745), .B(n33746), .C(n33747), .Y(n33744) );
  NOR2X1 U28225 ( .A(n33748), .B(n33749), .Y(n33747) );
  OAI22X1 U28226 ( .A(n30395), .B(n33612), .C(n30170), .D(n32765), .Y(n33749)
         );
  NAND2X1 U28227 ( .A(n30492), .B(n30117), .Y(n32765) );
  INVX1 U28228 ( .A(n29978), .Y(n30492) );
  NAND2X1 U28229 ( .A(reg_B[63]), .B(n30024), .Y(n29978) );
  NAND2X1 U28230 ( .A(n30117), .B(n30107), .Y(n33612) );
  INVX1 U28231 ( .A(n30103), .Y(n30107) );
  NAND2X1 U28232 ( .A(n30024), .B(n30028), .Y(n30103) );
  NAND2X1 U28233 ( .A(n29973), .B(n30293), .Y(n30223) );
  OAI21X1 U28234 ( .A(n30210), .B(n33273), .C(n33308), .Y(n33748) );
  NAND3X1 U28235 ( .A(n30298), .B(n29987), .C(reg_A[34]), .Y(n33308) );
  NAND2X1 U28236 ( .A(reg_A[35]), .B(n30298), .Y(n33273) );
  INVX1 U28237 ( .A(n29976), .Y(n30298) );
  NAND2X1 U28238 ( .A(n30117), .B(n29973), .Y(n29976) );
  AOI22X1 U28239 ( .A(n32420), .B(n33376), .C(n32724), .D(n32497), .Y(n33746)
         );
  NAND2X1 U28240 ( .A(n33750), .B(n33751), .Y(n32497) );
  AOI22X1 U28241 ( .A(reg_A[44]), .B(n30846), .C(n30212), .D(reg_A[45]), .Y(
        n33751) );
  AOI22X1 U28242 ( .A(reg_A[46]), .B(n29987), .C(n30847), .D(reg_A[47]), .Y(
        n33750) );
  INVX1 U28243 ( .A(n32041), .Y(n32724) );
  NAND2X1 U28244 ( .A(n30208), .B(reg_B[61]), .Y(n32041) );
  NAND2X1 U28245 ( .A(n33752), .B(n33753), .Y(n33376) );
  AOI22X1 U28246 ( .A(reg_A[36]), .B(n30846), .C(n30212), .D(reg_A[37]), .Y(
        n33753) );
  AOI22X1 U28247 ( .A(reg_A[38]), .B(n29987), .C(n30847), .D(reg_A[39]), .Y(
        n33752) );
  INVX1 U28248 ( .A(n32045), .Y(n32420) );
  NAND2X1 U28249 ( .A(n30117), .B(reg_B[61]), .Y(n32045) );
  INVX1 U28250 ( .A(n29994), .Y(n30117) );
  NAND2X1 U28251 ( .A(n30341), .B(n30853), .Y(n29994) );
  AOI22X1 U28252 ( .A(reg_B[59]), .B(n32000), .C(n30039), .D(n33346), .Y(
        n33745) );
  NAND2X1 U28253 ( .A(n33754), .B(n33755), .Y(n33346) );
  AOI22X1 U28254 ( .A(reg_A[40]), .B(n30846), .C(n30212), .D(reg_A[41]), .Y(
        n33755) );
  AOI22X1 U28255 ( .A(reg_A[42]), .B(n29987), .C(n30847), .D(reg_A[43]), .Y(
        n33754) );
  INVX1 U28256 ( .A(n32043), .Y(n30039) );
  NAND2X1 U28257 ( .A(n30208), .B(n29973), .Y(n32043) );
  INVX1 U28258 ( .A(n30109), .Y(n30208) );
  NAND2X1 U28259 ( .A(reg_B[60]), .B(n30341), .Y(n30109) );
  INVX1 U28260 ( .A(reg_B[59]), .Y(n30341) );
  NAND2X1 U28261 ( .A(n33756), .B(n33757), .Y(n32000) );
  AOI22X1 U28262 ( .A(n30323), .B(n31044), .C(n30324), .D(n31032), .Y(n33757)
         );
  NAND2X1 U28263 ( .A(n33758), .B(n33759), .Y(n31032) );
  AOI22X1 U28264 ( .A(reg_A[56]), .B(n30846), .C(n30212), .D(reg_A[57]), .Y(
        n33759) );
  AOI22X1 U28265 ( .A(reg_A[58]), .B(n29987), .C(n30847), .D(reg_A[59]), .Y(
        n33758) );
  INVX1 U28266 ( .A(n30136), .Y(n30324) );
  NAND2X1 U28267 ( .A(reg_B[60]), .B(n29973), .Y(n30136) );
  NAND2X1 U28268 ( .A(n33760), .B(n33761), .Y(n31044) );
  AOI22X1 U28269 ( .A(reg_A[60]), .B(n30846), .C(n30212), .D(reg_A[61]), .Y(
        n33761) );
  AOI22X1 U28270 ( .A(reg_A[62]), .B(n29987), .C(n30847), .D(reg_A[63]), .Y(
        n33760) );
  NOR2X1 U28271 ( .A(n30853), .B(n29973), .Y(n30323) );
  AOI22X1 U28272 ( .A(n30325), .B(n33344), .C(n30326), .D(n32427), .Y(n33756)
         );
  NAND2X1 U28273 ( .A(n33762), .B(n33763), .Y(n32427) );
  AOI22X1 U28274 ( .A(reg_A[52]), .B(n30846), .C(n30212), .D(reg_A[53]), .Y(
        n33763) );
  AOI22X1 U28275 ( .A(reg_A[54]), .B(n29987), .C(n30847), .D(reg_A[55]), .Y(
        n33762) );
  INVX1 U28276 ( .A(n30220), .Y(n30326) );
  NAND2X1 U28277 ( .A(reg_B[61]), .B(n30853), .Y(n30220) );
  NAND2X1 U28278 ( .A(n33764), .B(n33765), .Y(n33344) );
  AOI22X1 U28279 ( .A(n30846), .B(reg_A[48]), .C(n30212), .D(reg_A[49]), .Y(
        n33765) );
  NAND2X1 U28280 ( .A(reg_B[63]), .B(n30293), .Y(n30320) );
  NAND2X1 U28281 ( .A(n30293), .B(n30028), .Y(n29970) );
  INVX1 U28282 ( .A(reg_B[62]), .Y(n30293) );
  AOI22X1 U28283 ( .A(reg_A[50]), .B(n29987), .C(n30847), .D(reg_A[51]), .Y(
        n33764) );
  NAND2X1 U28284 ( .A(reg_B[63]), .B(reg_B[62]), .Y(n30210) );
  NAND2X1 U28285 ( .A(reg_B[62]), .B(n30028), .Y(n30038) );
  INVX1 U28286 ( .A(reg_B[63]), .Y(n30028) );
  INVX1 U28287 ( .A(n29975), .Y(n30325) );
  NAND2X1 U28288 ( .A(n30853), .B(n29973), .Y(n29975) );
  INVX1 U28289 ( .A(reg_B[61]), .Y(n29973) );
  INVX1 U28290 ( .A(reg_B[60]), .Y(n30853) );
  NAND2X1 U28291 ( .A(n33766), .B(n33767), .Y(n33726) );
  NOR2X1 U28292 ( .A(n33768), .B(n33769), .Y(n33767) );
  NAND3X1 U28293 ( .A(n33770), .B(n33771), .C(n33772), .Y(n33769) );
  NOR2X1 U28294 ( .A(n33773), .B(n33774), .Y(n33772) );
  OAI22X1 U28295 ( .A(n25316), .B(n30219), .C(n25318), .D(n29984), .Y(n33774)
         );
  INVX1 U28296 ( .A(reg_A[59]), .Y(n29984) );
  INVX1 U28297 ( .A(reg_A[58]), .Y(n30219) );
  OAI22X1 U28298 ( .A(n25320), .B(n30254), .C(n25322), .D(n29990), .Y(n33773)
         );
  INVX1 U28299 ( .A(reg_A[57]), .Y(n29990) );
  INVX1 U28300 ( .A(reg_A[56]), .Y(n30254) );
  AOI22X1 U28301 ( .A(reg_A[62]), .B(n25631), .C(reg_A[63]), .D(n25764), .Y(
        n33771) );
  AOI22X1 U28302 ( .A(reg_A[60]), .B(n25324), .C(reg_A[61]), .D(n25765), .Y(
        n33770) );
  NAND3X1 U28303 ( .A(n33775), .B(n33776), .C(n33777), .Y(n33768) );
  NOR2X1 U28304 ( .A(n33778), .B(n33779), .Y(n33777) );
  OAI22X1 U28305 ( .A(n25331), .B(n30008), .C(n25243), .D(n30009), .Y(n33779)
         );
  OAI22X1 U28306 ( .A(n25334), .B(n29655), .C(n25336), .D(n30174), .Y(n33778)
         );
  AOI22X1 U28307 ( .A(reg_A[54]), .B(n25242), .C(reg_A[55]), .D(n25338), .Y(
        n33776) );
  AOI22X1 U28308 ( .A(reg_A[52]), .B(n25339), .C(reg_A[53]), .D(n25257), .Y(
        n33775) );
  NOR2X1 U28309 ( .A(n33780), .B(n33781), .Y(n33766) );
  NAND3X1 U28310 ( .A(n33782), .B(n33783), .C(n33784), .Y(n33781) );
  NOR2X1 U28311 ( .A(n33785), .B(n33786), .Y(n33784) );
  OAI22X1 U28312 ( .A(n25043), .B(n30395), .C(n25039), .D(n30066), .Y(n33786)
         );
  OAI22X1 U28313 ( .A(n25064), .B(n30067), .C(n25065), .D(n30068), .Y(n33785)
         );
  AOI22X1 U28314 ( .A(reg_A[40]), .B(n25124), .C(reg_A[43]), .D(n25222), .Y(
        n33783) );
  AOI22X1 U28315 ( .A(reg_A[42]), .B(n25637), .C(reg_A[46]), .D(n25234), .Y(
        n33782) );
  NAND3X1 U28316 ( .A(n33787), .B(n33788), .C(n33789), .Y(n33780) );
  NOR2X1 U28317 ( .A(n33790), .B(n33791), .Y(n33789) );
  OAI22X1 U28318 ( .A(n25033), .B(n30060), .C(n25133), .D(n30394), .Y(n33791)
         );
  OAI22X1 U28319 ( .A(n25041), .B(n30393), .C(n25042), .D(n30170), .Y(n33790)
         );
  AOI22X1 U28320 ( .A(reg_A[39]), .B(n25628), .C(reg_A[36]), .D(n25068), .Y(
        n33788) );
  AOI22X1 U28321 ( .A(reg_A[37]), .B(n25123), .C(reg_A[41]), .D(n25629), .Y(
        n33787) );
  NAND3X1 U28322 ( .A(n33792), .B(n33793), .C(n33794), .Y(result[31]) );
  NOR2X1 U28323 ( .A(n33795), .B(n33796), .Y(n33794) );
  NAND3X1 U28324 ( .A(n33797), .B(n33798), .C(n33799), .Y(n33796) );
  AOI21X1 U28325 ( .A(n33800), .B(n25900), .C(n33801), .Y(n33799) );
  OAI22X1 U28326 ( .A(n29958), .B(n33802), .C(n25939), .D(n33803), .Y(n33801)
         );
  OAI21X1 U28327 ( .A(n33804), .B(n33805), .C(n33806), .Y(n33798) );
  OAI22X1 U28328 ( .A(n33807), .B(n26996), .C(n28105), .D(n33808), .Y(n33805)
         );
  AOI22X1 U28329 ( .A(n33809), .B(n33810), .C(n25840), .D(n33811), .Y(n33797)
         );
  NAND2X1 U28330 ( .A(n33812), .B(n33813), .Y(n33811) );
  NOR2X1 U28331 ( .A(n33814), .B(n33815), .Y(n33813) );
  NAND3X1 U28332 ( .A(n33816), .B(n33817), .C(n33818), .Y(n33815) );
  NOR2X1 U28333 ( .A(n33819), .B(n33820), .Y(n33818) );
  OAI22X1 U28334 ( .A(n25130), .B(n25499), .C(n26742), .D(n25852), .Y(n33820)
         );
  OAI22X1 U28335 ( .A(n25177), .B(n25854), .C(n29265), .D(n25316), .Y(n33819)
         );
  AOI22X1 U28336 ( .A(reg_A[10]), .B(n25257), .C(n25857), .D(reg_A[6]), .Y(
        n33817) );
  AOI22X1 U28337 ( .A(n25647), .B(reg_A[7]), .C(n25648), .D(reg_A[4]), .Y(
        n33816) );
  NAND3X1 U28338 ( .A(n33821), .B(n33822), .C(n33823), .Y(n33814) );
  NOR2X1 U28339 ( .A(n33824), .B(n33825), .Y(n33823) );
  OAI22X1 U28340 ( .A(n25038), .B(n25255), .C(n25334), .D(n29279), .Y(n33825)
         );
  OAI21X1 U28341 ( .A(n25047), .B(n25208), .C(n33826), .Y(n33824) );
  AOI22X1 U28342 ( .A(reg_A[13]), .B(n25241), .C(n25242), .D(reg_A[9]), .Y(
        n33822) );
  AOI22X1 U28343 ( .A(n25338), .B(reg_A[8]), .C(reg_A[11]), .D(n25339), .Y(
        n33821) );
  NOR2X1 U28344 ( .A(n33827), .B(n33828), .Y(n33812) );
  NAND3X1 U28345 ( .A(n33829), .B(n33830), .C(n33831), .Y(n33828) );
  NOR2X1 U28346 ( .A(n33832), .B(n33833), .Y(n33831) );
  OAI22X1 U28347 ( .A(n27954), .B(n25228), .C(n25224), .D(n25229), .Y(n33833)
         );
  OAI22X1 U28348 ( .A(n25220), .B(n25231), .C(n25250), .D(n25482), .Y(n33832)
         );
  AOI22X1 U28349 ( .A(reg_A[22]), .B(n25629), .C(reg_A[20]), .D(n25222), .Y(
        n33830) );
  AOI22X1 U28350 ( .A(reg_A[21]), .B(n25637), .C(n25234), .D(reg_A[17]), .Y(
        n33829) );
  NAND3X1 U28351 ( .A(n33834), .B(n33835), .C(n33836), .Y(n33827) );
  NOR2X1 U28352 ( .A(n33837), .B(n33838), .Y(n33836) );
  OAI22X1 U28353 ( .A(n25239), .B(n25133), .C(n25244), .D(n25254), .Y(n33838)
         );
  OAI22X1 U28354 ( .A(n29286), .B(n25784), .C(n25128), .D(n25498), .Y(n33837)
         );
  AOI22X1 U28355 ( .A(n25253), .B(reg_A[25]), .C(reg_A[24]), .D(n25628), .Y(
        n33835) );
  AOI22X1 U28356 ( .A(n25075), .B(reg_A[27]), .C(n25123), .D(reg_A[26]), .Y(
        n33834) );
  OAI21X1 U28357 ( .A(n25032), .B(n33839), .C(n33840), .Y(n33810) );
  AOI22X1 U28358 ( .A(n26504), .B(n33841), .C(n30616), .D(n33842), .Y(n33840)
         );
  NAND3X1 U28359 ( .A(n33843), .B(n33844), .C(n33845), .Y(n33795) );
  AOI21X1 U28360 ( .A(n26186), .B(n33846), .C(n33847), .Y(n33845) );
  OAI21X1 U28361 ( .A(n33848), .B(n33849), .C(n33850), .Y(n33847) );
  OAI21X1 U28362 ( .A(n33851), .B(n33852), .C(n25918), .Y(n33850) );
  NAND3X1 U28363 ( .A(n33853), .B(n33854), .C(n33855), .Y(n33852) );
  NOR2X1 U28364 ( .A(n33856), .B(n33857), .Y(n33855) );
  OAI22X1 U28365 ( .A(n25736), .B(n27954), .C(n25224), .D(n25737), .Y(n33857)
         );
  OAI22X1 U28366 ( .A(n25220), .B(n25738), .C(n25250), .D(n25739), .Y(n33856)
         );
  AOI22X1 U28367 ( .A(reg_A[23]), .B(n25615), .C(reg_A[20]), .D(n25616), .Y(
        n33854) );
  AOI22X1 U28368 ( .A(reg_A[21]), .B(n25607), .C(n25608), .D(reg_A[17]), .Y(
        n33853) );
  NAND3X1 U28369 ( .A(n33858), .B(n33859), .C(n33860), .Y(n33851) );
  NOR2X1 U28370 ( .A(n33861), .B(n33862), .Y(n33860) );
  OAI22X1 U28371 ( .A(n25061), .B(n27960), .C(n25746), .D(n25239), .Y(n33862)
         );
  OAI22X1 U28372 ( .A(n25747), .B(n25244), .C(n25748), .D(n29286), .Y(n33861)
         );
  AOI22X1 U28373 ( .A(reg_A[24]), .B(n25613), .C(n25749), .D(reg_A[27]), .Y(
        n33859) );
  AOI22X1 U28374 ( .A(n25750), .B(reg_A[26]), .C(reg_A[22]), .D(n25614), .Y(
        n33858) );
  NAND2X1 U28375 ( .A(n33863), .B(n25188), .Y(n33849) );
  NAND2X1 U28376 ( .A(reg_B[28]), .B(n32934), .Y(n33848) );
  OAI22X1 U28377 ( .A(n33864), .B(n33865), .C(n29305), .D(n33866), .Y(n33846)
         );
  MUX2X1 U28378 ( .B(reg_A[29]), .A(reg_A[25]), .S(reg_B[29]), .Y(n33866) );
  INVX1 U28379 ( .A(n33867), .Y(n33864) );
  NAND2X1 U28380 ( .A(n33868), .B(n28138), .Y(n33844) );
  AOI22X1 U28381 ( .A(reg_A[27]), .B(n33869), .C(n33870), .D(n25910), .Y(
        n33843) );
  INVX1 U28382 ( .A(n33871), .Y(n33870) );
  OAI21X1 U28383 ( .A(n33872), .B(n33873), .C(n28122), .Y(n33869) );
  NAND2X1 U28384 ( .A(n25170), .B(n33874), .Y(n33873) );
  NOR2X1 U28385 ( .A(n33875), .B(n33876), .Y(n33793) );
  OAI21X1 U28386 ( .A(n27961), .B(n32117), .C(n33877), .Y(n33876) );
  AOI22X1 U28387 ( .A(reg_A[31]), .B(n25952), .C(reg_B[30]), .D(n33878), .Y(
        n33877) );
  OAI21X1 U28388 ( .A(n25043), .B(n25835), .C(n30195), .Y(n25952) );
  INVX1 U28389 ( .A(n26044), .Y(n30195) );
  OAI21X1 U28390 ( .A(n33879), .B(n29286), .C(n33880), .Y(n33875) );
  AOI21X1 U28391 ( .A(n33881), .B(n27676), .C(n33882), .Y(n33880) );
  AOI21X1 U28392 ( .A(n33883), .B(n33884), .C(n25024), .Y(n33882) );
  AOI21X1 U28393 ( .A(n33885), .B(reg_B[31]), .C(n33886), .Y(n33884) );
  OAI21X1 U28394 ( .A(n33887), .B(n33888), .C(n33889), .Y(n33886) );
  NAND2X1 U28395 ( .A(n33890), .B(reg_B[27]), .Y(n33888) );
  INVX1 U28396 ( .A(n33891), .Y(n33885) );
  AOI22X1 U28397 ( .A(n33892), .B(n25258), .C(n33806), .D(n32933), .Y(n33883)
         );
  INVX1 U28398 ( .A(n33893), .Y(n33892) );
  INVX1 U28399 ( .A(n33894), .Y(n33879) );
  NOR2X1 U28400 ( .A(n33895), .B(n33896), .Y(n33792) );
  OAI21X1 U28401 ( .A(n33897), .B(n25697), .C(n33898), .Y(n33896) );
  OAI21X1 U28402 ( .A(n33899), .B(n33900), .C(n25999), .Y(n33898) );
  NAND2X1 U28403 ( .A(n33901), .B(n33902), .Y(n33900) );
  AOI22X1 U28404 ( .A(reg_A[24]), .B(n26002), .C(n26003), .D(reg_A[27]), .Y(
        n33902) );
  AOI22X1 U28405 ( .A(n25751), .B(reg_A[26]), .C(reg_A[31]), .D(n26004), .Y(
        n33901) );
  NAND2X1 U28406 ( .A(n33903), .B(n33904), .Y(n33899) );
  AOI22X1 U28407 ( .A(reg_A[30]), .B(n26007), .C(reg_A[28]), .D(n26008), .Y(
        n33904) );
  AOI22X1 U28408 ( .A(reg_A[29]), .B(n26009), .C(reg_A[25]), .D(n26010), .Y(
        n33903) );
  AOI21X1 U28409 ( .A(n25604), .B(n33905), .C(n33906), .Y(n33897) );
  OAI21X1 U28410 ( .A(n33907), .B(n31806), .C(n33908), .Y(n33906) );
  OAI21X1 U28411 ( .A(n33909), .B(n33910), .C(n25044), .Y(n33908) );
  OAI22X1 U28412 ( .A(n27954), .B(n33911), .C(n33912), .D(n33872), .Y(n33910)
         );
  INVX1 U28413 ( .A(n33913), .Y(n33912) );
  OAI21X1 U28414 ( .A(n33914), .B(n33915), .C(n33916), .Y(n33909) );
  INVX1 U28415 ( .A(n33917), .Y(n33916) );
  OAI21X1 U28416 ( .A(n29305), .B(n33918), .C(n33889), .Y(n33917) );
  NAND3X1 U28417 ( .A(reg_A[23]), .B(n33919), .C(n33890), .Y(n33889) );
  AOI21X1 U28418 ( .A(n33920), .B(reg_B[29]), .C(n33921), .Y(n33918) );
  AOI22X1 U28419 ( .A(n33922), .B(reg_A[7]), .C(n33923), .D(reg_A[15]), .Y(
        n33914) );
  OAI21X1 U28420 ( .A(n33924), .B(n29305), .C(n33925), .Y(n33905) );
  AOI22X1 U28421 ( .A(reg_B[28]), .B(n33926), .C(reg_B[31]), .D(n33927), .Y(
        n33925) );
  OAI22X1 U28422 ( .A(n26714), .B(n33915), .C(n25220), .D(n33872), .Y(n33926)
         );
  OAI21X1 U28423 ( .A(n25994), .B(n33928), .C(n33929), .Y(n33895) );
  AOI22X1 U28424 ( .A(n33930), .B(n32116), .C(n33931), .D(n26260), .Y(n33929)
         );
  INVX1 U28425 ( .A(n33932), .Y(n33931) );
  NAND3X1 U28426 ( .A(n33933), .B(n33934), .C(n33935), .Y(result[30]) );
  AND2X1 U28427 ( .A(n33936), .B(n33937), .Y(n33935) );
  NOR2X1 U28428 ( .A(n33938), .B(n33939), .Y(n33937) );
  OAI21X1 U28429 ( .A(n33907), .B(n31828), .C(n33940), .Y(n33939) );
  INVX1 U28430 ( .A(n33941), .Y(n33940) );
  OAI22X1 U28431 ( .A(n33942), .B(n26145), .C(n25244), .D(n26163), .Y(n33941)
         );
  NOR2X1 U28432 ( .A(n33943), .B(n27183), .Y(n26163) );
  AOI21X1 U28433 ( .A(n33944), .B(n33809), .C(n33945), .Y(n33907) );
  INVX1 U28434 ( .A(n33946), .Y(n33945) );
  AOI22X1 U28435 ( .A(n32934), .B(n33947), .C(reg_B[30]), .D(n33948), .Y(
        n33946) );
  NAND2X1 U28436 ( .A(n33949), .B(n33950), .Y(n33947) );
  AOI22X1 U28437 ( .A(n33922), .B(reg_A[6]), .C(n33923), .D(reg_A[14]), .Y(
        n33950) );
  AOI22X1 U28438 ( .A(reg_A[22]), .B(n33919), .C(reg_A[30]), .D(n32933), .Y(
        n33949) );
  OAI21X1 U28439 ( .A(n33951), .B(n29286), .C(n33952), .Y(n33938) );
  AOI22X1 U28440 ( .A(n26267), .B(n33953), .C(n25188), .D(n33954), .Y(n33952)
         );
  OAI22X1 U28441 ( .A(n33955), .B(n33956), .C(n33957), .D(n33958), .Y(n33954)
         );
  OAI22X1 U28442 ( .A(n33959), .B(n25264), .C(n33924), .D(n26758), .Y(n33953)
         );
  AOI21X1 U28443 ( .A(n33890), .B(n33804), .C(n26044), .Y(n33951) );
  OAI21X1 U28444 ( .A(n26943), .B(n29998), .C(n33960), .Y(n26044) );
  NOR2X1 U28445 ( .A(n26179), .B(n33961), .Y(n33960) );
  NOR2X1 U28446 ( .A(n33962), .B(n33963), .Y(n33936) );
  OAI22X1 U28447 ( .A(n33964), .B(n33891), .C(n27954), .D(n26136), .Y(n33963)
         );
  OAI21X1 U28448 ( .A(n33965), .B(n33966), .C(n33967), .Y(n33891) );
  AOI22X1 U28449 ( .A(n32934), .B(n33968), .C(reg_B[30]), .D(n33969), .Y(
        n33967) );
  OAI21X1 U28450 ( .A(reg_A[30]), .B(n33807), .C(n33970), .Y(n33968) );
  AOI22X1 U28451 ( .A(reg_B[27]), .B(n33971), .C(n33919), .D(n25230), .Y(
        n33970) );
  INVX1 U28452 ( .A(n33972), .Y(n33965) );
  OAI21X1 U28453 ( .A(n26421), .B(n33973), .C(n33974), .Y(n33962) );
  AOI22X1 U28454 ( .A(reg_A[29]), .B(n33894), .C(reg_A[27]), .D(n26161), .Y(
        n33974) );
  NAND2X1 U28455 ( .A(n26205), .B(n33975), .Y(n26161) );
  OAI21X1 U28456 ( .A(n33976), .B(n33977), .C(n26122), .Y(n33894) );
  INVX1 U28457 ( .A(n26016), .Y(n26122) );
  OAI21X1 U28458 ( .A(n27925), .B(n29998), .C(n33978), .Y(n26016) );
  NOR2X1 U28459 ( .A(n33979), .B(n33980), .Y(n33934) );
  OAI22X1 U28460 ( .A(n26012), .B(n33981), .C(n26525), .D(n33932), .Y(n33980)
         );
  OAI21X1 U28461 ( .A(n33982), .B(n26030), .C(n33983), .Y(n33932) );
  AOI22X1 U28462 ( .A(n26032), .B(n33984), .C(n25025), .D(n33985), .Y(n33983)
         );
  OAI21X1 U28463 ( .A(reg_A[30]), .B(n25063), .C(n33986), .Y(n33984) );
  AOI22X1 U28464 ( .A(n26038), .B(n25230), .C(reg_B[0]), .D(n33987), .Y(n33986) );
  OAI21X1 U28465 ( .A(n30226), .B(n27961), .C(n33988), .Y(n33979) );
  AOI22X1 U28466 ( .A(reg_A[24]), .B(n26043), .C(reg_A[25]), .D(n28282), .Y(
        n33988) );
  NOR2X1 U28467 ( .A(n33989), .B(n33990), .Y(n33933) );
  OAI21X1 U28468 ( .A(n29255), .B(n33991), .C(n33992), .Y(n33990) );
  MUX2X1 U28469 ( .B(n33993), .A(n33994), .S(reg_B[31]), .Y(n33992) );
  NAND3X1 U28470 ( .A(n33995), .B(n33996), .C(n33997), .Y(n33994) );
  AOI22X1 U28471 ( .A(n26186), .B(n33998), .C(n33999), .D(n25932), .Y(n33997)
         );
  NAND3X1 U28472 ( .A(reg_A[27]), .B(n33804), .C(n34000), .Y(n33996) );
  NAND3X1 U28473 ( .A(reg_A[25]), .B(n26504), .C(n33809), .Y(n33995) );
  NAND2X1 U28474 ( .A(n34001), .B(n34002), .Y(n33993) );
  AOI22X1 U28475 ( .A(n34003), .B(n34000), .C(n34004), .D(n33809), .Y(n34002)
         );
  NOR2X1 U28476 ( .A(n33976), .B(n25244), .Y(n34003) );
  INVX1 U28477 ( .A(n33804), .Y(n33976) );
  OAI21X1 U28478 ( .A(reg_B[28]), .B(n25794), .C(n25031), .Y(n33804) );
  AOI22X1 U28479 ( .A(n26186), .B(n33867), .C(n26267), .D(n33927), .Y(n34001)
         );
  NAND2X1 U28480 ( .A(n34005), .B(n34006), .Y(n33927) );
  MUX2X1 U28481 ( .B(n34007), .A(n34008), .S(reg_B[30]), .Y(n34006) );
  NOR2X1 U28482 ( .A(n27961), .B(n34009), .Y(n34007) );
  AOI22X1 U28483 ( .A(reg_B[28]), .B(n34010), .C(n34011), .D(reg_A[30]), .Y(
        n34005) );
  OAI22X1 U28484 ( .A(n34012), .B(n25230), .C(n25224), .D(n33966), .Y(n34010)
         );
  NAND2X1 U28485 ( .A(n34013), .B(n34014), .Y(n33867) );
  AOI22X1 U28486 ( .A(n34015), .B(reg_A[24]), .C(n34000), .D(reg_A[28]), .Y(
        n34014) );
  AOI22X1 U28487 ( .A(n33809), .B(reg_A[26]), .C(reg_A[30]), .D(n32934), .Y(
        n34013) );
  OAI21X1 U28488 ( .A(n34016), .B(n34017), .C(n34018), .Y(n33989) );
  AOI22X1 U28489 ( .A(n26045), .B(n34019), .C(n34020), .D(n34021), .Y(n34018)
         );
  NAND3X1 U28490 ( .A(n34022), .B(n34023), .C(n34024), .Y(n34019) );
  NOR2X1 U28491 ( .A(n34025), .B(n34026), .Y(n34024) );
  OAI22X1 U28492 ( .A(n25598), .B(n25244), .C(n25599), .D(n32918), .Y(n34026)
         );
  OAI21X1 U28493 ( .A(n25600), .B(n27960), .C(n34027), .Y(n34025) );
  OAI21X1 U28494 ( .A(n34028), .B(n34029), .C(n25604), .Y(n34027) );
  NAND2X1 U28495 ( .A(n34030), .B(n34031), .Y(n34029) );
  AOI22X1 U28496 ( .A(n25607), .B(reg_A[20]), .C(n25608), .D(reg_A[16]), .Y(
        n34031) );
  AOI22X1 U28497 ( .A(n25609), .B(reg_A[18]), .C(n25610), .D(reg_A[17]), .Y(
        n34030) );
  NAND2X1 U28498 ( .A(n34032), .B(n34033), .Y(n34028) );
  AOI22X1 U28499 ( .A(reg_A[23]), .B(n25613), .C(reg_A[21]), .D(n25614), .Y(
        n34033) );
  AOI22X1 U28500 ( .A(reg_A[22]), .B(n25615), .C(reg_A[19]), .D(n25616), .Y(
        n34032) );
  AOI21X1 U28501 ( .A(reg_A[29]), .B(n25617), .C(n34034), .Y(n34023) );
  OAI21X1 U28502 ( .A(n25619), .B(n29286), .C(n34035), .Y(n34034) );
  OAI21X1 U28503 ( .A(n34036), .B(n34037), .C(n25044), .Y(n34035) );
  NAND2X1 U28504 ( .A(n34038), .B(n34039), .Y(n34037) );
  NOR2X1 U28505 ( .A(n34040), .B(n34041), .Y(n34039) );
  OAI21X1 U28506 ( .A(n25034), .B(n25230), .C(n34042), .Y(n34041) );
  AOI22X1 U28507 ( .A(reg_A[23]), .B(n25628), .C(reg_A[21]), .D(n25629), .Y(
        n34042) );
  OAI21X1 U28508 ( .A(n25177), .B(n25498), .C(n34043), .Y(n34040) );
  AOI22X1 U28509 ( .A(n25631), .B(reg_A[0]), .C(n25324), .D(reg_A[2]), .Y(
        n34043) );
  NOR2X1 U28510 ( .A(n34044), .B(n34045), .Y(n34038) );
  OAI21X1 U28511 ( .A(n27953), .B(n25229), .C(n34046), .Y(n34045) );
  AOI22X1 U28512 ( .A(n25235), .B(reg_A[15]), .C(n25635), .D(reg_A[18]), .Y(
        n34046) );
  OAI21X1 U28513 ( .A(n25250), .B(n25475), .C(n34047), .Y(n34044) );
  AOI22X1 U28514 ( .A(reg_A[19]), .B(n25222), .C(n25637), .D(reg_A[20]), .Y(
        n34047) );
  NAND2X1 U28515 ( .A(n34048), .B(n34049), .Y(n34036) );
  NOR2X1 U28516 ( .A(n34050), .B(n34051), .Y(n34049) );
  OAI21X1 U28517 ( .A(n25132), .B(n25491), .C(n34052), .Y(n34051) );
  AOI22X1 U28518 ( .A(reg_A[12]), .B(n25241), .C(n25242), .D(reg_A[8]), .Y(
        n34052) );
  OAI21X1 U28519 ( .A(n25038), .B(n27967), .C(n34053), .Y(n34050) );
  AOI22X1 U28520 ( .A(reg_A[13]), .B(n25246), .C(reg_A[14]), .D(n25247), .Y(
        n34053) );
  NOR2X1 U28521 ( .A(n34054), .B(n34055), .Y(n34048) );
  OAI21X1 U28522 ( .A(n30569), .B(n25316), .C(n34056), .Y(n34055) );
  AOI22X1 U28523 ( .A(n25647), .B(reg_A[6]), .C(n25648), .D(reg_A[3]), .Y(
        n34056) );
  OAI21X1 U28524 ( .A(n29265), .B(n25322), .C(n34057), .Y(n34054) );
  AOI22X1 U28525 ( .A(reg_A[10]), .B(n25339), .C(n25257), .D(reg_A[9]), .Y(
        n34057) );
  AOI22X1 U28526 ( .A(reg_A[26]), .B(n25650), .C(reg_A[24]), .D(n25651), .Y(
        n34022) );
  NAND3X1 U28527 ( .A(n34058), .B(n34059), .C(n34060), .Y(result[2]) );
  NOR2X1 U28528 ( .A(n34061), .B(n34062), .Y(n34060) );
  NAND3X1 U28529 ( .A(n34063), .B(n34064), .C(n34065), .Y(n34062) );
  OAI21X1 U28530 ( .A(n34066), .B(n34067), .C(reg_A[0]), .Y(n34065) );
  OAI21X1 U28531 ( .A(n26032), .B(n26864), .C(n34068), .Y(n34067) );
  AOI21X1 U28532 ( .A(reg_B[30]), .B(n25932), .C(n34069), .Y(n34068) );
  AOI21X1 U28533 ( .A(n34070), .B(n33591), .C(n31658), .Y(n34069) );
  OR2X1 U28534 ( .A(n33394), .B(n26032), .Y(n33591) );
  NAND3X1 U28535 ( .A(n32940), .B(n29513), .C(n34071), .Y(n34066) );
  NAND2X1 U28536 ( .A(reg_B[6]), .B(n26504), .Y(n32940) );
  OAI21X1 U28537 ( .A(n34072), .B(n34073), .C(reg_A[1]), .Y(n34064) );
  OAI21X1 U28538 ( .A(n32947), .B(n33600), .C(n25566), .Y(n34073) );
  NAND2X1 U28539 ( .A(n29568), .B(n29565), .Y(n25566) );
  NOR2X1 U28540 ( .A(n25372), .B(n25170), .Y(n33600) );
  NOR2X1 U28541 ( .A(n25198), .B(n32950), .Y(n34072) );
  OAI21X1 U28542 ( .A(n34074), .B(n34075), .C(n25382), .Y(n34063) );
  OAI21X1 U28543 ( .A(n34076), .B(n29265), .C(n34077), .Y(n34075) );
  AOI22X1 U28544 ( .A(reg_A[4]), .B(n32998), .C(reg_A[3]), .D(n32999), .Y(
        n34077) );
  NAND2X1 U28545 ( .A(n34078), .B(n34079), .Y(n34074) );
  AOI22X1 U28546 ( .A(n32997), .B(n34080), .C(n28038), .D(n29232), .Y(n34079)
         );
  NAND2X1 U28547 ( .A(n34081), .B(n34082), .Y(n29232) );
  AOI22X1 U28548 ( .A(n26733), .B(reg_A[8]), .C(reg_A[7]), .D(n25172), .Y(
        n34082) );
  AOI22X1 U28549 ( .A(reg_A[9]), .B(n26734), .C(n25116), .D(reg_A[6]), .Y(
        n34081) );
  INVX1 U28550 ( .A(n29234), .Y(n34080) );
  AOI22X1 U28551 ( .A(reg_A[6]), .B(n27986), .C(reg_A[7]), .D(n28009), .Y(
        n29234) );
  AOI22X1 U28552 ( .A(n34083), .B(n29246), .C(n29245), .D(n29247), .Y(n34078)
         );
  NAND3X1 U28553 ( .A(n34084), .B(n32931), .C(n34085), .Y(n34061) );
  AOI22X1 U28554 ( .A(n30608), .B(n34086), .C(reg_A[2]), .D(n34087), .Y(n34085) );
  OAI21X1 U28555 ( .A(n34088), .B(n34089), .C(n34090), .Y(n34087) );
  NOR2X1 U28556 ( .A(n33602), .B(n26689), .Y(n34090) );
  INVX1 U28557 ( .A(n31788), .Y(n26689) );
  INVX1 U28558 ( .A(n25518), .Y(n33602) );
  NAND2X1 U28559 ( .A(n25284), .B(n29565), .Y(n25518) );
  INVX1 U28560 ( .A(n32961), .Y(n34086) );
  AOI22X1 U28561 ( .A(reg_A[0]), .B(n30613), .C(reg_A[2]), .D(n30612), .Y(
        n32961) );
  NOR2X1 U28562 ( .A(reg_B[5]), .B(reg_B[6]), .Y(n30612) );
  INVX1 U28563 ( .A(n30609), .Y(n30613) );
  NAND2X1 U28564 ( .A(reg_B[6]), .B(n31789), .Y(n30609) );
  INVX1 U28565 ( .A(n29319), .Y(n30608) );
  NAND2X1 U28566 ( .A(n26186), .B(n28041), .Y(n29319) );
  NAND3X1 U28567 ( .A(n32963), .B(n29302), .C(n26267), .Y(n34084) );
  OAI21X1 U28568 ( .A(n26742), .B(n25197), .C(n34091), .Y(n32963) );
  NAND3X1 U28569 ( .A(n31796), .B(n29256), .C(reg_A[2]), .Y(n34091) );
  INVX1 U28570 ( .A(n30551), .Y(n25197) );
  NOR2X1 U28571 ( .A(n29256), .B(n29304), .Y(n30551) );
  NOR2X1 U28572 ( .A(n34092), .B(n34093), .Y(n34059) );
  OAI22X1 U28573 ( .A(n25132), .B(n25652), .C(n26677), .D(n29782), .Y(n34093)
         );
  OAI22X1 U28574 ( .A(n29265), .B(n29765), .C(n30569), .D(n29766), .Y(n34092)
         );
  AOI21X1 U28575 ( .A(n26480), .B(n34094), .C(n34095), .Y(n34058) );
  OAI21X1 U28576 ( .A(n32967), .B(n31828), .C(n34096), .Y(n34095) );
  OAI21X1 U28577 ( .A(n34097), .B(n34098), .C(n25203), .Y(n34096) );
  NAND3X1 U28578 ( .A(n34099), .B(n34100), .C(n34101), .Y(n34098) );
  AOI21X1 U28579 ( .A(reg_A[2]), .B(n25434), .C(n34102), .Y(n34101) );
  OAI22X1 U28580 ( .A(n30569), .B(n25437), .C(n26677), .D(n25438), .Y(n34102)
         );
  AOI22X1 U28581 ( .A(n25439), .B(reg_A[12]), .C(n25440), .D(reg_A[8]), .Y(
        n34100) );
  AOI22X1 U28582 ( .A(reg_A[3]), .B(n25441), .C(n25442), .D(reg_A[5]), .Y(
        n34099) );
  NAND3X1 U28583 ( .A(n34103), .B(n34104), .C(n34105), .Y(n34097) );
  NOR2X1 U28584 ( .A(n34106), .B(n34107), .Y(n34105) );
  OAI22X1 U28585 ( .A(n25132), .B(n25449), .C(n25208), .D(n25451), .Y(n34107)
         );
  OAI21X1 U28586 ( .A(n29279), .B(n25453), .C(n34108), .Y(n34106) );
  OAI21X1 U28587 ( .A(n34109), .B(n34110), .C(n25044), .Y(n34108) );
  NAND3X1 U28588 ( .A(n34111), .B(n34112), .C(n34113), .Y(n34110) );
  NOR2X1 U28589 ( .A(n34114), .B(n34115), .Y(n34113) );
  OAI21X1 U28590 ( .A(n25128), .B(n25043), .C(n34116), .Y(n34115) );
  AOI22X1 U28591 ( .A(n25135), .B(reg_A[3]), .C(n25252), .D(reg_A[4]), .Y(
        n34116) );
  NAND2X1 U28592 ( .A(n34117), .B(n34118), .Y(n34114) );
  AOI22X1 U28593 ( .A(n25136), .B(reg_A[5]), .C(n25253), .D(reg_A[8]), .Y(
        n34118) );
  AOI22X1 U28594 ( .A(n25075), .B(reg_A[6]), .C(n25123), .D(reg_A[7]), .Y(
        n34117) );
  NOR2X1 U28595 ( .A(n34119), .B(n34120), .Y(n34112) );
  OAI22X1 U28596 ( .A(n25147), .B(n25467), .C(n25146), .D(n25129), .Y(n34120)
         );
  OAI22X1 U28597 ( .A(n25255), .B(n25219), .C(n27967), .D(n25223), .Y(n34119)
         );
  NOR2X1 U28598 ( .A(n34121), .B(n34122), .Y(n34111) );
  OAI22X1 U28599 ( .A(n25208), .B(n25231), .C(n25206), .D(n25473), .Y(n34122)
         );
  OAI22X1 U28600 ( .A(n29279), .B(n25229), .C(n25250), .D(n25475), .Y(n34121)
         );
  NAND3X1 U28601 ( .A(n34123), .B(n34124), .C(n34125), .Y(n34109) );
  NOR2X1 U28602 ( .A(n34126), .B(n34127), .Y(n34125) );
  OAI21X1 U28603 ( .A(n27953), .B(n25482), .C(n34128), .Y(n34127) );
  AOI22X1 U28604 ( .A(reg_A[19]), .B(n25246), .C(reg_A[18]), .D(n25247), .Y(
        n34128) );
  NAND2X1 U28605 ( .A(n34129), .B(n34130), .Y(n34126) );
  AOI22X1 U28606 ( .A(reg_A[21]), .B(n25487), .C(reg_A[20]), .D(n25241), .Y(
        n34130) );
  AOI22X1 U28607 ( .A(reg_A[22]), .B(n25339), .C(reg_A[23]), .D(n25257), .Y(
        n34129) );
  NOR2X1 U28608 ( .A(n34131), .B(n34132), .Y(n34124) );
  OAI22X1 U28609 ( .A(n27960), .B(n25491), .C(n25492), .D(n27962), .Y(n34132)
         );
  OAI22X1 U28610 ( .A(n27961), .B(n25320), .C(n32918), .D(n25322), .Y(n34131)
         );
  NOR2X1 U28611 ( .A(n34133), .B(n34134), .Y(n34123) );
  OAI22X1 U28612 ( .A(n25244), .B(n25316), .C(n25239), .D(n25318), .Y(n34134)
         );
  OAI22X1 U28613 ( .A(n27954), .B(n25498), .C(n29286), .D(n25499), .Y(n34133)
         );
  AOI22X1 U28614 ( .A(n25500), .B(reg_A[11]), .C(n25501), .D(reg_A[10]), .Y(
        n34104) );
  AOI22X1 U28615 ( .A(n25502), .B(reg_A[9]), .C(n25503), .D(reg_A[13]), .Y(
        n34103) );
  INVX1 U28616 ( .A(n34135), .Y(n32967) );
  OAI21X1 U28617 ( .A(n26742), .B(n31833), .C(n34136), .Y(n34135) );
  NAND3X1 U28618 ( .A(n32933), .B(n32934), .C(reg_A[2]), .Y(n34136) );
  NAND2X1 U28619 ( .A(n25110), .B(reg_B[30]), .Y(n31833) );
  NAND3X1 U28620 ( .A(n34137), .B(n34138), .C(n34139), .Y(n34094) );
  NOR2X1 U28621 ( .A(n34140), .B(n34141), .Y(n34139) );
  OAI22X1 U28622 ( .A(n34142), .B(n31782), .C(n29305), .D(n27944), .Y(n34141)
         );
  OAI22X1 U28623 ( .A(n34143), .B(n28033), .C(n25264), .D(n30620), .Y(n34140)
         );
  NAND2X1 U28624 ( .A(reg_A[5]), .B(n25110), .Y(n30620) );
  INVX1 U28625 ( .A(n29243), .Y(n34143) );
  NAND2X1 U28626 ( .A(n34144), .B(n34145), .Y(n29243) );
  AOI22X1 U28627 ( .A(n25156), .B(reg_A[6]), .C(n25142), .D(reg_A[7]), .Y(
        n34145) );
  AOI22X1 U28628 ( .A(n25258), .B(reg_A[8]), .C(reg_A[9]), .D(n26761), .Y(
        n34144) );
  AOI22X1 U28629 ( .A(n30644), .B(n34146), .C(n26772), .D(n34147), .Y(n34138)
         );
  AOI22X1 U28630 ( .A(reg_A[3]), .B(n32984), .C(n32985), .D(reg_A[2]), .Y(
        n34137) );
  NAND3X1 U28631 ( .A(n34148), .B(n34149), .C(n34150), .Y(result[29]) );
  NOR2X1 U28632 ( .A(n34151), .B(n34152), .Y(n34150) );
  OR2X1 U28633 ( .A(n34153), .B(n34154), .Y(n34152) );
  OAI22X1 U28634 ( .A(n29286), .B(n26136), .C(n27954), .D(n26812), .Y(n34154)
         );
  OAI21X1 U28635 ( .A(n26854), .B(n33928), .C(n34155), .Y(n34153) );
  AOI22X1 U28636 ( .A(n26269), .B(reg_A[25]), .C(reg_A[24]), .D(n34156), .Y(
        n34155) );
  NAND2X1 U28637 ( .A(n34157), .B(n34158), .Y(n33928) );
  AOI22X1 U28638 ( .A(n26313), .B(n25244), .C(n26314), .D(n25239), .Y(n34158)
         );
  AOI22X1 U28639 ( .A(reg_B[1]), .B(n34159), .C(reg_B[2]), .D(n34160), .Y(
        n34157) );
  INVX1 U28640 ( .A(n34161), .Y(n34159) );
  NAND3X1 U28641 ( .A(n34162), .B(n34163), .C(n34164), .Y(n34151) );
  AOI21X1 U28642 ( .A(n25170), .B(n34165), .C(n34166), .Y(n34164) );
  OAI21X1 U28643 ( .A(n34167), .B(n34168), .C(n34169), .Y(n34166) );
  NAND3X1 U28644 ( .A(n33998), .B(n33865), .C(n26186), .Y(n34169) );
  OAI21X1 U28645 ( .A(n34012), .B(n25239), .C(n34170), .Y(n33998) );
  AOI22X1 U28646 ( .A(n34000), .B(reg_A[27]), .C(n33809), .D(reg_A[25]), .Y(
        n34170) );
  NAND2X1 U28647 ( .A(n26504), .B(n33841), .Y(n34168) );
  MUX2X1 U28648 ( .B(n27961), .A(n32918), .S(n33865), .Y(n33841) );
  INVX1 U28649 ( .A(n34171), .Y(n34165) );
  AOI22X1 U28650 ( .A(n34172), .B(reg_B[31]), .C(n34021), .D(n34173), .Y(
        n34171) );
  NAND2X1 U28651 ( .A(n34174), .B(n34175), .Y(n34021) );
  AOI22X1 U28652 ( .A(n33921), .B(n34176), .C(n34000), .D(n33913), .Y(n34175)
         );
  NAND2X1 U28653 ( .A(n34177), .B(n34178), .Y(n33921) );
  AOI22X1 U28654 ( .A(n34179), .B(n34180), .C(n25103), .D(reg_A[13]), .Y(
        n34178) );
  NOR2X1 U28655 ( .A(n31782), .B(n29265), .Y(n34179) );
  AOI22X1 U28656 ( .A(reg_A[29]), .B(n25110), .C(n30644), .D(reg_A[21]), .Y(
        n34177) );
  AOI22X1 U28657 ( .A(n33809), .B(n33920), .C(n34015), .D(n34181), .Y(n34174)
         );
  OAI21X1 U28658 ( .A(n34182), .B(n34183), .C(n26267), .Y(n34163) );
  OAI22X1 U28659 ( .A(n34184), .B(n25264), .C(n33959), .D(n29305), .Y(n34183)
         );
  OAI22X1 U28660 ( .A(n34185), .B(n26758), .C(n33924), .D(n25262), .Y(n34182)
         );
  AND2X1 U28661 ( .A(n34186), .B(n34187), .Y(n33924) );
  AOI22X1 U28662 ( .A(n34188), .B(reg_A[17]), .C(n34180), .D(reg_A[21]), .Y(
        n34187) );
  AOI22X1 U28663 ( .A(n34189), .B(reg_A[29]), .C(n34190), .D(reg_A[25]), .Y(
        n34186) );
  AOI22X1 U28664 ( .A(n33930), .B(n32319), .C(n34191), .D(n34192), .Y(n34162)
         );
  AND2X1 U28665 ( .A(n34193), .B(n34194), .Y(n33930) );
  AOI22X1 U28666 ( .A(n26292), .B(n27960), .C(n26293), .D(n25239), .Y(n34194)
         );
  AOI22X1 U28667 ( .A(n26294), .B(n27962), .C(n26295), .D(n25244), .Y(n34193)
         );
  NOR2X1 U28668 ( .A(n34195), .B(n34196), .Y(n34149) );
  OAI21X1 U28669 ( .A(n25994), .B(n34197), .C(n34198), .Y(n34196) );
  INVX1 U28670 ( .A(n34199), .Y(n34198) );
  OAI22X1 U28671 ( .A(n33981), .B(n26525), .C(n34200), .D(n26012), .Y(n34199)
         );
  OAI21X1 U28672 ( .A(n34201), .B(n26208), .C(n34202), .Y(n33981) );
  AOI22X1 U28673 ( .A(n25026), .B(n33871), .C(n33803), .D(n26030), .Y(n34202)
         );
  INVX1 U28674 ( .A(n34203), .Y(n33803) );
  MUX2X1 U28675 ( .B(n34204), .A(n34205), .S(reg_B[2]), .Y(n34203) );
  OAI21X1 U28676 ( .A(reg_A[29]), .B(n25063), .C(n34206), .Y(n34204) );
  AOI22X1 U28677 ( .A(n26038), .B(n25232), .C(reg_B[0]), .D(n34207), .Y(n34206) );
  OAI21X1 U28678 ( .A(n26205), .B(n27961), .C(n34208), .Y(n34195) );
  AOI22X1 U28679 ( .A(n33999), .B(n30616), .C(reg_A[27]), .D(n33943), .Y(
        n34208) );
  INVX1 U28680 ( .A(n34209), .Y(n33999) );
  OAI21X1 U28681 ( .A(n34210), .B(n29255), .C(n34211), .Y(n34209) );
  AOI22X1 U28682 ( .A(n33893), .B(n34176), .C(n34000), .D(n34212), .Y(n34211)
         );
  NAND2X1 U28683 ( .A(n34213), .B(n34214), .Y(n33893) );
  MUX2X1 U28684 ( .B(n34215), .A(n34216), .S(reg_B[29]), .Y(n34214) );
  NOR2X1 U28685 ( .A(n34217), .B(n31782), .Y(n34215) );
  AOI22X1 U28686 ( .A(n25110), .B(n25239), .C(n30644), .D(n25232), .Y(n34213)
         );
  INVX1 U28687 ( .A(n30287), .Y(n26205) );
  NOR2X1 U28688 ( .A(n34218), .B(n34219), .Y(n34148) );
  OAI21X1 U28689 ( .A(n25239), .B(n30282), .C(n34220), .Y(n34219) );
  MUX2X1 U28690 ( .B(n33878), .A(n34221), .S(reg_B[30]), .Y(n34220) );
  NOR2X1 U28691 ( .A(n25032), .B(n34222), .Y(n34221) );
  OAI22X1 U28692 ( .A(n34223), .B(n34224), .C(n25342), .D(n34225), .Y(n33878)
         );
  MUX2X1 U28693 ( .B(n34226), .A(n34227), .S(reg_B[29]), .Y(n34225) );
  MUX2X1 U28694 ( .B(n27960), .A(n27962), .S(reg_B[31]), .Y(n34227) );
  OAI21X1 U28695 ( .A(n34228), .B(n33955), .C(n25188), .Y(n34224) );
  OAI22X1 U28696 ( .A(n34229), .B(n33957), .C(n34226), .D(n34230), .Y(n34223)
         );
  MUX2X1 U28697 ( .B(n25239), .A(n25244), .S(reg_B[31]), .Y(n34226) );
  OAI21X1 U28698 ( .A(n29255), .B(n33991), .C(n34231), .Y(n34218) );
  AOI22X1 U28699 ( .A(n26045), .B(n34232), .C(n25109), .D(n34233), .Y(n34231)
         );
  NAND3X1 U28700 ( .A(n34234), .B(n34235), .C(n34236), .Y(n34232) );
  NOR2X1 U28701 ( .A(n34237), .B(n34238), .Y(n34236) );
  OAI21X1 U28702 ( .A(n25204), .B(n25239), .C(n34239), .Y(n34238) );
  AOI22X1 U28703 ( .A(n27387), .B(reg_A[25]), .C(n28312), .D(reg_A[27]), .Y(
        n34239) );
  NAND2X1 U28704 ( .A(n34240), .B(n34241), .Y(n34237) );
  AOI22X1 U28705 ( .A(n25440), .B(reg_A[23]), .C(n34242), .D(n25610), .Y(
        n34241) );
  AOI22X1 U28706 ( .A(reg_A[28]), .B(n25441), .C(n25442), .D(reg_A[26]), .Y(
        n34240) );
  NOR2X1 U28707 ( .A(n34243), .B(n34244), .Y(n34235) );
  OAI22X1 U28708 ( .A(n30587), .B(n26229), .C(n27962), .D(n25449), .Y(n34244)
         );
  OAI21X1 U28709 ( .A(n27953), .B(n25451), .C(n34245), .Y(n34243) );
  OAI21X1 U28710 ( .A(n34246), .B(n34247), .C(n25044), .Y(n34245) );
  NAND3X1 U28711 ( .A(n34248), .B(n34249), .C(n34250), .Y(n34247) );
  NOR2X1 U28712 ( .A(n34251), .B(n34252), .Y(n34250) );
  OAI21X1 U28713 ( .A(n25239), .B(n25043), .C(n34253), .Y(n34252) );
  AOI22X1 U28714 ( .A(n25135), .B(reg_A[28]), .C(n25252), .D(reg_A[27]), .Y(
        n34253) );
  NAND2X1 U28715 ( .A(n34254), .B(n34255), .Y(n34251) );
  AOI22X1 U28716 ( .A(n25136), .B(reg_A[26]), .C(reg_A[23]), .D(n25253), .Y(
        n34255) );
  AOI22X1 U28717 ( .A(n25075), .B(reg_A[25]), .C(reg_A[24]), .D(n25123), .Y(
        n34254) );
  NOR2X1 U28718 ( .A(n34256), .B(n34257), .Y(n34249) );
  OAI22X1 U28719 ( .A(n25034), .B(n25232), .C(n25030), .D(n25230), .Y(n34257)
         );
  OAI22X1 U28720 ( .A(n25036), .B(n25220), .C(n25037), .D(n30587), .Y(n34256)
         );
  NOR2X1 U28721 ( .A(n34258), .B(n34259), .Y(n34248) );
  OAI22X1 U28722 ( .A(n27953), .B(n25231), .C(n25224), .D(n25473), .Y(n34259)
         );
  OAI22X1 U28723 ( .A(n25250), .B(n25229), .C(n29279), .D(n25475), .Y(n34258)
         );
  NAND3X1 U28724 ( .A(n34260), .B(n34261), .C(n34262), .Y(n34246) );
  NOR2X1 U28725 ( .A(n34263), .B(n34264), .Y(n34262) );
  OAI21X1 U28726 ( .A(n25208), .B(n25482), .C(n34265), .Y(n34264) );
  AOI22X1 U28727 ( .A(reg_A[12]), .B(n25246), .C(reg_A[13]), .D(n25247), .Y(
        n34265) );
  NAND2X1 U28728 ( .A(n34266), .B(n34267), .Y(n34263) );
  AOI22X1 U28729 ( .A(reg_A[10]), .B(n25487), .C(reg_A[11]), .D(n25241), .Y(
        n34267) );
  AOI22X1 U28730 ( .A(n25339), .B(reg_A[9]), .C(n25257), .D(reg_A[8]), .Y(
        n34266) );
  NOR2X1 U28731 ( .A(n34268), .B(n34269), .Y(n34261) );
  OAI22X1 U28732 ( .A(n26677), .B(n25491), .C(n25132), .D(n25492), .Y(n34269)
         );
  OAI22X1 U28733 ( .A(n29265), .B(n25320), .C(n30569), .D(n25322), .Y(n34268)
         );
  NOR2X1 U28734 ( .A(n34270), .B(n34271), .Y(n34260) );
  OAI22X1 U28735 ( .A(n25130), .B(n25316), .C(n25128), .D(n25318), .Y(n34271)
         );
  OAI22X1 U28736 ( .A(n26742), .B(n25498), .C(n25177), .D(n25499), .Y(n34270)
         );
  NOR2X1 U28737 ( .A(n34272), .B(n34273), .Y(n34234) );
  OAI22X1 U28738 ( .A(n25220), .B(n28362), .C(n25224), .D(n28363), .Y(n34273)
         );
  OAI22X1 U28739 ( .A(n25230), .B(n30443), .C(n25232), .D(n30444), .Y(n34272)
         );
  NAND3X1 U28740 ( .A(n34274), .B(n34275), .C(n34276), .Y(result[28]) );
  NOR2X1 U28741 ( .A(n34277), .B(n34278), .Y(n34276) );
  NAND3X1 U28742 ( .A(n34279), .B(n34280), .C(n34281), .Y(n34278) );
  AOI21X1 U28743 ( .A(reg_A[21]), .B(n34282), .C(n34283), .Y(n34281) );
  OAI22X1 U28744 ( .A(n34017), .B(n34284), .C(n25206), .D(n26625), .Y(n34283)
         );
  INVX1 U28745 ( .A(n34233), .Y(n34017) );
  NAND2X1 U28746 ( .A(n34285), .B(n30559), .Y(n34233) );
  AOI22X1 U28747 ( .A(reg_A[23]), .B(n26353), .C(reg_A[19]), .D(n26346), .Y(
        n34280) );
  AOI22X1 U28748 ( .A(reg_A[22]), .B(n26347), .C(reg_A[24]), .D(n26348), .Y(
        n34279) );
  NAND3X1 U28749 ( .A(n34286), .B(n34287), .C(n34288), .Y(n34277) );
  NOR2X1 U28750 ( .A(n34289), .B(n34290), .Y(n34288) );
  OAI22X1 U28751 ( .A(n26355), .B(n30587), .C(n26012), .D(n34291), .Y(n34290)
         );
  INVX1 U28752 ( .A(n26551), .Y(n26355) );
  OAI22X1 U28753 ( .A(n26525), .B(n34200), .C(n26526), .D(n25224), .Y(n34289)
         );
  OAI21X1 U28754 ( .A(n34292), .B(n26208), .C(n34293), .Y(n34200) );
  AOI22X1 U28755 ( .A(n25026), .B(n33985), .C(n34294), .D(n26030), .Y(n34293)
         );
  INVX1 U28756 ( .A(n33982), .Y(n34294) );
  MUX2X1 U28757 ( .B(n34295), .A(n34296), .S(reg_B[2]), .Y(n33982) );
  OAI21X1 U28758 ( .A(reg_A[28]), .B(n25063), .C(n34297), .Y(n34295) );
  AOI22X1 U28759 ( .A(n26038), .B(n30587), .C(reg_B[0]), .D(n34298), .Y(n34297) );
  AOI22X1 U28760 ( .A(n34192), .B(n30616), .C(reg_A[17]), .D(n26357), .Y(
        n34287) );
  INVX1 U28761 ( .A(n34299), .Y(n34192) );
  OAI21X1 U28762 ( .A(n34300), .B(n29255), .C(n34301), .Y(n34299) );
  AOI22X1 U28763 ( .A(n33969), .B(n34176), .C(n34000), .D(n33972), .Y(n34301)
         );
  NAND2X1 U28764 ( .A(n34302), .B(n34303), .Y(n33969) );
  MUX2X1 U28765 ( .B(n34304), .A(n34305), .S(reg_B[29]), .Y(n34303) );
  NOR2X1 U28766 ( .A(n34306), .B(n31782), .Y(n34304) );
  AOI22X1 U28767 ( .A(n25110), .B(n25244), .C(n30644), .D(n30587), .Y(n34302)
         );
  AOI22X1 U28768 ( .A(reg_A[28]), .B(n26398), .C(reg_A[27]), .D(n26358), .Y(
        n34286) );
  NOR2X1 U28769 ( .A(n34307), .B(n34308), .Y(n34275) );
  OR2X1 U28770 ( .A(n34309), .B(n34310), .Y(n34308) );
  OAI21X1 U28771 ( .A(n26370), .B(n25250), .C(n34311), .Y(n34310) );
  OAI21X1 U28772 ( .A(n34312), .B(n34313), .C(n25188), .Y(n34311) );
  OAI22X1 U28773 ( .A(n34009), .B(n34314), .C(n33957), .D(n34315), .Y(n34313)
         );
  OAI21X1 U28774 ( .A(n25262), .B(n34316), .C(n34317), .Y(n34312) );
  AOI21X1 U28775 ( .A(n34189), .B(n34318), .C(n34319), .Y(n34317) );
  OAI21X1 U28776 ( .A(n26373), .B(n27960), .C(n34320), .Y(n34309) );
  OAI21X1 U28777 ( .A(n34321), .B(n34322), .C(n26267), .Y(n34320) );
  OAI22X1 U28778 ( .A(n34323), .B(n25264), .C(n34184), .D(n29305), .Y(n34322)
         );
  OAI22X1 U28779 ( .A(n33959), .B(n26758), .C(n34185), .D(n25262), .Y(n34321)
         );
  INVX1 U28780 ( .A(n34008), .Y(n34185) );
  NAND3X1 U28781 ( .A(n34316), .B(n34324), .C(n34325), .Y(n34008) );
  AOI22X1 U28782 ( .A(n34190), .B(reg_A[24]), .C(n34180), .D(reg_A[20]), .Y(
        n34325) );
  NAND2X1 U28783 ( .A(n34189), .B(reg_A[28]), .Y(n34316) );
  NOR2X1 U28784 ( .A(n26472), .B(n28206), .Y(n26373) );
  NAND3X1 U28785 ( .A(n34326), .B(n34327), .C(n34328), .Y(n34307) );
  AOI22X1 U28786 ( .A(n34329), .B(n34172), .C(reg_B[31]), .D(n34330), .Y(
        n34328) );
  OAI21X1 U28787 ( .A(n34331), .B(n26151), .C(n34332), .Y(n34330) );
  AOI22X1 U28788 ( .A(n34333), .B(n25170), .C(n34334), .D(n25932), .Y(n34332)
         );
  INVX1 U28789 ( .A(n34335), .Y(n34334) );
  OAI21X1 U28790 ( .A(n34336), .B(n34167), .C(n34337), .Y(n34172) );
  AOI22X1 U28791 ( .A(n25097), .B(n34338), .C(n25589), .D(n34339), .Y(n34337)
         );
  OAI22X1 U28792 ( .A(n34012), .B(n25244), .C(n27962), .D(n33966), .Y(n34339)
         );
  INVX1 U28793 ( .A(n34340), .Y(n34338) );
  AOI22X1 U28794 ( .A(n34341), .B(n34015), .C(n34176), .D(n33948), .Y(n34340)
         );
  NAND2X1 U28795 ( .A(n34342), .B(n34343), .Y(n33948) );
  AOI21X1 U28796 ( .A(n25103), .B(reg_A[12]), .C(n34344), .Y(n34343) );
  OAI21X1 U28797 ( .A(n34345), .B(n33955), .C(n34346), .Y(n34344) );
  NAND3X1 U28798 ( .A(reg_A[4]), .B(reg_B[27]), .C(n34180), .Y(n34346) );
  INVX1 U28799 ( .A(n34347), .Y(n34345) );
  AOI22X1 U28800 ( .A(reg_A[28]), .B(n25110), .C(n30644), .D(reg_A[20]), .Y(
        n34342) );
  NAND3X1 U28801 ( .A(n34348), .B(n33955), .C(n26504), .Y(n34326) );
  OAI21X1 U28802 ( .A(n25262), .B(n25244), .C(n34349), .Y(n34348) );
  INVX1 U28803 ( .A(n34318), .Y(n34349) );
  OAI21X1 U28804 ( .A(n25264), .B(n27960), .C(n34350), .Y(n34318) );
  AOI22X1 U28805 ( .A(n25142), .B(reg_A[27]), .C(reg_A[26]), .D(n25258), .Y(
        n34350) );
  NOR2X1 U28806 ( .A(n34351), .B(n34352), .Y(n34274) );
  OAI21X1 U28807 ( .A(n25239), .B(n26136), .C(n34353), .Y(n34352) );
  AOI22X1 U28808 ( .A(n26451), .B(reg_A[31]), .C(n26310), .D(reg_A[30]), .Y(
        n34353) );
  OR2X1 U28809 ( .A(n34354), .B(n34355), .Y(n34351) );
  OAI22X1 U28810 ( .A(n26420), .B(n34356), .C(n26421), .D(n34357), .Y(n34355)
         );
  OAI21X1 U28811 ( .A(n26393), .B(n27961), .C(n34358), .Y(n34354) );
  OAI21X1 U28812 ( .A(n34359), .B(n34360), .C(n25840), .Y(n34358) );
  NAND3X1 U28813 ( .A(n34361), .B(n34362), .C(n34363), .Y(n34360) );
  NOR2X1 U28814 ( .A(n34364), .B(n34365), .Y(n34363) );
  OAI22X1 U28815 ( .A(n29279), .B(n25229), .C(n25208), .D(n25475), .Y(n34365)
         );
  OAI22X1 U28816 ( .A(n26431), .B(n27962), .C(n32918), .D(n25784), .Y(n34364)
         );
  AOI22X1 U28817 ( .A(n25647), .B(reg_A[4]), .C(n25648), .D(reg_A[1]), .Y(
        n34362) );
  AOI22X1 U28818 ( .A(n26432), .B(reg_A[2]), .C(n25324), .D(reg_A[0]), .Y(
        n34361) );
  NAND3X1 U28819 ( .A(n34366), .B(n34367), .C(n34368), .Y(n34359) );
  NOR2X1 U28820 ( .A(n34369), .B(n34370), .Y(n34368) );
  OAI22X1 U28821 ( .A(n26677), .B(n25492), .C(n25331), .D(n25147), .Y(n34370)
         );
  OAI21X1 U28822 ( .A(n25146), .B(n25243), .C(n34371), .Y(n34369) );
  AOI22X1 U28823 ( .A(reg_A[11]), .B(n25246), .C(reg_A[12]), .D(n25247), .Y(
        n34371) );
  AOI22X1 U28824 ( .A(n25338), .B(reg_A[5]), .C(n25339), .D(reg_A[8]), .Y(
        n34367) );
  AOI22X1 U28825 ( .A(n25257), .B(reg_A[7]), .C(n25857), .D(reg_A[3]), .Y(
        n34366) );
  NAND2X1 U28826 ( .A(n34372), .B(n34373), .Y(result[27]) );
  NOR2X1 U28827 ( .A(n34374), .B(n34375), .Y(n34373) );
  NAND3X1 U28828 ( .A(n34376), .B(n34377), .C(n34378), .Y(n34375) );
  NOR2X1 U28829 ( .A(n34379), .B(n34380), .Y(n34378) );
  OAI21X1 U28830 ( .A(n28586), .B(n27960), .C(n34381), .Y(n34380) );
  OAI21X1 U28831 ( .A(n34382), .B(n34383), .C(n26267), .Y(n34381) );
  OAI22X1 U28832 ( .A(n34384), .B(n25264), .C(n34323), .D(n29305), .Y(n34383)
         );
  OAI22X1 U28833 ( .A(n34184), .B(n26758), .C(n33959), .D(n25262), .Y(n34382)
         );
  INVX1 U28834 ( .A(n34385), .Y(n33959) );
  OAI21X1 U28835 ( .A(n26714), .B(n34009), .C(n34386), .Y(n34385) );
  AOI22X1 U28836 ( .A(n34180), .B(reg_A[19]), .C(n34189), .D(reg_A[27]), .Y(
        n34386) );
  OAI22X1 U28837 ( .A(n34387), .B(n34388), .C(n27954), .D(n30924), .Y(n34379)
         );
  INVX1 U28838 ( .A(n26482), .Y(n30924) );
  AOI22X1 U28839 ( .A(n28572), .B(reg_A[18]), .C(n28576), .D(reg_A[21]), .Y(
        n34377) );
  AOI22X1 U28840 ( .A(n25181), .B(reg_A[23]), .C(n28717), .D(reg_A[19]), .Y(
        n34376) );
  NAND3X1 U28841 ( .A(n34389), .B(n34390), .C(n34391), .Y(n34374) );
  NOR2X1 U28842 ( .A(n34392), .B(n34393), .Y(n34391) );
  OAI21X1 U28843 ( .A(n25032), .B(n34394), .C(n34395), .Y(n34393) );
  OAI21X1 U28844 ( .A(n26179), .B(n28835), .C(reg_A[27]), .Y(n34395) );
  INVX1 U28845 ( .A(n34396), .Y(n34394) );
  MUX2X1 U28846 ( .B(n34222), .A(n34397), .S(reg_B[30]), .Y(n34396) );
  OAI21X1 U28847 ( .A(n33863), .B(n34009), .C(n34398), .Y(n34222) );
  AOI21X1 U28848 ( .A(n33839), .B(n33955), .C(n34399), .Y(n34398) );
  INVX1 U28849 ( .A(n34400), .Y(n33839) );
  MUX2X1 U28850 ( .B(n34401), .A(n34402), .S(reg_B[31]), .Y(n34400) );
  MUX2X1 U28851 ( .B(reg_A[27]), .A(reg_A[19]), .S(reg_B[28]), .Y(n34401) );
  OAI21X1 U28852 ( .A(n34403), .B(n34404), .C(n34327), .Y(n34392) );
  AOI22X1 U28853 ( .A(n25382), .B(n33874), .C(n26480), .D(n32933), .Y(n34404)
         );
  AOI22X1 U28854 ( .A(n34333), .B(n34329), .C(n34004), .D(n34405), .Y(n34390)
         );
  INVX1 U28855 ( .A(n34406), .Y(n34329) );
  AOI21X1 U28856 ( .A(n34407), .B(n34408), .C(n25403), .Y(n34333) );
  AOI22X1 U28857 ( .A(n34409), .B(n34015), .C(n34181), .D(n33809), .Y(n34408)
         );
  AOI22X1 U28858 ( .A(n33920), .B(n34000), .C(n33913), .D(n32934), .Y(n34407)
         );
  NAND2X1 U28859 ( .A(n34410), .B(n34411), .Y(n33913) );
  AOI22X1 U28860 ( .A(n33922), .B(reg_A[3]), .C(n33923), .D(reg_A[11]), .Y(
        n34411) );
  AOI22X1 U28861 ( .A(reg_A[19]), .B(n33919), .C(reg_A[27]), .D(n32933), .Y(
        n34410) );
  AOI22X1 U28862 ( .A(n28549), .B(reg_A[16]), .C(n28649), .D(reg_A[17]), .Y(
        n34389) );
  NOR2X1 U28863 ( .A(n34412), .B(n34413), .Y(n34372) );
  NAND3X1 U28864 ( .A(n34414), .B(n34415), .C(n34416), .Y(n34413) );
  NOR2X1 U28865 ( .A(n34417), .B(n34418), .Y(n34416) );
  OAI21X1 U28866 ( .A(n25264), .B(n33991), .C(n34419), .Y(n34418) );
  MUX2X1 U28867 ( .B(n34420), .A(n34421), .S(reg_B[31]), .Y(n34419) );
  NOR2X1 U28868 ( .A(n34422), .B(n25697), .Y(n34421) );
  NOR2X1 U28869 ( .A(n28213), .B(n34331), .Y(n34420) );
  AOI22X1 U28870 ( .A(n32934), .B(reg_A[27]), .C(reg_A[25]), .D(n34000), .Y(
        n34331) );
  OAI22X1 U28871 ( .A(n30587), .B(n28562), .C(n25255), .D(n26625), .Y(n34417)
         );
  AOI22X1 U28872 ( .A(n34423), .B(n26028), .C(n34424), .D(n26260), .Y(n34415)
         );
  INVX1 U28873 ( .A(n34291), .Y(n34423) );
  NAND2X1 U28874 ( .A(n34425), .B(n34426), .Y(n34291) );
  AOI22X1 U28875 ( .A(n25025), .B(n34427), .C(n25026), .D(n34205), .Y(n34426)
         );
  AOI22X1 U28876 ( .A(n26032), .B(n33871), .C(n26530), .D(n34428), .Y(n34425)
         );
  OAI21X1 U28877 ( .A(reg_A[27]), .B(n25063), .C(n34429), .Y(n33871) );
  AOI22X1 U28878 ( .A(n26038), .B(n25220), .C(reg_B[0]), .D(n34430), .Y(n34429) );
  AOI22X1 U28879 ( .A(n34431), .B(n26262), .C(reg_A[26]), .D(n26626), .Y(
        n34414) );
  NAND3X1 U28880 ( .A(n34432), .B(n34433), .C(n34434), .Y(n34412) );
  NOR2X1 U28881 ( .A(n34435), .B(n34436), .Y(n34434) );
  OAI21X1 U28882 ( .A(n28664), .B(n27962), .C(n34437), .Y(n34436) );
  OAI21X1 U28883 ( .A(n34438), .B(n34439), .C(n25840), .Y(n34437) );
  NAND3X1 U28884 ( .A(n34440), .B(n34441), .C(n34442), .Y(n34439) );
  NOR2X1 U28885 ( .A(n34443), .B(n34444), .Y(n34442) );
  OAI21X1 U28886 ( .A(n32918), .B(n25228), .C(n34445), .Y(n34444) );
  AOI22X1 U28887 ( .A(n25635), .B(reg_A[15]), .C(n25325), .D(reg_A[14]), .Y(
        n34445) );
  OAI21X1 U28888 ( .A(n25206), .B(n25475), .C(n34446), .Y(n34443) );
  AOI22X1 U28889 ( .A(n25222), .B(reg_A[16]), .C(n25637), .D(reg_A[17]), .Y(
        n34446) );
  NOR2X1 U28890 ( .A(n34447), .B(n34448), .Y(n34441) );
  OAI22X1 U28891 ( .A(n26431), .B(n26714), .C(n25030), .D(n30587), .Y(n34448)
         );
  OAI22X1 U28892 ( .A(n25033), .B(n25232), .C(n27960), .D(n25133), .Y(n34447)
         );
  AOI21X1 U28893 ( .A(reg_A[19]), .B(n25124), .C(n34449), .Y(n34440) );
  OAI22X1 U28894 ( .A(n25037), .B(n25224), .C(n26703), .D(n25230), .Y(n34449)
         );
  NAND3X1 U28895 ( .A(n34450), .B(n34451), .C(n34452), .Y(n34438) );
  NOR2X1 U28896 ( .A(n34453), .B(n34454), .Y(n34452) );
  OAI21X1 U28897 ( .A(n25132), .B(n25238), .C(n34455), .Y(n34454) );
  AOI22X1 U28898 ( .A(n25242), .B(reg_A[5]), .C(n25338), .D(reg_A[4]), .Y(
        n34455) );
  NAND2X1 U28899 ( .A(n34456), .B(n34457), .Y(n34453) );
  AOI22X1 U28900 ( .A(reg_A[10]), .B(n25246), .C(reg_A[11]), .D(n25247), .Y(
        n34457) );
  AOI22X1 U28901 ( .A(n25487), .B(reg_A[8]), .C(n25241), .D(reg_A[9]), .Y(
        n34456) );
  NOR2X1 U28902 ( .A(n34458), .B(n34459), .Y(n34451) );
  OAI22X1 U28903 ( .A(n26742), .B(n25318), .C(n25130), .D(n25320), .Y(n34459)
         );
  OAI22X1 U28904 ( .A(n25128), .B(n25322), .C(n26677), .D(n26719), .Y(n34458)
         );
  AOI21X1 U28905 ( .A(reg_A[24]), .B(n25136), .C(n34460), .Y(n34450) );
  OAI22X1 U28906 ( .A(n27961), .B(n25784), .C(n25177), .D(n25316), .Y(n34460)
         );
  OAI22X1 U28907 ( .A(n33964), .B(n34335), .C(n25244), .D(n26136), .Y(n34435)
         );
  NAND2X1 U28908 ( .A(n34461), .B(n34462), .Y(n34335) );
  AOI22X1 U28909 ( .A(n32934), .B(n34212), .C(n34000), .D(n34216), .Y(n34462)
         );
  INVX1 U28910 ( .A(n33842), .Y(n34212) );
  AOI21X1 U28911 ( .A(n32918), .B(n32933), .C(n34463), .Y(n33842) );
  OAI22X1 U28912 ( .A(n31782), .B(n34464), .C(n34465), .D(reg_A[19]), .Y(
        n34463) );
  AOI22X1 U28913 ( .A(n33809), .B(n34466), .C(n34015), .D(n34467), .Y(n34461)
         );
  AOI22X1 U28914 ( .A(n25149), .B(reg_A[22]), .C(n26451), .D(reg_A[30]), .Y(
        n34433) );
  AOI22X1 U28915 ( .A(n34468), .B(n25150), .C(n26310), .D(reg_A[29]), .Y(
        n34432) );
  INVX1 U28916 ( .A(n34197), .Y(n34468) );
  OAI21X1 U28917 ( .A(reg_B[2]), .B(n33868), .C(n34469), .Y(n34197) );
  AOI22X1 U28918 ( .A(n26455), .B(n25250), .C(n26456), .D(n33802), .Y(n34469)
         );
  INVX1 U28919 ( .A(n34470), .Y(n33802) );
  AND2X1 U28920 ( .A(n34471), .B(n34472), .Y(n33868) );
  AOI22X1 U28921 ( .A(n26460), .B(n25220), .C(n26461), .D(n32918), .Y(n34472)
         );
  AOI22X1 U28922 ( .A(n26462), .B(n27961), .C(n26463), .D(n25224), .Y(n34471)
         );
  NAND2X1 U28923 ( .A(n34473), .B(n34474), .Y(result[26]) );
  NOR2X1 U28924 ( .A(n34475), .B(n34476), .Y(n34474) );
  NAND3X1 U28925 ( .A(n34477), .B(n34478), .C(n34479), .Y(n34476) );
  NOR2X1 U28926 ( .A(n34480), .B(n34481), .Y(n34479) );
  OAI21X1 U28927 ( .A(n26573), .B(n27962), .C(n34482), .Y(n34481) );
  OAI21X1 U28928 ( .A(n34483), .B(n34484), .C(n25188), .Y(n34482) );
  OAI21X1 U28929 ( .A(n34009), .B(n33958), .C(n34324), .Y(n34484) );
  INVX1 U28930 ( .A(n34319), .Y(n34324) );
  NOR2X1 U28931 ( .A(n34485), .B(n33955), .Y(n34319) );
  NAND2X1 U28932 ( .A(n34486), .B(n34487), .Y(n33958) );
  AOI22X1 U28933 ( .A(n25156), .B(n25230), .C(n25142), .D(n25232), .Y(n34487)
         );
  AOI22X1 U28934 ( .A(n25258), .B(n30587), .C(n26761), .D(n25220), .Y(n34486)
         );
  NOR2X1 U28935 ( .A(reg_B[29]), .B(n33956), .Y(n34483) );
  NAND2X1 U28936 ( .A(n34488), .B(n34489), .Y(n33956) );
  MUX2X1 U28937 ( .B(n34490), .A(n34491), .S(reg_B[28]), .Y(n34489) );
  NOR2X1 U28938 ( .A(reg_A[16]), .B(n34176), .Y(n34491) );
  OAI22X1 U28939 ( .A(reg_A[23]), .B(n25264), .C(reg_A[24]), .D(n29305), .Y(
        n34490) );
  AOI22X1 U28940 ( .A(n25156), .B(n34402), .C(n25142), .D(n34492), .Y(n34488)
         );
  MUX2X1 U28941 ( .B(reg_A[18]), .A(reg_A[26]), .S(n34493), .Y(n34402) );
  OAI21X1 U28942 ( .A(n34494), .B(n34495), .C(n34496), .Y(n34480) );
  OAI21X1 U28943 ( .A(n34497), .B(n34498), .C(n26267), .Y(n34496) );
  OAI22X1 U28944 ( .A(n34499), .B(n25264), .C(n34384), .D(n29305), .Y(n34498)
         );
  INVX1 U28945 ( .A(n34500), .Y(n34384) );
  INVX1 U28946 ( .A(n34501), .Y(n34499) );
  OAI22X1 U28947 ( .A(n34323), .B(n26758), .C(n34184), .D(n25262), .Y(n34497)
         );
  INVX1 U28948 ( .A(n34502), .Y(n34184) );
  OAI21X1 U28949 ( .A(n25230), .B(n34009), .C(n34503), .Y(n34502) );
  AOI22X1 U28950 ( .A(n34180), .B(reg_A[18]), .C(n34189), .D(reg_A[26]), .Y(
        n34503) );
  INVX1 U28951 ( .A(n34504), .Y(n34323) );
  AOI22X1 U28952 ( .A(reg_A[16]), .B(n26572), .C(reg_A[26]), .D(n26450), .Y(
        n34478) );
  AOI22X1 U28953 ( .A(n34505), .B(n28575), .C(n26451), .D(reg_A[29]), .Y(
        n34477) );
  INVX1 U28954 ( .A(n33973), .Y(n34505) );
  NAND3X1 U28955 ( .A(n34506), .B(n34507), .C(n34508), .Y(n34475) );
  NOR2X1 U28956 ( .A(n34509), .B(n34510), .Y(n34508) );
  OAI22X1 U28957 ( .A(n34016), .B(n34511), .C(n26584), .D(n33942), .Y(n34510)
         );
  NAND2X1 U28958 ( .A(n34512), .B(n34513), .Y(n33942) );
  AOI22X1 U28959 ( .A(n26593), .B(n25224), .C(n26594), .D(n25250), .Y(n34513)
         );
  AOI22X1 U28960 ( .A(n34514), .B(n26596), .C(n26597), .D(n34515), .Y(n34512)
         );
  OAI21X1 U28961 ( .A(reg_A[26]), .B(n26599), .C(n34516), .Y(n34514) );
  AOI22X1 U28962 ( .A(n26601), .B(n27962), .C(n26602), .D(n26714), .Y(n34516)
         );
  OAI21X1 U28963 ( .A(n34422), .B(n34406), .C(n34517), .Y(n34509) );
  AOI22X1 U28964 ( .A(n34518), .B(n34519), .C(reg_A[25]), .D(n34520), .Y(
        n34517) );
  OAI21X1 U28965 ( .A(n28213), .B(n33977), .C(n26483), .Y(n34520) );
  NOR2X1 U28966 ( .A(n34521), .B(n25697), .Y(n34518) );
  NAND2X1 U28967 ( .A(n25170), .B(n33865), .Y(n34406) );
  INVX1 U28968 ( .A(n34522), .Y(n34422) );
  OAI21X1 U28969 ( .A(n34336), .B(n34012), .C(n34523), .Y(n34522) );
  AOI22X1 U28970 ( .A(n34524), .B(n34000), .C(n25097), .D(n34525), .Y(n34523)
         );
  OAI21X1 U28971 ( .A(n34526), .B(n29255), .C(n34527), .Y(n34525) );
  AOI22X1 U28972 ( .A(n34000), .B(n34347), .C(n33809), .D(n34341), .Y(n34527)
         );
  INVX1 U28973 ( .A(n34528), .Y(n34526) );
  NOR2X1 U28974 ( .A(n26999), .B(n27962), .Y(n34524) );
  AOI22X1 U28975 ( .A(n25589), .B(reg_A[26]), .C(n33944), .D(n25097), .Y(
        n34336) );
  NAND2X1 U28976 ( .A(n34529), .B(n34530), .Y(n33944) );
  AOI22X1 U28977 ( .A(n33923), .B(reg_A[10]), .C(reg_A[26]), .D(n32933), .Y(
        n34530) );
  AOI22X1 U28978 ( .A(reg_A[18]), .B(n33919), .C(n33922), .D(reg_A[2]), .Y(
        n34529) );
  AOI22X1 U28979 ( .A(n34004), .B(n33890), .C(n30865), .D(reg_A[31]), .Y(
        n34507) );
  NOR2X1 U28980 ( .A(n27961), .B(n25031), .Y(n34004) );
  AOI22X1 U28981 ( .A(n26482), .B(reg_A[30]), .C(n34531), .D(n34191), .Y(
        n34506) );
  INVX1 U28982 ( .A(n34532), .Y(n34531) );
  NOR2X1 U28983 ( .A(n34533), .B(n34534), .Y(n34473) );
  NAND3X1 U28984 ( .A(n34535), .B(n34536), .C(n34537), .Y(n34534) );
  NOR2X1 U28985 ( .A(n34538), .B(n34539), .Y(n34537) );
  OAI22X1 U28986 ( .A(n26328), .B(n25220), .C(n32934), .D(n33991), .Y(n34539)
         );
  OAI22X1 U28987 ( .A(n27967), .B(n26625), .C(n25208), .D(n26917), .Y(n34538)
         );
  AOI22X1 U28988 ( .A(reg_A[23]), .B(n26472), .C(reg_A[17]), .D(n26346), .Y(
        n34536) );
  AOI22X1 U28989 ( .A(reg_A[20]), .B(n26347), .C(n26627), .D(reg_A[15]), .Y(
        n34535) );
  NAND3X1 U28990 ( .A(n34540), .B(n34541), .C(n34542), .Y(n34533) );
  NOR2X1 U28991 ( .A(n34543), .B(n34544), .Y(n34542) );
  OAI21X1 U28992 ( .A(n26534), .B(n25230), .C(n34545), .Y(n34544) );
  OAI21X1 U28993 ( .A(n34546), .B(n34547), .C(n25840), .Y(n34545) );
  NAND3X1 U28994 ( .A(n34548), .B(n34549), .C(n34550), .Y(n34547) );
  AOI21X1 U28995 ( .A(n25325), .B(reg_A[13]), .C(n34551), .Y(n34550) );
  OAI22X1 U28996 ( .A(n25255), .B(n25475), .C(n27960), .D(n25784), .Y(n34551)
         );
  AOI22X1 U28997 ( .A(n25257), .B(reg_A[5]), .C(n25857), .D(reg_A[1]), .Y(
        n34549) );
  AOI22X1 U28998 ( .A(n25647), .B(reg_A[2]), .C(n26432), .D(reg_A[0]), .Y(
        n34548) );
  NAND3X1 U28999 ( .A(n34552), .B(n34553), .C(n34554), .Y(n34546) );
  AOI21X1 U29000 ( .A(n25339), .B(reg_A[6]), .C(n34555), .Y(n34554) );
  OAI22X1 U29001 ( .A(n25130), .B(n25491), .C(n30569), .D(n25492), .Y(n34555)
         );
  AOI22X1 U29002 ( .A(n25246), .B(reg_A[9]), .C(reg_A[10]), .D(n25247), .Y(
        n34553) );
  AOI22X1 U29003 ( .A(n25487), .B(reg_A[7]), .C(n25241), .D(reg_A[8]), .Y(
        n34552) );
  OAI21X1 U29004 ( .A(n33964), .B(n34388), .C(n34556), .Y(n34543) );
  AOI22X1 U29005 ( .A(n26310), .B(reg_A[28]), .C(n26408), .D(reg_A[27]), .Y(
        n34556) );
  NAND2X1 U29006 ( .A(n34557), .B(n34558), .Y(n34388) );
  AOI22X1 U29007 ( .A(n32934), .B(n33972), .C(n34000), .D(n34305), .Y(n34558)
         );
  NAND2X1 U29008 ( .A(n34559), .B(n34560), .Y(n33972) );
  AOI22X1 U29009 ( .A(n33922), .B(n25128), .C(n33923), .D(n25147), .Y(n34560)
         );
  AOI22X1 U29010 ( .A(n33919), .B(n25224), .C(n32933), .D(n27961), .Y(n34559)
         );
  AOI22X1 U29011 ( .A(n33809), .B(n34561), .C(n34015), .D(n34562), .Y(n34557)
         );
  AOI22X1 U29012 ( .A(n34424), .B(n26028), .C(n34563), .D(n26260), .Y(n34541)
         );
  AND2X1 U29013 ( .A(n34564), .B(n34565), .Y(n34424) );
  AOI22X1 U29014 ( .A(n25025), .B(n34566), .C(n25026), .D(n34296), .Y(n34565)
         );
  AOI22X1 U29015 ( .A(n26032), .B(n33985), .C(n26530), .D(n34567), .Y(n34564)
         );
  NAND2X1 U29016 ( .A(n34568), .B(n34569), .Y(n33985) );
  AOI22X1 U29017 ( .A(n26662), .B(n25128), .C(n26663), .D(n25147), .Y(n34569)
         );
  AOI22X1 U29018 ( .A(n26038), .B(n25224), .C(n26664), .D(n27961), .Y(n34568)
         );
  AOI22X1 U29019 ( .A(reg_A[18]), .B(n26551), .C(reg_A[21]), .D(n26353), .Y(
        n34540) );
  NAND2X1 U29020 ( .A(n34570), .B(n34571), .Y(result[25]) );
  NOR2X1 U29021 ( .A(n34572), .B(n34573), .Y(n34571) );
  NAND3X1 U29022 ( .A(n34574), .B(n34575), .C(n34576), .Y(n34573) );
  AOI21X1 U29023 ( .A(n34431), .B(n25150), .C(n34577), .Y(n34576) );
  OAI21X1 U29024 ( .A(n25244), .B(n26418), .C(n34578), .Y(n34577) );
  OAI21X1 U29025 ( .A(n34579), .B(n34580), .C(n25188), .Y(n34578) );
  OAI21X1 U29026 ( .A(n29305), .B(n34581), .C(n34582), .Y(n34580) );
  INVX1 U29027 ( .A(n34583), .Y(n34582) );
  MUX2X1 U29028 ( .B(n34397), .A(n34485), .S(reg_B[30]), .Y(n34583) );
  OAI21X1 U29029 ( .A(reg_B[29]), .B(n34228), .C(n34584), .Y(n34397) );
  AOI21X1 U29030 ( .A(n34190), .B(n34585), .C(n34399), .Y(n34584) );
  AND2X1 U29031 ( .A(n34188), .B(n25250), .Y(n34399) );
  INVX1 U29032 ( .A(n34229), .Y(n34585) );
  MUX2X1 U29033 ( .B(n25232), .A(n30587), .S(reg_B[31]), .Y(n34229) );
  MUX2X1 U29034 ( .B(n34492), .A(n34586), .S(reg_B[31]), .Y(n34228) );
  MUX2X1 U29035 ( .B(reg_A[24]), .A(reg_A[16]), .S(reg_B[28]), .Y(n34586) );
  MUX2X1 U29036 ( .B(reg_A[17]), .A(reg_A[25]), .S(n34493), .Y(n34492) );
  OAI22X1 U29037 ( .A(n25264), .B(n34587), .C(n34588), .D(n34589), .Y(n34579)
         );
  INVX1 U29038 ( .A(n33863), .Y(n34588) );
  MUX2X1 U29039 ( .B(n26714), .A(n25230), .S(reg_B[31]), .Y(n33863) );
  AND2X1 U29040 ( .A(n34590), .B(n34591), .Y(n34431) );
  AOI22X1 U29041 ( .A(n26859), .B(n30587), .C(n26860), .D(n25232), .Y(n34591)
         );
  AOI22X1 U29042 ( .A(n26455), .B(n25250), .C(n34160), .D(n26452), .Y(n34590)
         );
  OAI21X1 U29043 ( .A(reg_A[16]), .B(n26861), .C(n34592), .Y(n34160) );
  AOI22X1 U29044 ( .A(n34515), .B(n26863), .C(n26462), .D(n27962), .Y(n34592)
         );
  MUX2X1 U29045 ( .B(reg_A[17]), .A(reg_A[25]), .S(n26596), .Y(n34515) );
  AOI22X1 U29046 ( .A(n34470), .B(n25166), .C(n34593), .D(n34191), .Y(n34575)
         );
  INVX1 U29047 ( .A(n34594), .Y(n34593) );
  AOI22X1 U29048 ( .A(n25203), .B(n34595), .C(n34596), .D(n25104), .Y(n34574)
         );
  OAI21X1 U29049 ( .A(n26895), .B(n25239), .C(n34597), .Y(n34595) );
  AOI22X1 U29050 ( .A(reg_A[31]), .B(n34598), .C(reg_A[30]), .D(n34599), .Y(
        n34597) );
  OR2X1 U29051 ( .A(n34600), .B(n34601), .Y(n34572) );
  NAND2X1 U29052 ( .A(n34602), .B(n34603), .Y(n34601) );
  AOI22X1 U29053 ( .A(reg_A[24]), .B(n34604), .C(reg_A[25]), .D(n34605), .Y(
        n34603) );
  OAI21X1 U29054 ( .A(n28213), .B(n33915), .C(n26569), .Y(n34605) );
  INVX1 U29055 ( .A(n26450), .Y(n26569) );
  INVX1 U29056 ( .A(n29315), .Y(n28213) );
  OAI21X1 U29057 ( .A(n33977), .B(n26151), .C(n28870), .Y(n34604) );
  NOR2X1 U29058 ( .A(n34606), .B(n32880), .Y(n28870) );
  AOI22X1 U29059 ( .A(n25170), .B(n34607), .C(n34608), .D(n25109), .Y(n34602)
         );
  OAI21X1 U29060 ( .A(n34521), .B(n32935), .C(n34609), .Y(n34607) );
  AOI21X1 U29061 ( .A(n34519), .B(n34610), .C(n34611), .Y(n34609) );
  AOI21X1 U29062 ( .A(n34612), .B(n34613), .C(n25415), .Y(n34611) );
  AOI22X1 U29063 ( .A(n25156), .B(n34504), .C(n25142), .D(n34500), .Y(n34613)
         );
  OAI21X1 U29064 ( .A(n25232), .B(n34009), .C(n34614), .Y(n34504) );
  AOI22X1 U29065 ( .A(n34180), .B(reg_A[17]), .C(n34189), .D(reg_A[25]), .Y(
        n34614) );
  AOI22X1 U29066 ( .A(n25258), .B(n34501), .C(n26761), .D(n34615), .Y(n34612)
         );
  AND2X1 U29067 ( .A(n34616), .B(n34617), .Y(n34521) );
  AOI22X1 U29068 ( .A(n32934), .B(n33920), .C(n34000), .D(n34181), .Y(n34617)
         );
  NAND2X1 U29069 ( .A(n34618), .B(n34619), .Y(n33920) );
  AOI22X1 U29070 ( .A(n33922), .B(reg_A[1]), .C(n33923), .D(reg_A[9]), .Y(
        n34619) );
  AOI22X1 U29071 ( .A(reg_A[17]), .B(n33919), .C(reg_A[25]), .D(n32933), .Y(
        n34618) );
  AOI22X1 U29072 ( .A(n33809), .B(n34409), .C(n34015), .D(n34620), .Y(n34616)
         );
  NAND3X1 U29073 ( .A(n34621), .B(n34327), .C(n34622), .Y(n34600) );
  AOI22X1 U29074 ( .A(reg_A[18]), .B(n34623), .C(reg_A[19]), .D(n34624), .Y(
        n34622) );
  OAI21X1 U29075 ( .A(n26864), .B(n25745), .C(n34625), .Y(n34624) );
  OAI21X1 U29076 ( .A(n26864), .B(n26936), .C(n26328), .Y(n34623) );
  NAND2X1 U29077 ( .A(n34626), .B(reg_B[29]), .Y(n34327) );
  OAI21X1 U29078 ( .A(n26866), .B(n26346), .C(reg_A[16]), .Y(n34621) );
  NOR2X1 U29079 ( .A(n34627), .B(n34628), .Y(n34570) );
  NAND3X1 U29080 ( .A(n34629), .B(n34630), .C(n34631), .Y(n34628) );
  AOI21X1 U29081 ( .A(n34626), .B(n25262), .C(n34632), .Y(n34631) );
  OAI22X1 U29082 ( .A(n25147), .B(n26625), .C(n25206), .D(n26917), .Y(n34632)
         );
  INVX1 U29083 ( .A(n33991), .Y(n34626) );
  NAND2X1 U29084 ( .A(reg_A[24]), .B(n26504), .Y(n33991) );
  AOI22X1 U29085 ( .A(reg_A[20]), .B(n26353), .C(reg_A[22]), .D(n26472), .Y(
        n34630) );
  AOI22X1 U29086 ( .A(reg_A[23]), .B(n34633), .C(n26627), .D(reg_A[14]), .Y(
        n34629) );
  NAND3X1 U29087 ( .A(n34634), .B(n34635), .C(n34636), .Y(n34627) );
  NOR2X1 U29088 ( .A(n34637), .B(n34638), .Y(n34636) );
  OAI21X1 U29089 ( .A(n33964), .B(n34532), .C(n34639), .Y(n34638) );
  OAI21X1 U29090 ( .A(n34640), .B(n34641), .C(n25840), .Y(n34639) );
  NAND3X1 U29091 ( .A(n34642), .B(n34643), .C(n34644), .Y(n34641) );
  AOI21X1 U29092 ( .A(n25325), .B(reg_A[12]), .C(n34645), .Y(n34644) );
  OAI22X1 U29093 ( .A(n27967), .B(n25475), .C(n29279), .D(n25219), .Y(n34645)
         );
  AOI22X1 U29094 ( .A(n25257), .B(reg_A[4]), .C(n25857), .D(reg_A[0]), .Y(
        n34643) );
  AOI22X1 U29095 ( .A(n25647), .B(reg_A[1]), .C(reg_A[24]), .D(n25135), .Y(
        n34642) );
  NAND3X1 U29096 ( .A(n34646), .B(n34647), .C(n34648), .Y(n34640) );
  AOI21X1 U29097 ( .A(n25339), .B(reg_A[5]), .C(n34649), .Y(n34648) );
  OAI22X1 U29098 ( .A(n25128), .B(n25491), .C(n25130), .D(n25492), .Y(n34649)
         );
  AOI22X1 U29099 ( .A(n25246), .B(reg_A[8]), .C(n25247), .D(reg_A[9]), .Y(
        n34647) );
  AOI22X1 U29100 ( .A(n25487), .B(reg_A[6]), .C(n25241), .D(reg_A[7]), .Y(
        n34646) );
  NAND2X1 U29101 ( .A(n34650), .B(n34651), .Y(n34532) );
  AOI22X1 U29102 ( .A(n32934), .B(n34216), .C(n34000), .D(n34466), .Y(n34651)
         );
  NAND2X1 U29103 ( .A(n34652), .B(n34653), .Y(n34216) );
  AOI22X1 U29104 ( .A(n33922), .B(n25177), .C(n33923), .D(n25146), .Y(n34653)
         );
  AOI22X1 U29105 ( .A(n33919), .B(n27953), .C(n32933), .D(n27960), .Y(n34652)
         );
  AOI22X1 U29106 ( .A(n33809), .B(n34467), .C(n34015), .D(n34654), .Y(n34650)
         );
  OAI22X1 U29107 ( .A(n27961), .B(n26136), .C(n32918), .D(n26812), .Y(n34637)
         );
  AOI22X1 U29108 ( .A(reg_A[21]), .B(n26636), .C(n34563), .D(n26028), .Y(
        n34635) );
  AND2X1 U29109 ( .A(n34655), .B(n34656), .Y(n34563) );
  AOI22X1 U29110 ( .A(n25025), .B(n34428), .C(n25026), .D(n34427), .Y(n34656)
         );
  AOI22X1 U29111 ( .A(n26032), .B(n34205), .C(n26530), .D(n34657), .Y(n34655)
         );
  NAND2X1 U29112 ( .A(n34658), .B(n34659), .Y(n34205) );
  AOI22X1 U29113 ( .A(n26662), .B(n25177), .C(n26663), .D(n25146), .Y(n34659)
         );
  AOI22X1 U29114 ( .A(n26038), .B(n27953), .C(n26664), .D(n27960), .Y(n34658)
         );
  AOI22X1 U29115 ( .A(n34660), .B(n26260), .C(reg_A[17]), .D(n26551), .Y(
        n34634) );
  NAND3X1 U29116 ( .A(n34661), .B(n34662), .C(n34663), .Y(result[24]) );
  NOR2X1 U29117 ( .A(n34664), .B(n34665), .Y(n34663) );
  NAND3X1 U29118 ( .A(n34666), .B(n34667), .C(n34668), .Y(n34665) );
  AOI22X1 U29119 ( .A(n25918), .B(n34669), .C(n25730), .D(n34670), .Y(n34668)
         );
  NAND3X1 U29120 ( .A(n34671), .B(n34672), .C(n34673), .Y(n34670) );
  NOR2X1 U29121 ( .A(n34674), .B(n34675), .Y(n34673) );
  OAI22X1 U29122 ( .A(n25061), .B(n29286), .C(n27961), .D(n25746), .Y(n34675)
         );
  OAI22X1 U29123 ( .A(n25747), .B(n32918), .C(n25748), .D(n27960), .Y(n34674)
         );
  AOI22X1 U29124 ( .A(n25613), .B(reg_A[31]), .C(n25749), .D(reg_A[28]), .Y(
        n34672) );
  AOI22X1 U29125 ( .A(n25750), .B(reg_A[29]), .C(reg_A[24]), .D(n26924), .Y(
        n34671) );
  NAND3X1 U29126 ( .A(n34676), .B(n34677), .C(n34678), .Y(n34669) );
  NOR2X1 U29127 ( .A(n34679), .B(n34680), .Y(n34678) );
  OAI22X1 U29128 ( .A(n26936), .B(n27953), .C(n25745), .D(n25224), .Y(n34680)
         );
  OAI21X1 U29129 ( .A(n25062), .B(n25230), .C(n34681), .Y(n34679) );
  AOI22X1 U29130 ( .A(reg_A[23]), .B(n26803), .C(reg_A[21]), .D(n26804), .Y(
        n34681) );
  AOI22X1 U29131 ( .A(reg_A[20]), .B(n25749), .C(reg_A[19]), .D(n25750), .Y(
        n34677) );
  AOI22X1 U29132 ( .A(n25615), .B(reg_A[16]), .C(reg_A[24]), .D(n26924), .Y(
        n34676) );
  OAI21X1 U29133 ( .A(n34682), .B(n34683), .C(n26928), .Y(n34667) );
  NAND2X1 U29134 ( .A(n34684), .B(n34685), .Y(n34683) );
  AOI22X1 U29135 ( .A(n26002), .B(reg_A[31]), .C(n26003), .D(reg_A[28]), .Y(
        n34685) );
  AOI22X1 U29136 ( .A(n25751), .B(reg_A[29]), .C(reg_A[24]), .D(n26004), .Y(
        n34684) );
  NAND2X1 U29137 ( .A(n34686), .B(n34687), .Y(n34682) );
  AOI22X1 U29138 ( .A(reg_A[25]), .B(n26007), .C(reg_A[27]), .D(n26008), .Y(
        n34687) );
  AOI22X1 U29139 ( .A(n26009), .B(reg_A[26]), .C(reg_A[30]), .D(n26010), .Y(
        n34686) );
  AOI22X1 U29140 ( .A(n26519), .B(reg_A[12]), .C(n26349), .D(reg_A[9]), .Y(
        n34666) );
  NAND2X1 U29141 ( .A(n34688), .B(n34689), .Y(n34664) );
  AOI21X1 U29142 ( .A(n34660), .B(n26028), .C(n34690), .Y(n34689) );
  OAI21X1 U29143 ( .A(n34691), .B(n31828), .C(n34692), .Y(n34690) );
  OAI21X1 U29144 ( .A(n34693), .B(n34694), .C(n25840), .Y(n34692) );
  NAND3X1 U29145 ( .A(n34695), .B(n34696), .C(n34697), .Y(n34694) );
  NOR2X1 U29146 ( .A(n34698), .B(n34699), .Y(n34697) );
  OAI21X1 U29147 ( .A(n29279), .B(n25223), .C(n34700), .Y(n34699) );
  AOI22X1 U29148 ( .A(reg_A[20]), .B(n25073), .C(reg_A[19]), .D(n25123), .Y(
        n34700) );
  OAI21X1 U29149 ( .A(n25030), .B(n27953), .C(n34701), .Y(n34698) );
  AOI22X1 U29150 ( .A(reg_A[22]), .B(n25252), .C(reg_A[18]), .D(n25253), .Y(
        n34701) );
  AOI21X1 U29151 ( .A(n25234), .B(reg_A[10]), .C(n34702), .Y(n34696) );
  OAI22X1 U29152 ( .A(n25208), .B(n25219), .C(n25250), .D(n25467), .Y(n34702)
         );
  AOI22X1 U29153 ( .A(n25325), .B(reg_A[11]), .C(n25125), .D(reg_A[24]), .Y(
        n34695) );
  NAND3X1 U29154 ( .A(n34703), .B(n34704), .C(n34705), .Y(n34693) );
  NOR2X1 U29155 ( .A(n34706), .B(n34707), .Y(n34705) );
  OAI21X1 U29156 ( .A(n25177), .B(n25491), .C(n34708), .Y(n34707) );
  AOI22X1 U29157 ( .A(n25241), .B(reg_A[6]), .C(n25242), .D(reg_A[2]), .Y(
        n34708) );
  OAI21X1 U29158 ( .A(n29265), .B(n25243), .C(n34709), .Y(n34706) );
  AOI22X1 U29159 ( .A(n25246), .B(reg_A[7]), .C(n25247), .D(reg_A[8]), .Y(
        n34709) );
  AOI21X1 U29160 ( .A(n25647), .B(reg_A[0]), .C(n34710), .Y(n34704) );
  OAI22X1 U29161 ( .A(n25130), .B(n26719), .C(n30569), .D(n25238), .Y(n34710)
         );
  AOI22X1 U29162 ( .A(reg_A[23]), .B(n25135), .C(reg_A[21]), .D(n25136), .Y(
        n34703) );
  INVX1 U29163 ( .A(n34610), .Y(n34691) );
  NAND2X1 U29164 ( .A(n34711), .B(n34712), .Y(n34610) );
  AOI22X1 U29165 ( .A(n32934), .B(n34347), .C(n34000), .D(n34341), .Y(n34712)
         );
  NAND2X1 U29166 ( .A(n34713), .B(n34714), .Y(n34347) );
  AOI22X1 U29167 ( .A(n33922), .B(reg_A[0]), .C(n33923), .D(reg_A[8]), .Y(
        n34714) );
  AOI22X1 U29168 ( .A(reg_A[16]), .B(n33919), .C(reg_A[24]), .D(n32933), .Y(
        n34713) );
  AOI22X1 U29169 ( .A(n33809), .B(n34528), .C(n34015), .D(n34715), .Y(n34711)
         );
  AND2X1 U29170 ( .A(n34716), .B(n34717), .Y(n34660) );
  AOI22X1 U29171 ( .A(n25025), .B(n34567), .C(n25026), .D(n34566), .Y(n34717)
         );
  AOI22X1 U29172 ( .A(n26032), .B(n34296), .C(n26530), .D(n34718), .Y(n34716)
         );
  OR2X1 U29173 ( .A(n34719), .B(n34720), .Y(n34296) );
  OAI22X1 U29174 ( .A(reg_A[24]), .B(n25063), .C(reg_A[16]), .D(n26981), .Y(
        n34720) );
  OAI21X1 U29175 ( .A(reg_A[8]), .B(n26982), .C(n34721), .Y(n34719) );
  AOI21X1 U29176 ( .A(n26627), .B(reg_A[13]), .C(n34722), .Y(n34688) );
  OAI22X1 U29177 ( .A(n25250), .B(n26985), .C(n26012), .D(n34723), .Y(n34722)
         );
  NOR2X1 U29178 ( .A(n34724), .B(n34725), .Y(n34662) );
  OAI21X1 U29179 ( .A(n34726), .B(n34495), .C(n34727), .Y(n34725) );
  AOI22X1 U29180 ( .A(n34728), .B(n27008), .C(n26267), .D(n34729), .Y(n34727)
         );
  NAND2X1 U29181 ( .A(n34730), .B(n34731), .Y(n34729) );
  AOI22X1 U29182 ( .A(n25156), .B(n34500), .C(n25142), .D(n34501), .Y(n34731)
         );
  OAI21X1 U29183 ( .A(n30587), .B(n34009), .C(n34732), .Y(n34500) );
  AOI22X1 U29184 ( .A(n34180), .B(reg_A[16]), .C(n34189), .D(reg_A[24]), .Y(
        n34732) );
  AOI22X1 U29185 ( .A(n25258), .B(n34615), .C(n26761), .D(n34733), .Y(n34730)
         );
  INVX1 U29186 ( .A(n34734), .Y(n34733) );
  INVX1 U29187 ( .A(n34356), .Y(n34728) );
  NAND2X1 U29188 ( .A(n34735), .B(n34736), .Y(n34356) );
  AOI22X1 U29189 ( .A(n26601), .B(n25230), .C(n26602), .D(n25232), .Y(n34736)
         );
  AOI22X1 U29190 ( .A(n27012), .B(n27962), .C(n26597), .D(n26714), .Y(n34735)
         );
  INVX1 U29191 ( .A(n34596), .Y(n34495) );
  OAI21X1 U29192 ( .A(n34737), .B(n34738), .C(n34285), .Y(n34596) );
  NAND3X1 U29193 ( .A(n33874), .B(n33955), .C(n25382), .Y(n34285) );
  NAND2X1 U29194 ( .A(n25382), .B(n34189), .Y(n34738) );
  OAI21X1 U29195 ( .A(n34387), .B(n34739), .C(n34740), .Y(n34724) );
  AOI22X1 U29196 ( .A(reg_A[24]), .B(n34741), .C(n34608), .D(n26777), .Y(
        n34740) );
  INVX1 U29197 ( .A(n34511), .Y(n34608) );
  NAND2X1 U29198 ( .A(n25382), .B(n34742), .Y(n34511) );
  OAI22X1 U29199 ( .A(n34009), .B(n34737), .C(n33808), .D(n33955), .Y(n34742)
         );
  INVX1 U29200 ( .A(n33874), .Y(n33808) );
  OAI21X1 U29201 ( .A(reg_B[28]), .B(n25415), .C(n26999), .Y(n33874) );
  OAI21X1 U29202 ( .A(n26151), .B(n33915), .C(n34743), .Y(n34741) );
  INVX1 U29203 ( .A(n27032), .Y(n34743) );
  NOR2X1 U29204 ( .A(n34744), .B(n34745), .Y(n34661) );
  OAI22X1 U29205 ( .A(n34746), .B(n30547), .C(n33964), .D(n34594), .Y(n34745)
         );
  NAND2X1 U29206 ( .A(n34747), .B(n34748), .Y(n34594) );
  AOI22X1 U29207 ( .A(n32934), .B(n34305), .C(n34000), .D(n34561), .Y(n34748)
         );
  OR2X1 U29208 ( .A(n34749), .B(n34750), .Y(n34305) );
  OAI22X1 U29209 ( .A(reg_A[24]), .B(n33807), .C(reg_A[16]), .D(n34465), .Y(
        n34750) );
  OAI21X1 U29210 ( .A(reg_A[8]), .B(n34751), .C(n34752), .Y(n34749) );
  AOI22X1 U29211 ( .A(n33809), .B(n34562), .C(n34015), .D(n34753), .Y(n34747)
         );
  OAI21X1 U29212 ( .A(n26420), .B(n34357), .C(n34754), .Y(n34744) );
  AOI22X1 U29213 ( .A(n25188), .B(n34755), .C(n25310), .D(n34756), .Y(n34754)
         );
  NAND3X1 U29214 ( .A(n34757), .B(n34758), .C(n34759), .Y(n34756) );
  AOI21X1 U29215 ( .A(n25123), .B(reg_A[29]), .C(n34760), .Y(n34759) );
  OAI22X1 U29216 ( .A(n25244), .B(n26431), .C(n27954), .D(n25129), .Y(n34760)
         );
  AOI22X1 U29217 ( .A(n25135), .B(reg_A[25]), .C(n25136), .D(reg_A[27]), .Y(
        n34758) );
  AOI22X1 U29218 ( .A(n25252), .B(reg_A[26]), .C(n25253), .D(reg_A[30]), .Y(
        n34757) );
  OAI21X1 U29219 ( .A(n34230), .B(n34314), .C(n34761), .Y(n34755) );
  INVX1 U29220 ( .A(n34762), .Y(n34761) );
  OAI21X1 U29221 ( .A(n34315), .B(n34009), .C(n34485), .Y(n34762) );
  NAND2X1 U29222 ( .A(n34763), .B(n34764), .Y(n34315) );
  AOI22X1 U29223 ( .A(n25156), .B(n30587), .C(n25142), .D(n25220), .Y(n34764)
         );
  AOI22X1 U29224 ( .A(n25258), .B(n25224), .C(n26761), .D(n27953), .Y(n34763)
         );
  NAND2X1 U29225 ( .A(n34765), .B(n34766), .Y(n34314) );
  AOI22X1 U29226 ( .A(n25156), .B(n27962), .C(n25142), .D(n26714), .Y(n34766)
         );
  AOI22X1 U29227 ( .A(n25258), .B(n25230), .C(n26761), .D(n25232), .Y(n34765)
         );
  OR2X1 U29228 ( .A(n34767), .B(n34768), .Y(result[23]) );
  NAND3X1 U29229 ( .A(n34769), .B(n34770), .C(n34771), .Y(n34768) );
  NOR2X1 U29230 ( .A(n34772), .B(n34773), .Y(n34771) );
  OAI22X1 U29231 ( .A(n26525), .B(n34723), .C(n33964), .D(n34739), .Y(n34773)
         );
  NAND2X1 U29232 ( .A(n34774), .B(n34775), .Y(n34739) );
  AOI22X1 U29233 ( .A(n32934), .B(n34466), .C(n34000), .D(n34467), .Y(n34775)
         );
  INVX1 U29234 ( .A(n34210), .Y(n34466) );
  NOR2X1 U29235 ( .A(n34776), .B(n34777), .Y(n34210) );
  OAI22X1 U29236 ( .A(reg_A[23]), .B(n33807), .C(reg_A[15]), .D(n34465), .Y(
        n34777) );
  OAI21X1 U29237 ( .A(reg_A[7]), .B(n34751), .C(n34752), .Y(n34776) );
  AOI22X1 U29238 ( .A(n33809), .B(n34654), .C(n34015), .D(n34778), .Y(n34774)
         );
  INVX1 U29239 ( .A(n34779), .Y(n34778) );
  INVX1 U29240 ( .A(n34780), .Y(n34654) );
  NAND2X1 U29241 ( .A(n34781), .B(n34782), .Y(n34723) );
  AOI22X1 U29242 ( .A(n25025), .B(n34657), .C(n25026), .D(n34428), .Y(n34782)
         );
  INVX1 U29243 ( .A(n34783), .Y(n34657) );
  AOI22X1 U29244 ( .A(n26032), .B(n34427), .C(n26530), .D(n34784), .Y(n34781)
         );
  INVX1 U29245 ( .A(n34201), .Y(n34427) );
  NOR2X1 U29246 ( .A(n34785), .B(n34786), .Y(n34201) );
  OAI22X1 U29247 ( .A(reg_A[23]), .B(n25063), .C(reg_A[15]), .D(n26981), .Y(
        n34786) );
  OAI21X1 U29248 ( .A(reg_A[7]), .B(n26982), .C(n34721), .Y(n34785) );
  OAI21X1 U29249 ( .A(n25945), .B(n34787), .C(n34788), .Y(n34772) );
  AOI22X1 U29250 ( .A(n27132), .B(reg_A[19]), .C(reg_A[16]), .D(n27051), .Y(
        n34788) );
  AOI22X1 U29251 ( .A(n34789), .B(n26260), .C(n25730), .D(n34790), .Y(n34770)
         );
  NAND3X1 U29252 ( .A(n34791), .B(n34792), .C(n34793), .Y(n34790) );
  NOR2X1 U29253 ( .A(n34794), .B(n34795), .Y(n34793) );
  OAI22X1 U29254 ( .A(n29286), .B(n26936), .C(n25745), .D(n25239), .Y(n34795)
         );
  OAI21X1 U29255 ( .A(n27960), .B(n25746), .C(n34796), .Y(n34794) );
  AOI22X1 U29256 ( .A(reg_A[24]), .B(n26803), .C(n26804), .D(reg_A[26]), .Y(
        n34796) );
  AOI22X1 U29257 ( .A(n25749), .B(reg_A[27]), .C(n25750), .D(reg_A[28]), .Y(
        n34792) );
  AOI22X1 U29258 ( .A(n25615), .B(reg_A[31]), .C(reg_A[23]), .D(n26924), .Y(
        n34791) );
  INVX1 U29259 ( .A(n34797), .Y(n34789) );
  AOI22X1 U29260 ( .A(n34798), .B(n28037), .C(n25310), .D(n34799), .Y(n34769)
         );
  NAND3X1 U29261 ( .A(n34800), .B(n34801), .C(n34802), .Y(n34799) );
  NOR2X1 U29262 ( .A(n34803), .B(n34804), .Y(n34802) );
  OAI22X1 U29263 ( .A(n29286), .B(n25129), .C(n25239), .D(n25131), .Y(n34804)
         );
  OAI21X1 U29264 ( .A(n27960), .B(n25133), .C(n34805), .Y(n34803) );
  AOI22X1 U29265 ( .A(reg_A[24]), .B(n25135), .C(n25136), .D(reg_A[26]), .Y(
        n34805) );
  AOI22X1 U29266 ( .A(n25075), .B(reg_A[27]), .C(n25123), .D(reg_A[28]), .Y(
        n34801) );
  AOI22X1 U29267 ( .A(n25124), .B(reg_A[31]), .C(n25125), .D(reg_A[23]), .Y(
        n34800) );
  OAI21X1 U29268 ( .A(n34806), .B(n34009), .C(n34807), .Y(n28037) );
  AOI22X1 U29269 ( .A(n33806), .B(reg_B[28]), .C(n34189), .D(n34808), .Y(
        n34807) );
  INVX1 U29270 ( .A(n34809), .Y(n34806) );
  NAND2X1 U29271 ( .A(n34810), .B(n34811), .Y(n34767) );
  NOR2X1 U29272 ( .A(n34812), .B(n34813), .Y(n34811) );
  OAI21X1 U29273 ( .A(n34814), .B(n26714), .C(n34815), .Y(n34813) );
  OAI21X1 U29274 ( .A(n34816), .B(n34817), .C(n25170), .Y(n34815) );
  OAI21X1 U29275 ( .A(n34746), .B(n32935), .C(n34818), .Y(n34817) );
  MUX2X1 U29276 ( .B(n34819), .A(n34820), .S(reg_B[23]), .Y(n34818) );
  NOR2X1 U29277 ( .A(n34821), .B(n26999), .Y(n34820) );
  OAI21X1 U29278 ( .A(n25232), .B(n34822), .C(n34823), .Y(n34819) );
  AOI22X1 U29279 ( .A(n34824), .B(n34825), .C(n34826), .D(reg_A[23]), .Y(
        n34823) );
  MUX2X1 U29280 ( .B(n25220), .A(n27953), .S(reg_B[22]), .Y(n34824) );
  AND2X1 U29281 ( .A(n34827), .B(n34828), .Y(n34746) );
  AOI22X1 U29282 ( .A(n32934), .B(n34181), .C(n34000), .D(n34409), .Y(n34828)
         );
  OAI21X1 U29283 ( .A(n33807), .B(n26714), .C(n34829), .Y(n34181) );
  AOI22X1 U29284 ( .A(n33923), .B(reg_A[7]), .C(reg_A[15]), .D(n33919), .Y(
        n34829) );
  AOI22X1 U29285 ( .A(n33809), .B(n34620), .C(n34015), .D(n34830), .Y(n34827)
         );
  OAI21X1 U29286 ( .A(n34831), .B(n31806), .C(n34832), .Y(n34816) );
  OAI21X1 U29287 ( .A(n34833), .B(n34834), .C(n25604), .Y(n34832) );
  NOR2X1 U29288 ( .A(n34835), .B(n25264), .Y(n34833) );
  INVX1 U29289 ( .A(n34836), .Y(n34814) );
  OAI21X1 U29290 ( .A(n34837), .B(n25087), .C(n34838), .Y(n34836) );
  NAND3X1 U29291 ( .A(n34839), .B(n34840), .C(n34841), .Y(n34812) );
  OAI21X1 U29292 ( .A(n34834), .B(n34842), .C(n25188), .Y(n34841) );
  OAI21X1 U29293 ( .A(n34843), .B(n25264), .C(n34485), .Y(n34842) );
  AOI21X1 U29294 ( .A(reg_A[16]), .B(reg_B[29]), .C(n34844), .Y(n34843) );
  OAI21X1 U29295 ( .A(n34734), .B(n29305), .C(n34845), .Y(n34834) );
  AOI22X1 U29296 ( .A(n25156), .B(n34501), .C(n25142), .D(n34615), .Y(n34845)
         );
  OAI21X1 U29297 ( .A(n26714), .B(n34230), .C(n34581), .Y(n34501) );
  NAND2X1 U29298 ( .A(n34190), .B(reg_A[19]), .Y(n34581) );
  OAI21X1 U29299 ( .A(n34846), .B(n34847), .C(n25840), .Y(n34840) );
  NAND2X1 U29300 ( .A(n34848), .B(n34849), .Y(n34847) );
  NOR2X1 U29301 ( .A(n34850), .B(n34851), .Y(n34849) );
  OAI21X1 U29302 ( .A(n26714), .B(n25043), .C(n34852), .Y(n34851) );
  AOI22X1 U29303 ( .A(reg_A[22]), .B(n25135), .C(reg_A[21]), .D(n25252), .Y(
        n34852) );
  OAI21X1 U29304 ( .A(n25028), .B(n25224), .C(n34853), .Y(n34850) );
  AOI22X1 U29305 ( .A(reg_A[20]), .B(n25136), .C(reg_A[19]), .D(n25068), .Y(
        n34853) );
  NOR2X1 U29306 ( .A(n34854), .B(n34855), .Y(n34848) );
  OAI21X1 U29307 ( .A(n29279), .B(n25467), .C(n34856), .Y(n34855) );
  AOI22X1 U29308 ( .A(reg_A[17]), .B(n25253), .C(reg_A[16]), .D(n25628), .Y(
        n34856) );
  OAI21X1 U29309 ( .A(n25206), .B(n25219), .C(n34857), .Y(n34854) );
  AOI22X1 U29310 ( .A(n25629), .B(reg_A[14]), .C(n25222), .D(reg_A[12]), .Y(
        n34857) );
  NAND2X1 U29311 ( .A(n34858), .B(n34859), .Y(n34846) );
  NOR2X1 U29312 ( .A(n34860), .B(n34861), .Y(n34859) );
  OAI21X1 U29313 ( .A(n25147), .B(n25229), .C(n34862), .Y(n34861) );
  AOI22X1 U29314 ( .A(n25234), .B(reg_A[9]), .C(n25635), .D(reg_A[11]), .Y(
        n34862) );
  OAI21X1 U29315 ( .A(n26701), .B(n25482), .C(n34863), .Y(n34860) );
  AOI22X1 U29316 ( .A(n25246), .B(reg_A[6]), .C(n25247), .D(reg_A[7]), .Y(
        n34863) );
  NOR2X1 U29317 ( .A(n34864), .B(n34865), .Y(n34858) );
  OAI21X1 U29318 ( .A(n25130), .B(n25238), .C(n34866), .Y(n34865) );
  AOI22X1 U29319 ( .A(n25487), .B(reg_A[4]), .C(n25241), .D(reg_A[5]), .Y(
        n34866) );
  OAI21X1 U29320 ( .A(n25128), .B(n26719), .C(n34867), .Y(n34864) );
  AOI22X1 U29321 ( .A(n25242), .B(reg_A[1]), .C(n25338), .D(reg_A[0]), .Y(
        n34867) );
  OAI21X1 U29322 ( .A(n34868), .B(n34869), .C(n27067), .Y(n34839) );
  OAI21X1 U29323 ( .A(n25060), .B(n26714), .C(n34870), .Y(n34869) );
  AOI22X1 U29324 ( .A(reg_A[19]), .B(n25749), .C(reg_A[18]), .D(n25750), .Y(
        n34870) );
  NAND2X1 U29325 ( .A(n34871), .B(n34872), .Y(n34868) );
  AOI22X1 U29326 ( .A(reg_A[22]), .B(n26803), .C(reg_A[20]), .D(n26804), .Y(
        n34872) );
  AOI22X1 U29327 ( .A(reg_A[21]), .B(n26927), .C(reg_A[17]), .D(n26878), .Y(
        n34871) );
  NOR2X1 U29328 ( .A(n34873), .B(n34874), .Y(n34810) );
  OAI21X1 U29329 ( .A(n34875), .B(n25342), .C(n34876), .Y(n34874) );
  OAI21X1 U29330 ( .A(n34877), .B(n34878), .C(n25999), .Y(n34876) );
  OAI22X1 U29331 ( .A(n25754), .B(n27953), .C(n31144), .D(n25232), .Y(n34878)
         );
  OAI22X1 U29332 ( .A(n30090), .B(n30587), .C(n27925), .D(n25230), .Y(n34877)
         );
  NOR2X1 U29333 ( .A(n34879), .B(n34880), .Y(n34875) );
  OAI21X1 U29334 ( .A(n34881), .B(n34882), .C(n34883), .Y(n34880) );
  NAND3X1 U29335 ( .A(reg_B[21]), .B(reg_A[19]), .C(n34884), .Y(n34883) );
  INVX1 U29336 ( .A(n34885), .Y(n34882) );
  MUX2X1 U29337 ( .B(n34886), .A(n34887), .S(reg_B[23]), .Y(n34879) );
  NAND2X1 U29338 ( .A(n34888), .B(reg_A[23]), .Y(n34886) );
  OAI21X1 U29339 ( .A(n25224), .B(n27108), .C(n34889), .Y(n34873) );
  AOI22X1 U29340 ( .A(n34470), .B(n27110), .C(n34890), .D(n34191), .Y(n34889)
         );
  MUX2X1 U29341 ( .B(n26714), .A(n25230), .S(reg_B[4]), .Y(n34470) );
  NAND3X1 U29342 ( .A(n34891), .B(n34892), .C(n34893), .Y(result[22]) );
  NOR2X1 U29343 ( .A(n34894), .B(n34895), .Y(n34893) );
  NAND3X1 U29344 ( .A(n34896), .B(n34897), .C(n34898), .Y(n34895) );
  AOI21X1 U29345 ( .A(n34020), .B(n34899), .C(n34900), .Y(n34898) );
  OAI22X1 U29346 ( .A(n34901), .B(n34902), .C(n34821), .D(n34903), .Y(n34900)
         );
  AOI21X1 U29347 ( .A(reg_B[21]), .B(n34904), .C(n34905), .Y(n34821) );
  INVX1 U29348 ( .A(n29244), .Y(n34901) );
  OAI21X1 U29349 ( .A(n34906), .B(n34230), .C(n34907), .Y(n29244) );
  AOI22X1 U29350 ( .A(n34180), .B(n34908), .C(n34190), .D(n34909), .Y(n34907)
         );
  AOI22X1 U29351 ( .A(n34910), .B(n34911), .C(n27402), .D(reg_A[23]), .Y(
        n34896) );
  NAND3X1 U29352 ( .A(n34912), .B(n34913), .C(n34914), .Y(n34894) );
  NOR2X1 U29353 ( .A(n34915), .B(n34916), .Y(n34914) );
  OAI22X1 U29354 ( .A(n26012), .B(n34917), .C(n26525), .D(n34797), .Y(n34916)
         );
  NAND2X1 U29355 ( .A(n34918), .B(n34919), .Y(n34797) );
  AOI22X1 U29356 ( .A(n25025), .B(n34718), .C(n25026), .D(n34567), .Y(n34919)
         );
  INVX1 U29357 ( .A(n34920), .Y(n34718) );
  AOI22X1 U29358 ( .A(n26032), .B(n34566), .C(n26530), .D(n34921), .Y(n34918)
         );
  INVX1 U29359 ( .A(n34292), .Y(n34566) );
  NOR2X1 U29360 ( .A(n34922), .B(n34923), .Y(n34292) );
  OAI22X1 U29361 ( .A(reg_A[22]), .B(n25063), .C(reg_A[14]), .D(n26981), .Y(
        n34923) );
  OAI21X1 U29362 ( .A(reg_A[6]), .B(n26982), .C(n34721), .Y(n34922) );
  OAI22X1 U29363 ( .A(n34924), .B(n27953), .C(n34831), .D(n31828), .Y(n34915)
         );
  AND2X1 U29364 ( .A(n34925), .B(n34926), .Y(n34831) );
  AOI22X1 U29365 ( .A(n32934), .B(n34341), .C(n34000), .D(n34528), .Y(n34926)
         );
  OAI21X1 U29366 ( .A(n33807), .B(n25230), .C(n34927), .Y(n34341) );
  AOI22X1 U29367 ( .A(n33923), .B(reg_A[6]), .C(reg_A[14]), .D(n33919), .Y(
        n34927) );
  AOI22X1 U29368 ( .A(n33809), .B(n34715), .C(n34015), .D(n34928), .Y(n34925)
         );
  INVX1 U29369 ( .A(n27256), .Y(n34924) );
  OAI21X1 U29370 ( .A(n34929), .B(n34930), .C(n25310), .Y(n34913) );
  OR2X1 U29371 ( .A(n34931), .B(n34932), .Y(n34930) );
  OAI22X1 U29372 ( .A(n25230), .B(n25228), .C(n29286), .D(n25467), .Y(n34932)
         );
  OAI21X1 U29373 ( .A(n27954), .B(n25223), .C(n34933), .Y(n34931) );
  AOI22X1 U29374 ( .A(n25075), .B(reg_A[26]), .C(n25123), .D(reg_A[27]), .Y(
        n34933) );
  OR2X1 U29375 ( .A(n34934), .B(n34935), .Y(n34929) );
  OAI22X1 U29376 ( .A(n25239), .B(n25129), .C(n25244), .D(n25131), .Y(n34935)
         );
  OAI21X1 U29377 ( .A(n25040), .B(n27962), .C(n34936), .Y(n34934) );
  AOI22X1 U29378 ( .A(reg_A[23]), .B(n25135), .C(n25136), .D(reg_A[25]), .Y(
        n34936) );
  AOI22X1 U29379 ( .A(n26045), .B(n34937), .C(n25730), .D(n34938), .Y(n34912)
         );
  NAND3X1 U29380 ( .A(n34939), .B(n34940), .C(n34941), .Y(n34938) );
  NOR2X1 U29381 ( .A(n34942), .B(n34943), .Y(n34941) );
  OAI22X1 U29382 ( .A(n25239), .B(n26936), .C(n25745), .D(n25244), .Y(n34943)
         );
  OAI21X1 U29383 ( .A(n25062), .B(n27962), .C(n34944), .Y(n34942) );
  AOI22X1 U29384 ( .A(reg_A[23]), .B(n26803), .C(n26804), .D(reg_A[25]), .Y(
        n34944) );
  AOI21X1 U29385 ( .A(n25614), .B(reg_A[31]), .C(n34945), .Y(n34940) );
  OAI22X1 U29386 ( .A(n32918), .B(n26800), .C(n27961), .D(n26801), .Y(n34945)
         );
  AOI22X1 U29387 ( .A(n25615), .B(reg_A[30]), .C(reg_A[22]), .D(n26924), .Y(
        n34939) );
  NAND3X1 U29388 ( .A(n34946), .B(n34947), .C(n34948), .Y(n34937) );
  NOR2X1 U29389 ( .A(n34949), .B(n34950), .Y(n34948) );
  OAI22X1 U29390 ( .A(n27218), .B(n25232), .C(n25207), .D(n27953), .Y(n34950)
         );
  OAI21X1 U29391 ( .A(n27219), .B(n25250), .C(n34951), .Y(n34949) );
  OAI21X1 U29392 ( .A(n34952), .B(n34953), .C(n25044), .Y(n34951) );
  NAND3X1 U29393 ( .A(n34954), .B(n34955), .C(n34956), .Y(n34953) );
  NOR2X1 U29394 ( .A(n34957), .B(n34958), .Y(n34956) );
  OAI21X1 U29395 ( .A(n25255), .B(n25219), .C(n34959), .Y(n34958) );
  AOI22X1 U29396 ( .A(n25124), .B(reg_A[14]), .C(n25222), .D(reg_A[11]), .Y(
        n34959) );
  OAI21X1 U29397 ( .A(n25206), .B(n25223), .C(n34960), .Y(n34957) );
  AOI22X1 U29398 ( .A(reg_A[18]), .B(n25073), .C(reg_A[17]), .D(n25123), .Y(
        n34960) );
  AOI21X1 U29399 ( .A(n25635), .B(reg_A[10]), .C(n34961), .Y(n34955) );
  OAI22X1 U29400 ( .A(n25132), .B(n25482), .C(n26701), .D(n25475), .Y(n34961)
         );
  AOI22X1 U29401 ( .A(n25325), .B(reg_A[9]), .C(n25125), .D(reg_A[22]), .Y(
        n34954) );
  NAND2X1 U29402 ( .A(n34962), .B(n34963), .Y(n34952) );
  NOR2X1 U29403 ( .A(n34964), .B(n34965), .Y(n34963) );
  OAI21X1 U29404 ( .A(n25128), .B(n25238), .C(n34966), .Y(n34965) );
  AOI22X1 U29405 ( .A(n25241), .B(reg_A[4]), .C(n25242), .D(reg_A[0]), .Y(
        n34966) );
  OAI21X1 U29406 ( .A(n25130), .B(n25243), .C(n34967), .Y(n34964) );
  AOI22X1 U29407 ( .A(n25246), .B(reg_A[5]), .C(n25247), .D(reg_A[6]), .Y(
        n34967) );
  NOR2X1 U29408 ( .A(n34968), .B(n34969), .Y(n34962) );
  OAI21X1 U29409 ( .A(n29279), .B(n25129), .C(n34970), .Y(n34969) );
  AOI22X1 U29410 ( .A(reg_A[20]), .B(n25252), .C(reg_A[16]), .D(n25253), .Y(
        n34970) );
  OAI21X1 U29411 ( .A(n25041), .B(n25220), .C(n34971), .Y(n34968) );
  AOI22X1 U29412 ( .A(n25257), .B(reg_A[1]), .C(reg_A[21]), .D(n25135), .Y(
        n34971) );
  AOI22X1 U29413 ( .A(reg_A[19]), .B(n27241), .C(reg_A[18]), .D(n27242), .Y(
        n34947) );
  AOI22X1 U29414 ( .A(reg_A[20]), .B(n27243), .C(reg_A[22]), .D(n25434), .Y(
        n34946) );
  NOR2X1 U29415 ( .A(n34972), .B(n34973), .Y(n34892) );
  OAI21X1 U29416 ( .A(n27190), .B(n33973), .C(n34974), .Y(n34973) );
  AOI22X1 U29417 ( .A(n27204), .B(reg_A[19]), .C(n34975), .D(n34976), .Y(
        n34974) );
  NAND2X1 U29418 ( .A(n34977), .B(n34978), .Y(n33973) );
  AOI22X1 U29419 ( .A(n26601), .B(n30587), .C(n26602), .D(n25220), .Y(n34978)
         );
  AOI22X1 U29420 ( .A(n27012), .B(n25230), .C(n26597), .D(n25232), .Y(n34977)
         );
  NAND2X1 U29421 ( .A(n34979), .B(n34980), .Y(n34972) );
  INVX1 U29422 ( .A(n34981), .Y(n34980) );
  OAI22X1 U29423 ( .A(n34982), .B(n27354), .C(n34983), .D(n25342), .Y(n34981)
         );
  MUX2X1 U29424 ( .B(n34905), .A(n34911), .S(reg_B[23]), .Y(n34983) );
  OAI21X1 U29425 ( .A(n30587), .B(n34984), .C(n34887), .Y(n34905) );
  AOI22X1 U29426 ( .A(reg_A[22]), .B(n34888), .C(reg_A[18]), .D(n34985), .Y(
        n34887) );
  AOI22X1 U29427 ( .A(n34986), .B(reg_B[31]), .C(n34615), .D(n25156), .Y(
        n34982) );
  OAI21X1 U29428 ( .A(n25230), .B(n34230), .C(n34587), .Y(n34615) );
  NAND2X1 U29429 ( .A(n34190), .B(reg_A[18]), .Y(n34587) );
  AOI22X1 U29430 ( .A(n25258), .B(n34987), .C(reg_A[16]), .D(n34988), .Y(
        n34979) );
  OAI21X1 U29431 ( .A(n25032), .B(n29255), .C(n31325), .Y(n34988) );
  INVX1 U29432 ( .A(n27192), .Y(n31325) );
  OAI22X1 U29433 ( .A(n25794), .B(n34989), .C(n34835), .D(n26147), .Y(n34987)
         );
  NOR2X1 U29434 ( .A(n34990), .B(n34991), .Y(n34891) );
  OAI21X1 U29435 ( .A(n27173), .B(n25224), .C(n34992), .Y(n34991) );
  AOI22X1 U29436 ( .A(reg_A[22]), .B(n27184), .C(n34890), .D(n30616), .Y(
        n34992) );
  AND2X1 U29437 ( .A(n34993), .B(n34994), .Y(n34890) );
  AOI22X1 U29438 ( .A(n32934), .B(n34561), .C(n34000), .D(n34562), .Y(n34994)
         );
  INVX1 U29439 ( .A(n34300), .Y(n34561) );
  NOR2X1 U29440 ( .A(n34995), .B(n34996), .Y(n34300) );
  OAI22X1 U29441 ( .A(reg_A[22]), .B(n33807), .C(reg_A[14]), .D(n34465), .Y(
        n34996) );
  OAI21X1 U29442 ( .A(reg_A[6]), .B(n34751), .C(n34752), .Y(n34995) );
  AOI22X1 U29443 ( .A(n34015), .B(n34997), .C(n33809), .D(n34753), .Y(n34993)
         );
  INVX1 U29444 ( .A(n34998), .Y(n34753) );
  NAND2X1 U29445 ( .A(n25795), .B(n34999), .Y(n27184) );
  OAI21X1 U29446 ( .A(n30587), .B(n31351), .C(n35000), .Y(n34990) );
  AOI22X1 U29447 ( .A(n35001), .B(n34191), .C(n27188), .D(reg_A[21]), .Y(
        n35000) );
  INVX1 U29448 ( .A(n34387), .Y(n34191) );
  INVX1 U29449 ( .A(n35002), .Y(n35001) );
  OR2X1 U29450 ( .A(n35003), .B(n35004), .Y(result[21]) );
  NAND3X1 U29451 ( .A(n35005), .B(n35006), .C(n35007), .Y(n35004) );
  NOR2X1 U29452 ( .A(n35008), .B(n35009), .Y(n35007) );
  OAI21X1 U29453 ( .A(n35010), .B(n34902), .C(n35011), .Y(n35009) );
  AOI22X1 U29454 ( .A(n30617), .B(n34899), .C(n35012), .D(n34911), .Y(n35011)
         );
  OAI21X1 U29455 ( .A(n25232), .B(n35013), .C(n35014), .Y(n34911) );
  AOI22X1 U29456 ( .A(n34985), .B(reg_A[17]), .C(n35015), .D(reg_A[19]), .Y(
        n35014) );
  NAND2X1 U29457 ( .A(n35016), .B(n35017), .Y(n34899) );
  AOI22X1 U29458 ( .A(n32934), .B(n34409), .C(n34000), .D(n34620), .Y(n35017)
         );
  OAI21X1 U29459 ( .A(n33807), .B(n25232), .C(n35018), .Y(n34409) );
  AOI22X1 U29460 ( .A(n33923), .B(reg_A[5]), .C(reg_A[13]), .D(n33919), .Y(
        n35018) );
  AOI22X1 U29461 ( .A(n33809), .B(n34830), .C(n34015), .D(n35019), .Y(n35016)
         );
  INVX1 U29462 ( .A(n30645), .Y(n35010) );
  OAI21X1 U29463 ( .A(n35020), .B(n33957), .C(n35021), .Y(n30645) );
  AOI22X1 U29464 ( .A(n34189), .B(n35022), .C(n34190), .D(n25104), .Y(n35021)
         );
  OAI21X1 U29465 ( .A(n35023), .B(n27152), .C(n35024), .Y(n35008) );
  AOI22X1 U29466 ( .A(reg_A[20]), .B(n27513), .C(n27358), .D(n35025), .Y(
        n35024) );
  NAND3X1 U29467 ( .A(n35026), .B(n35027), .C(n35028), .Y(n35025) );
  NOR2X1 U29468 ( .A(n35029), .B(n35030), .Y(n35028) );
  OAI22X1 U29469 ( .A(n27374), .B(n34787), .C(n25250), .D(n27375), .Y(n35030)
         );
  NAND2X1 U29470 ( .A(n35031), .B(n34161), .Y(n34787) );
  AOI22X1 U29471 ( .A(n30587), .B(n26295), .C(n25232), .D(n26293), .Y(n34161)
         );
  AOI22X1 U29472 ( .A(n26292), .B(n27953), .C(n26294), .D(n25250), .Y(n35031)
         );
  OAI22X1 U29473 ( .A(n27377), .B(n34917), .C(n27379), .D(n35032), .Y(n35029)
         );
  OAI21X1 U29474 ( .A(n35033), .B(n26030), .C(n35034), .Y(n34917) );
  AOI22X1 U29475 ( .A(n25025), .B(n34784), .C(n26032), .D(n34428), .Y(n35034)
         );
  OR2X1 U29476 ( .A(n35035), .B(n35036), .Y(n34428) );
  OAI22X1 U29477 ( .A(reg_A[21]), .B(n25063), .C(reg_A[13]), .D(n26981), .Y(
        n35036) );
  OAI21X1 U29478 ( .A(reg_A[5]), .B(n26982), .C(n34721), .Y(n35035) );
  INVX1 U29479 ( .A(n35037), .Y(n34784) );
  INVX1 U29480 ( .A(n35038), .Y(n35033) );
  AOI22X1 U29481 ( .A(n27386), .B(reg_A[18]), .C(n27387), .D(reg_A[17]), .Y(
        n35027) );
  AOI22X1 U29482 ( .A(n27388), .B(reg_A[19]), .C(n27389), .D(reg_A[21]), .Y(
        n35026) );
  AND2X1 U29483 ( .A(n35039), .B(n35040), .Y(n35023) );
  NOR2X1 U29484 ( .A(n35041), .B(n35042), .Y(n35040) );
  OAI21X1 U29485 ( .A(n27960), .B(n26801), .C(n35043), .Y(n35042) );
  AOI22X1 U29486 ( .A(reg_A[27]), .B(n26878), .C(n25613), .D(reg_A[28]), .Y(
        n35043) );
  OAI21X1 U29487 ( .A(n25062), .B(n26714), .C(n35044), .Y(n35041) );
  AOI22X1 U29488 ( .A(reg_A[22]), .B(n26803), .C(reg_A[24]), .D(n26804), .Y(
        n35044) );
  NOR2X1 U29489 ( .A(n35045), .B(n35046), .Y(n35039) );
  OAI22X1 U29490 ( .A(n25736), .B(n25232), .C(n27954), .D(n31398), .Y(n35046)
         );
  OAI21X1 U29491 ( .A(n25239), .B(n27252), .C(n35047), .Y(n35045) );
  AOI22X1 U29492 ( .A(n25750), .B(reg_A[26]), .C(n25614), .D(reg_A[30]), .Y(
        n35047) );
  INVX1 U29493 ( .A(n35048), .Y(n35006) );
  OAI21X1 U29494 ( .A(n25719), .B(n25230), .C(n35049), .Y(n35048) );
  AOI22X1 U29495 ( .A(n35050), .B(n34910), .C(n35051), .D(n34020), .Y(n35049)
         );
  NOR2X1 U29496 ( .A(n35052), .B(n35053), .Y(n35005) );
  OAI21X1 U29497 ( .A(n26714), .B(n25717), .C(n34897), .Y(n35053) );
  INVX1 U29498 ( .A(n35054), .Y(n34897) );
  OAI21X1 U29499 ( .A(n25032), .B(n34485), .C(n35055), .Y(n35054) );
  NAND3X1 U29500 ( .A(reg_B[21]), .B(n26504), .C(n34904), .Y(n35055) );
  NAND2X1 U29501 ( .A(reg_A[16]), .B(reg_B[28]), .Y(n34485) );
  MUX2X1 U29502 ( .B(n35056), .A(n35057), .S(reg_B[31]), .Y(n35052) );
  NAND2X1 U29503 ( .A(n26267), .B(n35058), .Y(n35057) );
  NAND2X1 U29504 ( .A(n34986), .B(n27155), .Y(n35056) );
  OAI22X1 U29505 ( .A(reg_B[30]), .B(n34734), .C(n25220), .D(n34589), .Y(
        n34986) );
  AOI22X1 U29506 ( .A(reg_A[21]), .B(n34189), .C(reg_A[17]), .D(n34190), .Y(
        n34734) );
  NAND3X1 U29507 ( .A(n35059), .B(n35060), .C(n35061), .Y(n35003) );
  NOR2X1 U29508 ( .A(n35062), .B(n35063), .Y(n35061) );
  OAI21X1 U29509 ( .A(n27418), .B(n25220), .C(n35064), .Y(n35063) );
  AOI22X1 U29510 ( .A(reg_A[21]), .B(n27303), .C(reg_A[18]), .D(n27396), .Y(
        n35064) );
  NAND2X1 U29511 ( .A(n35065), .B(n35066), .Y(n27303) );
  INVX1 U29512 ( .A(n27397), .Y(n27418) );
  OAI21X1 U29513 ( .A(n33964), .B(n35002), .C(n35067), .Y(n35062) );
  AOI22X1 U29514 ( .A(n25310), .B(n35068), .C(reg_A[16]), .D(n27316), .Y(
        n35067) );
  OAI22X1 U29515 ( .A(n25207), .B(n27523), .C(n31658), .D(n35069), .Y(n27316)
         );
  NAND3X1 U29516 ( .A(n35070), .B(n35071), .C(n35072), .Y(n35068) );
  NOR2X1 U29517 ( .A(n35073), .B(n35074), .Y(n35072) );
  OAI22X1 U29518 ( .A(n27954), .B(n25219), .C(n25239), .D(n25467), .Y(n35074)
         );
  OAI21X1 U29519 ( .A(n29286), .B(n25223), .C(n35075), .Y(n35073) );
  AOI22X1 U29520 ( .A(n25075), .B(reg_A[25]), .C(n25123), .D(reg_A[26]), .Y(
        n35075) );
  AOI21X1 U29521 ( .A(reg_A[23]), .B(n25252), .C(n35076), .Y(n35071) );
  OAI22X1 U29522 ( .A(n25041), .B(n27962), .C(n25042), .D(n25230), .Y(n35076)
         );
  AOI22X1 U29523 ( .A(n25253), .B(reg_A[27]), .C(n25628), .D(reg_A[28]), .Y(
        n35070) );
  OAI21X1 U29524 ( .A(n34779), .B(n33966), .C(n35077), .Y(n35002) );
  AOI22X1 U29525 ( .A(n32934), .B(n34467), .C(reg_B[30]), .D(n35078), .Y(
        n35077) );
  OR2X1 U29526 ( .A(n35079), .B(n35080), .Y(n34467) );
  OAI22X1 U29527 ( .A(reg_A[21]), .B(n33807), .C(reg_A[13]), .D(n34465), .Y(
        n35080) );
  OAI21X1 U29528 ( .A(reg_A[5]), .B(n34751), .C(n34752), .Y(n35079) );
  AOI21X1 U29529 ( .A(n34975), .B(n35081), .C(n35082), .Y(n35060) );
  OAI21X1 U29530 ( .A(n35083), .B(n25342), .C(n35084), .Y(n35082) );
  OAI21X1 U29531 ( .A(n35085), .B(n35086), .C(n25840), .Y(n35084) );
  NAND3X1 U29532 ( .A(n35087), .B(n35088), .C(n35089), .Y(n35086) );
  NOR2X1 U29533 ( .A(n35090), .B(n35091), .Y(n35089) );
  OAI21X1 U29534 ( .A(n27967), .B(n25219), .C(n35092), .Y(n35091) );
  AOI22X1 U29535 ( .A(n25124), .B(reg_A[13]), .C(n25222), .D(reg_A[10]), .Y(
        n35092) );
  OAI21X1 U29536 ( .A(n25255), .B(n25223), .C(n35093), .Y(n35090) );
  AOI22X1 U29537 ( .A(reg_A[17]), .B(n25073), .C(n25123), .D(reg_A[16]), .Y(
        n35093) );
  AOI21X1 U29538 ( .A(n25635), .B(reg_A[9]), .C(n35094), .Y(n35088) );
  OAI22X1 U29539 ( .A(n26677), .B(n25482), .C(n25132), .D(n25475), .Y(n35094)
         );
  AOI22X1 U29540 ( .A(n25325), .B(reg_A[8]), .C(n25125), .D(reg_A[21]), .Y(
        n35087) );
  NAND3X1 U29541 ( .A(n35095), .B(n35096), .C(n35097), .Y(n35085) );
  NOR2X1 U29542 ( .A(n35098), .B(n35099), .Y(n35097) );
  OAI21X1 U29543 ( .A(n26742), .B(n26719), .C(n35100), .Y(n35099) );
  AOI22X1 U29544 ( .A(n25241), .B(reg_A[3]), .C(n25339), .D(reg_A[1]), .Y(
        n35100) );
  OAI21X1 U29545 ( .A(n25128), .B(n25243), .C(n35101), .Y(n35098) );
  AOI22X1 U29546 ( .A(n25246), .B(reg_A[4]), .C(n25247), .D(reg_A[5]), .Y(
        n35101) );
  AOI21X1 U29547 ( .A(reg_A[19]), .B(n25252), .C(n35102), .Y(n35096) );
  OAI22X1 U29548 ( .A(n25041), .B(n25224), .C(n25042), .D(n30587), .Y(n35102)
         );
  AOI22X1 U29549 ( .A(reg_A[15]), .B(n25253), .C(reg_A[14]), .D(n25628), .Y(
        n35095) );
  AOI22X1 U29550 ( .A(n35103), .B(n35015), .C(n34885), .D(n34881), .Y(n35083)
         );
  MUX2X1 U29551 ( .B(n35104), .A(n35105), .S(reg_B[23]), .Y(n34885) );
  MUX2X1 U29552 ( .B(reg_A[20]), .A(reg_A[16]), .S(reg_B[21]), .Y(n35105) );
  MUX2X1 U29553 ( .B(reg_A[21]), .A(reg_A[17]), .S(reg_B[21]), .Y(n35104) );
  MUX2X1 U29554 ( .B(n25220), .A(n25224), .S(reg_B[23]), .Y(n35103) );
  INVX1 U29555 ( .A(n35106), .Y(n35081) );
  AOI21X1 U29556 ( .A(n25188), .B(n35107), .C(n35108), .Y(n35059) );
  OAI22X1 U29557 ( .A(n27953), .B(n27431), .C(n34387), .D(n35109), .Y(n35108)
         );
  NAND2X1 U29558 ( .A(reg_B[31]), .B(n25932), .Y(n34387) );
  OAI21X1 U29559 ( .A(n30587), .B(n35110), .C(n35111), .Y(n35107) );
  AOI22X1 U29560 ( .A(n35112), .B(n34189), .C(n35113), .D(reg_A[16]), .Y(
        n35111) );
  INVX1 U29561 ( .A(n30648), .Y(n35113) );
  NOR2X1 U29562 ( .A(n25264), .B(n25224), .Y(n35112) );
  NAND3X1 U29563 ( .A(n35114), .B(n35115), .C(n35116), .Y(result[20]) );
  NOR2X1 U29564 ( .A(n35117), .B(n35118), .Y(n35116) );
  NAND3X1 U29565 ( .A(n35119), .B(n35120), .C(n35121), .Y(n35118) );
  AOI21X1 U29566 ( .A(n34910), .B(n35122), .C(n35123), .Y(n35121) );
  OAI22X1 U29567 ( .A(n35124), .B(n30547), .C(n31781), .D(n34902), .Y(n35123)
         );
  INVX1 U29568 ( .A(n34798), .Y(n34902) );
  OAI21X1 U29569 ( .A(reg_B[27]), .B(n26996), .C(n27500), .Y(n34798) );
  INVX1 U29570 ( .A(n35125), .Y(n31781) );
  OAI21X1 U29571 ( .A(n35126), .B(n34230), .C(n35127), .Y(n35125) );
  AOI22X1 U29572 ( .A(n34190), .B(n26778), .C(n34180), .D(n26777), .Y(n35127)
         );
  AOI22X1 U29573 ( .A(reg_A[27]), .B(n25293), .C(reg_A[21]), .D(n25282), .Y(
        n35120) );
  AOI22X1 U29574 ( .A(n30617), .B(n35051), .C(n35012), .D(n35050), .Y(n35119)
         );
  OAI21X1 U29575 ( .A(n30587), .B(n35013), .C(n35128), .Y(n35050) );
  AOI22X1 U29576 ( .A(n34985), .B(reg_A[16]), .C(n35015), .D(reg_A[18]), .Y(
        n35128) );
  NOR2X1 U29577 ( .A(n35129), .B(reg_B[22]), .Y(n34985) );
  NAND2X1 U29578 ( .A(n35130), .B(n35131), .Y(n35051) );
  AOI22X1 U29579 ( .A(n32934), .B(n34528), .C(n34000), .D(n34715), .Y(n35131)
         );
  OAI21X1 U29580 ( .A(n33807), .B(n30587), .C(n35132), .Y(n34528) );
  AOI22X1 U29581 ( .A(n33923), .B(reg_A[4]), .C(reg_A[12]), .D(n33919), .Y(
        n35132) );
  AOI22X1 U29582 ( .A(n33809), .B(n34928), .C(n34015), .D(n35133), .Y(n35130)
         );
  NAND3X1 U29583 ( .A(n35134), .B(n35135), .C(n35136), .Y(n35117) );
  NOR2X1 U29584 ( .A(n35137), .B(n35138), .Y(n35136) );
  OAI22X1 U29585 ( .A(n25295), .B(n27961), .C(n25297), .D(n27960), .Y(n35138)
         );
  OAI22X1 U29586 ( .A(n27511), .B(n27962), .C(n27512), .D(n25244), .Y(n35137)
         );
  AOI22X1 U29587 ( .A(reg_A[19]), .B(n27513), .C(reg_A[30]), .D(n25299), .Y(
        n35135) );
  AOI22X1 U29588 ( .A(reg_A[31]), .B(n25300), .C(reg_A[29]), .D(n25301), .Y(
        n35134) );
  NOR2X1 U29589 ( .A(n35139), .B(n35140), .Y(n35115) );
  NAND2X1 U29590 ( .A(n35141), .B(n35142), .Y(n35140) );
  AOI22X1 U29591 ( .A(reg_A[17]), .B(n35143), .C(reg_A[20]), .D(n35144), .Y(
        n35142) );
  OAI21X1 U29592 ( .A(n25032), .B(n35145), .C(n27423), .Y(n35144) );
  INVX1 U29593 ( .A(n31520), .Y(n27423) );
  OAI21X1 U29594 ( .A(n34822), .B(n35146), .C(n27419), .Y(n35143) );
  INVX1 U29595 ( .A(n27396), .Y(n27419) );
  NAND2X1 U29596 ( .A(reg_B[23]), .B(n25372), .Y(n35146) );
  AOI22X1 U29597 ( .A(n35147), .B(n35148), .C(n34975), .D(n35149), .Y(n35141)
         );
  NOR2X1 U29598 ( .A(n25523), .B(reg_B[21]), .Y(n34975) );
  INVX1 U29599 ( .A(n35078), .Y(n35148) );
  NAND3X1 U29600 ( .A(n35150), .B(n35151), .C(n35152), .Y(n35139) );
  AOI22X1 U29601 ( .A(n35153), .B(n35154), .C(n35155), .D(reg_B[31]), .Y(
        n35152) );
  NOR2X1 U29602 ( .A(n27354), .B(n35156), .Y(n35155) );
  INVX1 U29603 ( .A(n27155), .Y(n27354) );
  NAND2X1 U29604 ( .A(n25032), .B(n25023), .Y(n27155) );
  MUX2X1 U29605 ( .B(n30587), .A(n25220), .S(reg_B[23]), .Y(n35154) );
  NOR2X1 U29606 ( .A(n25031), .B(n35013), .Y(n35153) );
  OAI21X1 U29607 ( .A(n35157), .B(n35158), .C(n25840), .Y(n35151) );
  NAND3X1 U29608 ( .A(n35159), .B(n35160), .C(n35161), .Y(n35158) );
  NOR2X1 U29609 ( .A(n35162), .B(n35163), .Y(n35161) );
  OAI22X1 U29610 ( .A(n30587), .B(n25228), .C(n25132), .D(n25229), .Y(n35163)
         );
  OAI21X1 U29611 ( .A(n26701), .B(n25231), .C(n35164), .Y(n35162) );
  AOI22X1 U29612 ( .A(n25234), .B(reg_A[6]), .C(n25235), .D(reg_A[5]), .Y(
        n35164) );
  AOI21X1 U29613 ( .A(n25124), .B(reg_A[12]), .C(n35165), .Y(n35160) );
  OAI22X1 U29614 ( .A(n27967), .B(n25223), .C(n29279), .D(n26703), .Y(n35165)
         );
  AOI22X1 U29615 ( .A(n25222), .B(reg_A[9]), .C(n25637), .D(reg_A[10]), .Y(
        n35159) );
  NAND3X1 U29616 ( .A(n35166), .B(n35167), .C(n35168), .Y(n35157) );
  NOR2X1 U29617 ( .A(n35169), .B(n35170), .Y(n35168) );
  OAI21X1 U29618 ( .A(n25042), .B(n25220), .C(n35171), .Y(n35170) );
  AOI22X1 U29619 ( .A(n25241), .B(reg_A[2]), .C(n25339), .D(reg_A[0]), .Y(
        n35171) );
  OAI21X1 U29620 ( .A(n25177), .B(n25243), .C(n35172), .Y(n35169) );
  AOI22X1 U29621 ( .A(n25246), .B(reg_A[3]), .C(n25247), .D(reg_A[4]), .Y(
        n35172) );
  AOI21X1 U29622 ( .A(reg_A[14]), .B(n25253), .C(n35173), .Y(n35167) );
  OAI22X1 U29623 ( .A(n25040), .B(n25224), .C(n25254), .D(n27953), .Y(n35173)
         );
  AOI22X1 U29624 ( .A(reg_A[13]), .B(n25628), .C(n25070), .D(reg_A[16]), .Y(
        n35166) );
  OAI21X1 U29625 ( .A(n35174), .B(n35175), .C(n27358), .Y(n35150) );
  OAI22X1 U29626 ( .A(n30587), .B(n27442), .C(n27443), .D(n35176), .Y(n35175)
         );
  OAI21X1 U29627 ( .A(n35177), .B(n25403), .C(n35178), .Y(n35174) );
  INVX1 U29628 ( .A(n35179), .Y(n35178) );
  OAI22X1 U29629 ( .A(n27448), .B(n25250), .C(n34357), .D(n27449), .Y(n35179)
         );
  NAND2X1 U29630 ( .A(n35180), .B(n35181), .Y(n34357) );
  AOI22X1 U29631 ( .A(n26601), .B(n25224), .C(n26602), .D(n27953), .Y(n35181)
         );
  AOI22X1 U29632 ( .A(n27012), .B(n30587), .C(n26597), .D(n25220), .Y(n35180)
         );
  AOI21X1 U29633 ( .A(n35182), .B(n26863), .C(n35183), .Y(n35177) );
  OAI22X1 U29634 ( .A(n27454), .B(n35038), .C(n27455), .D(n35184), .Y(n35183)
         );
  INVX1 U29635 ( .A(n35032), .Y(n35182) );
  OAI21X1 U29636 ( .A(n35185), .B(n26030), .C(n35186), .Y(n35032) );
  AOI22X1 U29637 ( .A(n25025), .B(n34921), .C(n26032), .D(n34567), .Y(n35186)
         );
  OR2X1 U29638 ( .A(n35187), .B(n35188), .Y(n34567) );
  OAI22X1 U29639 ( .A(reg_A[20]), .B(n25063), .C(reg_A[12]), .D(n26981), .Y(
        n35188) );
  OAI21X1 U29640 ( .A(reg_A[4]), .B(n26982), .C(n34721), .Y(n35187) );
  NOR2X1 U29641 ( .A(n35189), .B(n35190), .Y(n35114) );
  OAI21X1 U29642 ( .A(n25360), .B(n26714), .C(n35191), .Y(n35190) );
  AOI22X1 U29643 ( .A(n35192), .B(n30616), .C(reg_A[22]), .D(n25364), .Y(
        n35191) );
  INVX1 U29644 ( .A(n33964), .Y(n30616) );
  INVX1 U29645 ( .A(n35109), .Y(n35192) );
  OAI21X1 U29646 ( .A(n35193), .B(n34176), .C(n35194), .Y(n35109) );
  AOI22X1 U29647 ( .A(n32934), .B(n34562), .C(n33809), .D(n34997), .Y(n35194)
         );
  OR2X1 U29648 ( .A(n35195), .B(n35196), .Y(n34562) );
  OAI22X1 U29649 ( .A(reg_A[20]), .B(n33807), .C(reg_A[12]), .D(n34465), .Y(
        n35196) );
  OAI21X1 U29650 ( .A(reg_A[4]), .B(n34751), .C(n34752), .Y(n35195) );
  INVX1 U29651 ( .A(n35197), .Y(n35193) );
  OR2X1 U29652 ( .A(n35198), .B(n35199), .Y(n35189) );
  OAI21X1 U29653 ( .A(n27943), .B(n35200), .C(n35201), .Y(n35199) );
  OAI21X1 U29654 ( .A(n27397), .B(n35202), .C(reg_A[18]), .Y(n35201) );
  OAI21X1 U29655 ( .A(n34230), .B(n35203), .C(n35204), .Y(n35202) );
  NAND3X1 U29656 ( .A(n25372), .B(n35205), .C(n35206), .Y(n35204) );
  NAND2X1 U29657 ( .A(n25188), .B(n25258), .Y(n35203) );
  OAI21X1 U29658 ( .A(n35207), .B(n35208), .C(n35209), .Y(n35198) );
  OAI21X1 U29659 ( .A(n35210), .B(n35211), .C(reg_A[16]), .Y(n35209) );
  OAI21X1 U29660 ( .A(n25031), .B(n35129), .C(n27431), .Y(n35211) );
  NOR2X1 U29661 ( .A(n34189), .B(n25032), .Y(n35210) );
  INVX1 U29662 ( .A(n35058), .Y(n35207) );
  OAI22X1 U29663 ( .A(reg_B[30]), .B(n34835), .C(n25224), .D(n34589), .Y(
        n35058) );
  INVX1 U29664 ( .A(n35212), .Y(n34589) );
  AOI21X1 U29665 ( .A(reg_A[16]), .B(n34190), .C(n34844), .Y(n34835) );
  INVX1 U29666 ( .A(n34989), .Y(n34844) );
  NAND2X1 U29667 ( .A(n34189), .B(reg_A[20]), .Y(n34989) );
  NAND2X1 U29668 ( .A(n35213), .B(n35214), .Y(result[1]) );
  AOI21X1 U29669 ( .A(reg_A[0]), .B(n35215), .C(n35216), .Y(n35214) );
  OAI21X1 U29670 ( .A(n35217), .B(n25177), .C(n32931), .Y(n35216) );
  NAND3X1 U29671 ( .A(n25372), .B(n35218), .C(reg_A[0]), .Y(n32931) );
  OAI21X1 U29672 ( .A(n31796), .B(n25415), .C(n35219), .Y(n35218) );
  AOI21X1 U29673 ( .A(n25044), .B(n26775), .C(n32997), .Y(n35219) );
  NOR2X1 U29674 ( .A(n35220), .B(n35221), .Y(n35217) );
  OAI21X1 U29675 ( .A(n34088), .B(n25517), .C(n35222), .Y(n35221) );
  OAI21X1 U29676 ( .A(n29566), .B(n31658), .C(n31788), .Y(n35220) );
  NAND2X1 U29677 ( .A(n32985), .B(n25932), .Y(n31788) );
  INVX1 U29678 ( .A(n25284), .Y(n29566) );
  NAND3X1 U29679 ( .A(n35223), .B(n35224), .C(n35225), .Y(n35215) );
  NOR2X1 U29680 ( .A(n35226), .B(n35227), .Y(n35225) );
  OAI22X1 U29681 ( .A(n25156), .B(n27438), .C(n27986), .D(n25342), .Y(n35227)
         );
  OAI21X1 U29682 ( .A(n25125), .B(n25835), .C(n29366), .Y(n35226) );
  AOI22X1 U29683 ( .A(n25170), .B(n32999), .C(n25699), .D(n32984), .Y(n35224)
         );
  INVX1 U29684 ( .A(n35228), .Y(n35223) );
  OAI21X1 U29685 ( .A(n25032), .B(n25116), .C(n35229), .Y(n35228) );
  AOI22X1 U29686 ( .A(n25382), .B(n35230), .C(n25203), .D(n35231), .Y(n35213)
         );
  NAND3X1 U29687 ( .A(n35232), .B(n35233), .C(n35234), .Y(n35231) );
  NOR2X1 U29688 ( .A(n35235), .B(n35236), .Y(n35234) );
  OAI22X1 U29689 ( .A(n26895), .B(n29265), .C(n26893), .D(n26677), .Y(n35236)
         );
  INVX1 U29690 ( .A(n34599), .Y(n26893) );
  OAI21X1 U29691 ( .A(n26894), .B(n25132), .C(n35237), .Y(n35235) );
  OAI21X1 U29692 ( .A(n35238), .B(n35239), .C(n25604), .Y(n35237) );
  NAND2X1 U29693 ( .A(n35240), .B(n35241), .Y(n35239) );
  AOI22X1 U29694 ( .A(n25607), .B(reg_A[11]), .C(n25608), .D(reg_A[15]), .Y(
        n35241) );
  AOI22X1 U29695 ( .A(n25609), .B(reg_A[13]), .C(n25610), .D(reg_A[14]), .Y(
        n35240) );
  NAND2X1 U29696 ( .A(n35242), .B(n35243), .Y(n35238) );
  AOI22X1 U29697 ( .A(n25613), .B(reg_A[8]), .C(n25614), .D(reg_A[10]), .Y(
        n35243) );
  AOI22X1 U29698 ( .A(n25615), .B(reg_A[9]), .C(n25616), .D(reg_A[12]), .Y(
        n35242) );
  AOI21X1 U29699 ( .A(reg_A[3]), .B(n29349), .C(n35244), .Y(n35233) );
  OAI21X1 U29700 ( .A(n35245), .B(n30569), .C(n35246), .Y(n35244) );
  OAI21X1 U29701 ( .A(n35247), .B(n35248), .C(n25044), .Y(n35246) );
  NAND2X1 U29702 ( .A(n35249), .B(n35250), .Y(n35248) );
  NOR2X1 U29703 ( .A(n35251), .B(n35252), .Y(n35250) );
  OAI21X1 U29704 ( .A(n25146), .B(n25467), .C(n35253), .Y(n35252) );
  AOI22X1 U29705 ( .A(n25628), .B(reg_A[8]), .C(n25629), .D(reg_A[10]), .Y(
        n35253) );
  OAI21X1 U29706 ( .A(n29286), .B(n25498), .C(n35254), .Y(n35251) );
  AOI22X1 U29707 ( .A(n25631), .B(reg_A[31]), .C(n25324), .D(reg_A[29]), .Y(
        n35254) );
  NOR2X1 U29708 ( .A(n35255), .B(n35256), .Y(n35249) );
  OAI21X1 U29709 ( .A(n25208), .B(n25229), .C(n35257), .Y(n35256) );
  AOI22X1 U29710 ( .A(n25235), .B(reg_A[16]), .C(n25635), .D(reg_A[13]), .Y(
        n35257) );
  OAI21X1 U29711 ( .A(n29279), .B(n25475), .C(n35258), .Y(n35255) );
  AOI22X1 U29712 ( .A(n25222), .B(reg_A[12]), .C(n25637), .D(reg_A[11]), .Y(
        n35258) );
  NAND2X1 U29713 ( .A(n35259), .B(n35260), .Y(n35247) );
  NOR2X1 U29714 ( .A(n35261), .B(n35262), .Y(n35260) );
  OAI21X1 U29715 ( .A(n27962), .B(n25491), .C(n35263), .Y(n35262) );
  AOI22X1 U29716 ( .A(reg_A[19]), .B(n25241), .C(reg_A[23]), .D(n25242), .Y(
        n35263) );
  OAI21X1 U29717 ( .A(n25038), .B(n30587), .C(n35264), .Y(n35261) );
  AOI22X1 U29718 ( .A(reg_A[18]), .B(n25246), .C(reg_A[17]), .D(n25247), .Y(
        n35264) );
  NOR2X1 U29719 ( .A(n35265), .B(n35266), .Y(n35259) );
  OAI21X1 U29720 ( .A(n32918), .B(n25316), .C(n35267), .Y(n35266) );
  AOI22X1 U29721 ( .A(n25647), .B(reg_A[25]), .C(n25648), .D(reg_A[28]), .Y(
        n35267) );
  OAI21X1 U29722 ( .A(n27961), .B(n25322), .C(n35268), .Y(n35265) );
  AOI22X1 U29723 ( .A(reg_A[21]), .B(n25339), .C(reg_A[22]), .D(n25257), .Y(
        n35268) );
  INVX1 U29724 ( .A(n29346), .Y(n35245) );
  AOI22X1 U29725 ( .A(reg_A[1]), .B(n27639), .C(reg_A[2]), .D(n25617), .Y(
        n35232) );
  NAND3X1 U29726 ( .A(n35269), .B(n35270), .C(n35271), .Y(n35230) );
  NOR2X1 U29727 ( .A(n35272), .B(n35273), .Y(n35271) );
  OAI21X1 U29728 ( .A(n25092), .B(n35274), .C(n35275), .Y(n35273) );
  OAI21X1 U29729 ( .A(n35276), .B(n35277), .C(n25044), .Y(n35275) );
  NAND2X1 U29730 ( .A(n35278), .B(n35279), .Y(n35277) );
  AOI22X1 U29731 ( .A(reg_B[27]), .B(n35280), .C(n26772), .D(n25102), .Y(
        n35279) );
  AOI22X1 U29732 ( .A(reg_A[2]), .B(n32984), .C(n32985), .D(reg_A[1]), .Y(
        n35278) );
  INVX1 U29733 ( .A(n33911), .Y(n32985) );
  NAND2X1 U29734 ( .A(n35281), .B(n35282), .Y(n35276) );
  AOI22X1 U29735 ( .A(n35283), .B(n25258), .C(n29317), .D(n26761), .Y(n35282)
         );
  INVX1 U29736 ( .A(n27944), .Y(n29317) );
  NAND2X1 U29737 ( .A(n25110), .B(reg_A[4]), .Y(n27944) );
  NOR2X1 U29738 ( .A(n25130), .B(n26775), .Y(n35283) );
  AOI22X1 U29739 ( .A(n25101), .B(n30570), .C(n30644), .D(n25111), .Y(n35281)
         );
  NAND2X1 U29740 ( .A(n35284), .B(n35285), .Y(n25111) );
  AOI22X1 U29741 ( .A(n25156), .B(reg_A[9]), .C(n25142), .D(reg_A[10]), .Y(
        n35285) );
  AOI22X1 U29742 ( .A(reg_A[11]), .B(n25258), .C(reg_A[12]), .D(n26761), .Y(
        n35284) );
  NAND2X1 U29743 ( .A(n35286), .B(n35287), .Y(n30570) );
  AOI22X1 U29744 ( .A(n25156), .B(reg_A[5]), .C(n25142), .D(reg_A[6]), .Y(
        n35287) );
  AOI22X1 U29745 ( .A(n25258), .B(reg_A[7]), .C(n26761), .D(reg_A[8]), .Y(
        n35286) );
  INVX1 U29746 ( .A(n35288), .Y(n25092) );
  OAI21X1 U29747 ( .A(n30630), .B(n32976), .C(n35289), .Y(n35272) );
  AOI22X1 U29748 ( .A(n29245), .B(n25090), .C(n32997), .D(n30633), .Y(n35289)
         );
  OAI21X1 U29749 ( .A(n29265), .B(n31786), .C(n35290), .Y(n30633) );
  AOI22X1 U29750 ( .A(n28009), .B(reg_A[6]), .C(n27985), .D(reg_A[7]), .Y(
        n35290) );
  NAND2X1 U29751 ( .A(n35291), .B(n35292), .Y(n25090) );
  AOI22X1 U29752 ( .A(reg_A[11]), .B(n26733), .C(reg_A[10]), .D(n25172), .Y(
        n35292) );
  AOI22X1 U29753 ( .A(reg_A[12]), .B(n26734), .C(n25116), .D(reg_A[9]), .Y(
        n35291) );
  AND2X1 U29754 ( .A(n35293), .B(n35294), .Y(n30630) );
  AOI22X1 U29755 ( .A(n26733), .B(reg_A[7]), .C(reg_A[6]), .D(n25172), .Y(
        n35294) );
  AOI22X1 U29756 ( .A(n26734), .B(reg_A[8]), .C(n25116), .D(reg_A[5]), .Y(
        n35293) );
  AOI22X1 U29757 ( .A(reg_A[3]), .B(n32998), .C(reg_A[2]), .D(n32999), .Y(
        n35270) );
  INVX1 U29758 ( .A(n32947), .Y(n32999) );
  INVX1 U29759 ( .A(n35295), .Y(n32998) );
  AOI22X1 U29760 ( .A(reg_A[4]), .B(n33000), .C(reg_A[1]), .D(n28040), .Y(
        n35269) );
  OR2X1 U29761 ( .A(n35296), .B(n35297), .Y(result[19]) );
  NAND3X1 U29762 ( .A(n35298), .B(n35299), .C(n35300), .Y(n35297) );
  NOR2X1 U29763 ( .A(n35301), .B(n35302), .Y(n35300) );
  OAI21X1 U29764 ( .A(n32946), .B(n25220), .C(n35303), .Y(n35302) );
  AOI22X1 U29765 ( .A(reg_A[26]), .B(n25293), .C(reg_A[20]), .D(n25282), .Y(
        n35303) );
  OAI21X1 U29766 ( .A(n25295), .B(n27960), .C(n35304), .Y(n35301) );
  AOI22X1 U29767 ( .A(reg_A[27]), .B(n25302), .C(reg_A[24]), .D(n29030), .Y(
        n35304) );
  AOI21X1 U29768 ( .A(n26045), .B(n35305), .C(n35306), .Y(n35299) );
  OAI21X1 U29769 ( .A(n35307), .B(n31658), .C(n35308), .Y(n35306) );
  OAI21X1 U29770 ( .A(n35309), .B(n35310), .C(n25372), .Y(n35308) );
  NAND3X1 U29771 ( .A(n35311), .B(n35312), .C(n35313), .Y(n35310) );
  MUX2X1 U29772 ( .B(n35314), .A(n35315), .S(reg_B[23]), .Y(n35313) );
  NOR2X1 U29773 ( .A(n35316), .B(n26999), .Y(n35314) );
  MUX2X1 U29774 ( .B(n35317), .A(n35318), .S(reg_B[30]), .Y(n35311) );
  OAI21X1 U29775 ( .A(n32935), .B(n35200), .C(n35319), .Y(n35318) );
  OAI21X1 U29776 ( .A(n35320), .B(n35321), .C(n34519), .Y(n35319) );
  NOR2X1 U29777 ( .A(reg_B[27]), .B(n35322), .Y(n35320) );
  OAI22X1 U29778 ( .A(n31806), .B(n35197), .C(n32935), .D(n35078), .Y(n35317)
         );
  OAI21X1 U29779 ( .A(reg_B[29]), .B(n34780), .C(n35323), .Y(n35078) );
  AOI21X1 U29780 ( .A(n35324), .B(n33887), .C(n35325), .Y(n35323) );
  INVX1 U29781 ( .A(n35326), .Y(n33887) );
  NOR2X1 U29782 ( .A(n35327), .B(n35328), .Y(n34780) );
  OAI22X1 U29783 ( .A(reg_A[19]), .B(n33807), .C(reg_A[11]), .D(n34465), .Y(
        n35328) );
  OAI21X1 U29784 ( .A(reg_A[3]), .B(n34751), .C(n34752), .Y(n35327) );
  OAI21X1 U29785 ( .A(n25264), .B(n35176), .C(n35329), .Y(n35309) );
  AOI22X1 U29786 ( .A(n35330), .B(n25604), .C(reg_A[18]), .D(n35331), .Y(
        n35329) );
  NOR2X1 U29787 ( .A(reg_B[31]), .B(n35156), .Y(n35330) );
  NOR2X1 U29788 ( .A(n35332), .B(n35333), .Y(n35307) );
  OAI21X1 U29789 ( .A(n26701), .B(n25438), .C(n35334), .Y(n35333) );
  INVX1 U29790 ( .A(n35305), .Y(n35334) );
  OAI21X1 U29791 ( .A(n27564), .B(n25250), .C(n35335), .Y(n35332) );
  OAI21X1 U29792 ( .A(n35336), .B(n35337), .C(n25044), .Y(n35335) );
  OAI22X1 U29793 ( .A(n27454), .B(n35338), .C(n26599), .D(n35038), .Y(n35337)
         );
  OAI21X1 U29794 ( .A(reg_B[2]), .B(n34783), .C(n35339), .Y(n35038) );
  AOI21X1 U29795 ( .A(n27570), .B(n35340), .C(n35341), .Y(n35339) );
  NOR2X1 U29796 ( .A(n35342), .B(n35343), .Y(n34783) );
  OAI22X1 U29797 ( .A(reg_A[19]), .B(n25063), .C(reg_A[11]), .D(n26981), .Y(
        n35343) );
  OAI21X1 U29798 ( .A(reg_A[3]), .B(n26982), .C(n34721), .Y(n35342) );
  OAI21X1 U29799 ( .A(n27575), .B(n35184), .C(n35344), .Y(n35336) );
  AOI22X1 U29800 ( .A(n35345), .B(n27577), .C(n27579), .D(reg_A[0]), .Y(n35344) );
  NOR2X1 U29801 ( .A(n35346), .B(n33393), .Y(n27564) );
  INVX1 U29802 ( .A(n35347), .Y(n33393) );
  OAI21X1 U29803 ( .A(n26010), .B(n35348), .C(n25604), .Y(n35347) );
  OAI21X1 U29804 ( .A(n25204), .B(n25220), .C(n35349), .Y(n35305) );
  AOI22X1 U29805 ( .A(reg_A[18]), .B(n25441), .C(reg_A[17]), .D(n27243), .Y(
        n35349) );
  AOI21X1 U29806 ( .A(n34910), .B(n35350), .C(n35351), .Y(n35298) );
  OAI22X1 U29807 ( .A(n35316), .B(n34903), .C(n35124), .D(n31828), .Y(n35351)
         );
  AND2X1 U29808 ( .A(n35352), .B(n35353), .Y(n35124) );
  AOI22X1 U29809 ( .A(n32934), .B(n34620), .C(n34000), .D(n34830), .Y(n35353)
         );
  OAI21X1 U29810 ( .A(n33807), .B(n25220), .C(n35354), .Y(n34620) );
  AOI22X1 U29811 ( .A(n33923), .B(reg_A[3]), .C(reg_A[11]), .D(n33919), .Y(
        n35354) );
  AOI22X1 U29812 ( .A(n33809), .B(n35019), .C(n34015), .D(n35355), .Y(n35352)
         );
  INVX1 U29813 ( .A(n35122), .Y(n35316) );
  OAI22X1 U29814 ( .A(n25220), .B(n35013), .C(n27953), .D(n34984), .Y(n35122)
         );
  INVX1 U29815 ( .A(n35356), .Y(n34910) );
  NAND3X1 U29816 ( .A(n35357), .B(n35358), .C(n35359), .Y(n35296) );
  NOR2X1 U29817 ( .A(n35360), .B(n35361), .Y(n35359) );
  OAI21X1 U29818 ( .A(n31590), .B(n25244), .C(n35362), .Y(n35361) );
  AOI22X1 U29819 ( .A(reg_A[29]), .B(n25299), .C(reg_A[30]), .D(n25300), .Y(
        n35362) );
  OAI21X1 U29820 ( .A(n25360), .B(n25230), .C(n35363), .Y(n35360) );
  AOI22X1 U29821 ( .A(reg_A[31]), .B(n25363), .C(reg_A[21]), .D(n25364), .Y(
        n35363) );
  NOR2X1 U29822 ( .A(n35364), .B(n35365), .Y(n35358) );
  OAI22X1 U29823 ( .A(n25250), .B(n27587), .C(n35156), .D(n35208), .Y(n35365)
         );
  AOI22X1 U29824 ( .A(reg_A[17]), .B(n35212), .C(reg_A[19]), .D(n34011), .Y(
        n35156) );
  OAI21X1 U29825 ( .A(n26147), .B(n35366), .C(n35367), .Y(n35364) );
  OAI21X1 U29826 ( .A(n35368), .B(n35369), .C(n25840), .Y(n35367) );
  NAND3X1 U29827 ( .A(n35370), .B(n35371), .C(n35372), .Y(n35369) );
  NOR2X1 U29828 ( .A(n35373), .B(n35374), .Y(n35372) );
  OAI22X1 U29829 ( .A(n25220), .B(n25228), .C(n26677), .D(n25229), .Y(n35374)
         );
  OAI21X1 U29830 ( .A(n25132), .B(n25231), .C(n35375), .Y(n35373) );
  AOI22X1 U29831 ( .A(n25234), .B(reg_A[5]), .C(n25235), .D(reg_A[4]), .Y(
        n35375) );
  AOI21X1 U29832 ( .A(n25124), .B(reg_A[11]), .C(n35376), .Y(n35371) );
  OAI22X1 U29833 ( .A(n25147), .B(n25223), .C(n26703), .D(n25208), .Y(n35376)
         );
  AOI22X1 U29834 ( .A(n25222), .B(reg_A[8]), .C(n25637), .D(reg_A[9]), .Y(
        n35370) );
  NAND3X1 U29835 ( .A(n35377), .B(n35378), .C(n35379), .Y(n35368) );
  NOR2X1 U29836 ( .A(n35380), .B(n35381), .Y(n35379) );
  OAI22X1 U29837 ( .A(n25042), .B(n25224), .C(n25177), .D(n25331), .Y(n35381)
         );
  OAI21X1 U29838 ( .A(n26742), .B(n25243), .C(n35382), .Y(n35380) );
  AOI22X1 U29839 ( .A(n25246), .B(reg_A[2]), .C(n25247), .D(reg_A[3]), .Y(
        n35382) );
  AOI21X1 U29840 ( .A(reg_A[13]), .B(n25253), .C(n35383), .Y(n35378) );
  OAI22X1 U29841 ( .A(n25040), .B(n27953), .C(n25041), .D(n25250), .Y(n35383)
         );
  AOI22X1 U29842 ( .A(n25628), .B(reg_A[12]), .C(n25070), .D(reg_A[15]), .Y(
        n35377) );
  OR2X1 U29843 ( .A(n33865), .B(n35384), .Y(n35366) );
  AOI21X1 U29844 ( .A(n34020), .B(n35385), .C(n35386), .Y(n35357) );
  OAI21X1 U29845 ( .A(n32909), .B(n26714), .C(n35387), .Y(n35386) );
  OAI21X1 U29846 ( .A(n35388), .B(n35389), .C(n25382), .Y(n35387) );
  OAI21X1 U29847 ( .A(n35390), .B(n35391), .C(n35392), .Y(n35389) );
  NAND3X1 U29848 ( .A(n34825), .B(reg_A[23]), .C(n34884), .Y(n35392) );
  INVX1 U29849 ( .A(n32989), .Y(n35390) );
  OAI21X1 U29850 ( .A(n34403), .B(n34493), .C(n35393), .Y(n32989) );
  AOI22X1 U29851 ( .A(n34189), .B(n35394), .C(n34190), .D(n34808), .Y(n35393)
         );
  MUX2X1 U29852 ( .B(n35395), .A(n35396), .S(reg_B[23]), .Y(n35388) );
  AOI22X1 U29853 ( .A(n34826), .B(reg_A[20]), .C(n35206), .D(reg_A[22]), .Y(
        n35396) );
  OR2X1 U29854 ( .A(n35397), .B(n35398), .Y(result[18]) );
  NAND3X1 U29855 ( .A(n35399), .B(n35400), .C(n35401), .Y(n35398) );
  NOR2X1 U29856 ( .A(n35402), .B(n35403), .Y(n35401) );
  OAI21X1 U29857 ( .A(n35404), .B(n30547), .C(n35405), .Y(n35403) );
  OAI21X1 U29858 ( .A(n35406), .B(n35407), .C(n25203), .Y(n35405) );
  NAND3X1 U29859 ( .A(n35408), .B(n35409), .C(n35410), .Y(n35407) );
  AOI21X1 U29860 ( .A(reg_A[20]), .B(n27637), .C(n35411), .Y(n35410) );
  OAI22X1 U29861 ( .A(n25599), .B(n25232), .C(n25600), .D(n26714), .Y(n35411)
         );
  AOI22X1 U29862 ( .A(reg_A[18]), .B(n27639), .C(reg_A[19]), .D(n25617), .Y(
        n35409) );
  AOI22X1 U29863 ( .A(reg_A[22]), .B(n25650), .C(reg_A[24]), .D(n25651), .Y(
        n35408) );
  NAND3X1 U29864 ( .A(n35412), .B(n35413), .C(n35414), .Y(n35406) );
  AOI21X1 U29865 ( .A(reg_A[29]), .B(n27643), .C(n35415), .Y(n35414) );
  OAI22X1 U29866 ( .A(n27645), .B(n25244), .C(n27646), .D(n32918), .Y(n35415)
         );
  AOI22X1 U29867 ( .A(reg_A[30]), .B(n27647), .C(reg_A[31]), .D(n27648), .Y(
        n35413) );
  AOI22X1 U29868 ( .A(reg_A[25]), .B(n27649), .C(reg_A[26]), .D(n27650), .Y(
        n35412) );
  OAI21X1 U29869 ( .A(n35416), .B(n35417), .C(n35418), .Y(n35402) );
  OAI21X1 U29870 ( .A(n35419), .B(n35420), .C(n25372), .Y(n35418) );
  NAND2X1 U29871 ( .A(n35421), .B(n35312), .Y(n35420) );
  AOI22X1 U29872 ( .A(reg_A[18]), .B(n35422), .C(n34242), .D(reg_B[30]), .Y(
        n35421) );
  OAI21X1 U29873 ( .A(n35423), .B(n25403), .C(n35424), .Y(n35419) );
  AOI21X1 U29874 ( .A(reg_A[17]), .B(n35331), .C(n35315), .Y(n35424) );
  NOR2X1 U29875 ( .A(n35425), .B(n26999), .Y(n35315) );
  OAI22X1 U29876 ( .A(n35426), .B(n35205), .C(n25415), .D(n35110), .Y(n35331)
         );
  NOR2X1 U29877 ( .A(n35427), .B(n35428), .Y(n35423) );
  OAI22X1 U29878 ( .A(n26758), .B(n35200), .C(n25262), .D(n35197), .Y(n35428)
         );
  OAI21X1 U29879 ( .A(reg_B[29]), .B(n34998), .C(n35429), .Y(n35197) );
  AOI21X1 U29880 ( .A(n35324), .B(n33971), .C(n35325), .Y(n35429) );
  NOR2X1 U29881 ( .A(n35430), .B(n35431), .Y(n34998) );
  OAI22X1 U29882 ( .A(reg_A[18]), .B(n33807), .C(reg_A[10]), .D(n34465), .Y(
        n35431) );
  OAI21X1 U29883 ( .A(reg_A[2]), .B(n34751), .C(n34752), .Y(n35430) );
  OAI21X1 U29884 ( .A(n29305), .B(n35432), .C(n35433), .Y(n35427) );
  OAI21X1 U29885 ( .A(n35434), .B(n35321), .C(n26761), .Y(n35433) );
  NOR2X1 U29886 ( .A(reg_B[27]), .B(n35435), .Y(n35434) );
  MUX2X1 U29887 ( .B(n35436), .A(n35437), .S(reg_B[29]), .Y(n35432) );
  OAI21X1 U29888 ( .A(reg_B[27]), .B(n35438), .C(n35439), .Y(n35437) );
  INVX1 U29889 ( .A(n34997), .Y(n35436) );
  OAI21X1 U29890 ( .A(reg_A[0]), .B(n31782), .C(n35440), .Y(n34997) );
  AOI22X1 U29891 ( .A(n33919), .B(n26701), .C(n32933), .D(n25250), .Y(n35440)
         );
  NAND2X1 U29892 ( .A(n35441), .B(n27676), .Y(n35417) );
  AOI22X1 U29893 ( .A(n26597), .B(n35184), .C(n26009), .D(n34921), .Y(n35441)
         );
  OAI21X1 U29894 ( .A(reg_A[0]), .B(n27677), .C(n35442), .Y(n34921) );
  AOI22X1 U29895 ( .A(n26038), .B(n26701), .C(n26664), .D(n25250), .Y(n35442)
         );
  OAI21X1 U29896 ( .A(n35185), .B(n26599), .C(n35443), .Y(n35416) );
  AOI22X1 U29897 ( .A(n27680), .B(n26742), .C(n35444), .D(n27677), .Y(n35443)
         );
  OAI21X1 U29898 ( .A(n35445), .B(n25754), .C(n35446), .Y(n35444) );
  AOI22X1 U29899 ( .A(n26002), .B(n34430), .C(n26008), .D(n35340), .Y(n35446)
         );
  INVX1 U29900 ( .A(n35338), .Y(n35185) );
  OAI21X1 U29901 ( .A(reg_B[2]), .B(n34920), .C(n35447), .Y(n35338) );
  AOI21X1 U29902 ( .A(n27570), .B(n33987), .C(n35341), .Y(n35447) );
  NOR2X1 U29903 ( .A(n35448), .B(n35449), .Y(n34920) );
  OAI22X1 U29904 ( .A(reg_A[18]), .B(n26036), .C(reg_A[10]), .D(n26981), .Y(
        n35449) );
  OAI21X1 U29905 ( .A(reg_A[2]), .B(n26982), .C(n34721), .Y(n35448) );
  AOI22X1 U29906 ( .A(n25509), .B(reg_A[23]), .C(n30617), .D(n35385), .Y(
        n35400) );
  NAND2X1 U29907 ( .A(n35450), .B(n35451), .Y(n35385) );
  AOI22X1 U29908 ( .A(n32934), .B(n34715), .C(n34000), .D(n34928), .Y(n35451)
         );
  OAI21X1 U29909 ( .A(n33807), .B(n25224), .C(n35452), .Y(n34715) );
  AOI22X1 U29910 ( .A(n33923), .B(reg_A[2]), .C(reg_A[10]), .D(n33919), .Y(
        n35452) );
  AOI22X1 U29911 ( .A(n34015), .B(n35453), .C(n33809), .D(n35133), .Y(n35450)
         );
  AOI22X1 U29912 ( .A(reg_A[18]), .B(n27687), .C(n35012), .D(n35350), .Y(
        n35399) );
  OAI22X1 U29913 ( .A(n25224), .B(n35013), .C(reg_B[21]), .D(n35425), .Y(
        n35350) );
  INVX1 U29914 ( .A(n34904), .Y(n35425) );
  NOR2X1 U29915 ( .A(n34881), .B(n25250), .Y(n34904) );
  INVX1 U29916 ( .A(n34903), .Y(n35012) );
  NAND3X1 U29917 ( .A(n35454), .B(n35455), .C(n35456), .Y(n35397) );
  NOR2X1 U29918 ( .A(n35457), .B(n35458), .Y(n35456) );
  OAI21X1 U29919 ( .A(n27698), .B(n25250), .C(n35459), .Y(n35458) );
  OAI21X1 U29920 ( .A(n35460), .B(n35461), .C(n25382), .Y(n35459) );
  OAI22X1 U29921 ( .A(n35462), .B(n35463), .C(n34142), .D(n35391), .Y(n35461)
         );
  AND2X1 U29922 ( .A(n35464), .B(n35465), .Y(n34142) );
  AOI22X1 U29923 ( .A(n34188), .B(n34908), .C(n34180), .D(n34909), .Y(n35465)
         );
  AOI22X1 U29924 ( .A(n34190), .B(n35466), .C(n34189), .D(n35467), .Y(n35464)
         );
  INVX1 U29925 ( .A(n34976), .Y(n35462) );
  OAI21X1 U29926 ( .A(n25230), .B(n35468), .C(n35469), .Y(n34976) );
  NAND3X1 U29927 ( .A(reg_A[23]), .B(n34881), .C(reg_B[23]), .Y(n35469) );
  MUX2X1 U29928 ( .B(n35470), .A(n35395), .S(reg_B[23]), .Y(n35460) );
  AOI22X1 U29929 ( .A(reg_A[21]), .B(n35206), .C(reg_A[19]), .D(n34826), .Y(
        n35395) );
  INVX1 U29930 ( .A(n35471), .Y(n27698) );
  OAI21X1 U29931 ( .A(n35472), .B(n31658), .C(n35473), .Y(n35471) );
  AOI21X1 U29932 ( .A(n25589), .B(n35474), .C(n35475), .Y(n35472) );
  NAND2X1 U29933 ( .A(n33592), .B(n35476), .Y(n35475) );
  OAI21X1 U29934 ( .A(reg_B[3]), .B(n35348), .C(n25604), .Y(n33592) );
  OAI21X1 U29935 ( .A(n35384), .B(n35208), .C(n35477), .Y(n35457) );
  AND2X1 U29936 ( .A(n35478), .B(n35479), .Y(n35477) );
  OAI21X1 U29937 ( .A(n35480), .B(n35481), .C(n25840), .Y(n35479) );
  NAND3X1 U29938 ( .A(n35482), .B(n35483), .C(n35484), .Y(n35481) );
  NOR2X1 U29939 ( .A(n35485), .B(n35486), .Y(n35484) );
  OAI22X1 U29940 ( .A(n30569), .B(n25475), .C(n26701), .D(n25219), .Y(n35486)
         );
  OAI21X1 U29941 ( .A(n25132), .B(n25473), .C(n35487), .Y(n35485) );
  AOI22X1 U29942 ( .A(n25629), .B(reg_A[9]), .C(n25124), .D(reg_A[10]), .Y(
        n35487) );
  AOI22X1 U29943 ( .A(n25235), .B(reg_A[3]), .C(n25635), .D(reg_A[6]), .Y(
        n35483) );
  AOI22X1 U29944 ( .A(n25325), .B(reg_A[5]), .C(n25125), .D(reg_A[18]), .Y(
        n35482) );
  NAND3X1 U29945 ( .A(n35488), .B(n35489), .C(n35490), .Y(n35480) );
  NOR2X1 U29946 ( .A(n35491), .B(n35492), .Y(n35490) );
  OAI22X1 U29947 ( .A(n25206), .B(n26703), .C(n26431), .D(n25208), .Y(n35492)
         );
  OAI21X1 U29948 ( .A(n27967), .B(n25129), .C(n35493), .Y(n35491) );
  AOI22X1 U29949 ( .A(reg_A[16]), .B(n25252), .C(n25253), .D(reg_A[12]), .Y(
        n35493) );
  AOI21X1 U29950 ( .A(n25241), .B(reg_A[0]), .C(n35494), .Y(n35489) );
  OAI22X1 U29951 ( .A(n25128), .B(n25334), .C(n25177), .D(n25336), .Y(n35494)
         );
  AOI22X1 U29952 ( .A(reg_A[17]), .B(n25135), .C(reg_A[15]), .D(n25136), .Y(
        n35488) );
  OAI21X1 U29953 ( .A(n27725), .B(n35495), .C(reg_A[17]), .Y(n35478) );
  INVX1 U29954 ( .A(n31718), .Y(n27725) );
  NAND2X1 U29955 ( .A(n26267), .B(n33865), .Y(n35208) );
  AOI22X1 U29956 ( .A(reg_A[16]), .B(n35212), .C(reg_A[18]), .D(n34011), .Y(
        n35384) );
  NOR2X1 U29957 ( .A(n34012), .B(reg_B[28]), .Y(n34011) );
  NOR2X1 U29958 ( .A(n34230), .B(n34176), .Y(n35212) );
  AOI22X1 U29959 ( .A(n25369), .B(reg_A[8]), .C(n25506), .D(reg_A[20]), .Y(
        n35455) );
  AOI22X1 U29960 ( .A(n25507), .B(reg_A[21]), .C(n25508), .D(reg_A[22]), .Y(
        n35454) );
  INVX1 U29961 ( .A(n29765), .Y(n25507) );
  NAND3X1 U29962 ( .A(n35496), .B(n35497), .C(n35498), .Y(result[17]) );
  NOR2X1 U29963 ( .A(n35499), .B(n35500), .Y(n35498) );
  NAND3X1 U29964 ( .A(n35501), .B(n35502), .C(n35503), .Y(n35500) );
  AOI21X1 U29965 ( .A(n29779), .B(reg_A[23]), .C(n35504), .Y(n35503) );
  OAI22X1 U29966 ( .A(n27826), .B(n35340), .C(n27825), .D(n35184), .Y(n35504)
         );
  OAI21X1 U29967 ( .A(reg_B[2]), .B(n35037), .C(n35505), .Y(n35184) );
  AOI21X1 U29968 ( .A(n27570), .B(n34207), .C(n35341), .Y(n35505) );
  AND2X1 U29969 ( .A(n27828), .B(n26742), .Y(n35341) );
  NOR2X1 U29970 ( .A(n35506), .B(n35507), .Y(n35037) );
  OAI22X1 U29971 ( .A(reg_A[17]), .B(n26036), .C(reg_A[9]), .D(n26981), .Y(
        n35507) );
  OAI21X1 U29972 ( .A(reg_A[1]), .B(n26982), .C(n34721), .Y(n35506) );
  NAND2X1 U29973 ( .A(n26662), .B(n26742), .Y(n34721) );
  OAI21X1 U29974 ( .A(n35508), .B(n35509), .C(n25382), .Y(n35502) );
  OAI22X1 U29975 ( .A(n35510), .B(n35391), .C(n35106), .D(n35463), .Y(n35509)
         );
  MUX2X1 U29976 ( .B(n35511), .A(n35512), .S(reg_B[23]), .Y(n35106) );
  NOR2X1 U29977 ( .A(reg_B[22]), .B(n25230), .Y(n35512) );
  INVX1 U29978 ( .A(n35280), .Y(n35510) );
  NAND2X1 U29979 ( .A(n35513), .B(n35514), .Y(n35280) );
  AOI22X1 U29980 ( .A(n34188), .B(n25109), .C(n34190), .D(n35022), .Y(n35514)
         );
  AOI22X1 U29981 ( .A(n34180), .B(n25104), .C(n34189), .D(n30643), .Y(n35513)
         );
  MUX2X1 U29982 ( .B(n35515), .A(n35470), .S(reg_B[23]), .Y(n35508) );
  AOI22X1 U29983 ( .A(reg_A[20]), .B(n35206), .C(reg_A[18]), .D(n34826), .Y(
        n35470) );
  INVX1 U29984 ( .A(n34822), .Y(n35206) );
  INVX1 U29985 ( .A(n35516), .Y(n35515) );
  OAI21X1 U29986 ( .A(n35495), .B(n35517), .C(reg_A[16]), .Y(n35501) );
  OAI21X1 U29987 ( .A(n34884), .B(n25342), .C(n27767), .Y(n35517) );
  NAND2X1 U29988 ( .A(n27358), .B(n33618), .Y(n27767) );
  OAI21X1 U29989 ( .A(n26004), .B(n26999), .C(n35518), .Y(n33618) );
  INVX1 U29990 ( .A(n35519), .Y(n35518) );
  OAI21X1 U29991 ( .A(n25415), .B(n27012), .C(n35476), .Y(n35519) );
  INVX1 U29992 ( .A(n35468), .Y(n34884) );
  OAI21X1 U29993 ( .A(n35013), .B(n35356), .C(n35520), .Y(n35495) );
  AOI21X1 U29994 ( .A(n35521), .B(n26267), .C(n27770), .Y(n35520) );
  INVX1 U29995 ( .A(n35110), .Y(n35521) );
  NAND2X1 U29996 ( .A(n34405), .B(n34493), .Y(n35110) );
  NAND2X1 U29997 ( .A(reg_B[23]), .B(n26186), .Y(n35356) );
  NAND3X1 U29998 ( .A(n35522), .B(n35523), .C(n35524), .Y(n35499) );
  INVX1 U29999 ( .A(n35525), .Y(n35524) );
  OAI22X1 U30000 ( .A(n34430), .B(n27820), .C(n35526), .D(n27821), .Y(n35525)
         );
  INVX1 U30001 ( .A(n35527), .Y(n34430) );
  OAI21X1 U30002 ( .A(n27687), .B(n35528), .C(reg_A[17]), .Y(n35523) );
  AND2X1 U30003 ( .A(n35529), .B(n35530), .Y(n35522) );
  OAI21X1 U30004 ( .A(n35531), .B(n35532), .C(n25840), .Y(n35530) );
  NAND3X1 U30005 ( .A(n35533), .B(n35534), .C(n35535), .Y(n35532) );
  NOR2X1 U30006 ( .A(n35536), .B(n35537), .Y(n35535) );
  OAI22X1 U30007 ( .A(n25130), .B(n25475), .C(n25132), .D(n25219), .Y(n35537)
         );
  OAI21X1 U30008 ( .A(n26677), .B(n25473), .C(n35538), .Y(n35536) );
  AOI22X1 U30009 ( .A(n25629), .B(reg_A[8]), .C(n25124), .D(reg_A[9]), .Y(
        n35538) );
  AOI22X1 U30010 ( .A(n25235), .B(reg_A[2]), .C(n25635), .D(reg_A[5]), .Y(
        n35534) );
  AOI22X1 U30011 ( .A(n25325), .B(reg_A[4]), .C(n25125), .D(reg_A[17]), .Y(
        n35533) );
  NAND3X1 U30012 ( .A(n35539), .B(n35540), .C(n35541), .Y(n35531) );
  NOR2X1 U30013 ( .A(n35542), .B(n35543), .Y(n35541) );
  OAI22X1 U30014 ( .A(n25040), .B(n29279), .C(n25041), .D(n25208), .Y(n35543)
         );
  OAI21X1 U30015 ( .A(n25042), .B(n25250), .C(n35544), .Y(n35542) );
  AOI22X1 U30016 ( .A(n25246), .B(reg_A[0]), .C(n25247), .D(reg_A[1]), .Y(
        n35544) );
  AOI22X1 U30017 ( .A(n25253), .B(reg_A[11]), .C(n25628), .D(reg_A[10]), .Y(
        n35540) );
  AOI22X1 U30018 ( .A(reg_A[13]), .B(n25073), .C(n25123), .D(reg_A[12]), .Y(
        n35539) );
  OAI21X1 U30019 ( .A(n35545), .B(n35546), .C(n25372), .Y(n35529) );
  OAI21X1 U30020 ( .A(n25156), .B(n35176), .C(n35312), .Y(n35546) );
  AOI22X1 U30021 ( .A(reg_A[16]), .B(n34825), .C(n34230), .D(n34242), .Y(
        n35312) );
  INVX1 U30022 ( .A(n35176), .Y(n34242) );
  INVX1 U30023 ( .A(n35463), .Y(n34825) );
  NAND2X1 U30024 ( .A(reg_A[16]), .B(n25604), .Y(n35176) );
  OAI21X1 U30025 ( .A(n35547), .B(n27953), .C(n35548), .Y(n35545) );
  AOI22X1 U30026 ( .A(n34519), .B(n35549), .C(n34173), .D(n35550), .Y(n35548)
         );
  OAI21X1 U30027 ( .A(reg_B[27]), .B(n35551), .C(n35552), .Y(n35550) );
  INVX1 U30028 ( .A(n35553), .Y(n35552) );
  MUX2X1 U30029 ( .B(n35200), .A(n35439), .S(reg_B[30]), .Y(n35553) );
  OAI21X1 U30030 ( .A(reg_B[29]), .B(n34779), .C(n35554), .Y(n35200) );
  AOI21X1 U30031 ( .A(n35324), .B(n35555), .C(n35325), .Y(n35554) );
  INVX1 U30032 ( .A(n35556), .Y(n35325) );
  NAND3X1 U30033 ( .A(reg_B[27]), .B(n26742), .C(reg_B[29]), .Y(n35556) );
  INVX1 U30034 ( .A(n34217), .Y(n35555) );
  NOR2X1 U30035 ( .A(n33955), .B(reg_B[27]), .Y(n35324) );
  NOR2X1 U30036 ( .A(n35557), .B(n35558), .Y(n34779) );
  OAI22X1 U30037 ( .A(reg_A[17]), .B(n33807), .C(reg_A[9]), .D(n34465), .Y(
        n35558) );
  OAI21X1 U30038 ( .A(reg_A[1]), .B(n34751), .C(n34752), .Y(n35557) );
  NAND2X1 U30039 ( .A(n33922), .B(n26742), .Y(n34752) );
  NOR2X1 U30040 ( .A(n34493), .B(n31782), .Y(n33922) );
  AOI22X1 U30041 ( .A(n34464), .B(n34015), .C(n35326), .D(n34000), .Y(n35551)
         );
  INVX1 U30042 ( .A(n32935), .Y(n34173) );
  OAI21X1 U30043 ( .A(reg_B[27]), .B(n35559), .C(n35439), .Y(n35549) );
  INVX1 U30044 ( .A(n31806), .Y(n34519) );
  INVX1 U30045 ( .A(n35422), .Y(n35547) );
  OAI21X1 U30046 ( .A(n25415), .B(n35145), .C(n34837), .Y(n35422) );
  NOR2X1 U30047 ( .A(n35560), .B(n35561), .Y(n35497) );
  OAI22X1 U30048 ( .A(n25232), .B(n29782), .C(n30587), .D(n29765), .Y(n35561)
         );
  OAI21X1 U30049 ( .A(n25220), .B(n29766), .C(n35562), .Y(n35560) );
  AOI22X1 U30050 ( .A(reg_A[0]), .B(n27778), .C(n25369), .D(reg_A[8]), .Y(
        n35562) );
  INVX1 U30051 ( .A(n25583), .Y(n25369) );
  NAND2X1 U30052 ( .A(n27387), .B(n27358), .Y(n25583) );
  OAI22X1 U30053 ( .A(n27677), .B(n26012), .C(n26030), .D(n31636), .Y(n27778)
         );
  NOR2X1 U30054 ( .A(n35563), .B(n35564), .Y(n35496) );
  OAI21X1 U30055 ( .A(n35404), .B(n31828), .C(n35565), .Y(n35564) );
  OAI21X1 U30056 ( .A(n35566), .B(n35567), .C(n25203), .Y(n35565) );
  NAND3X1 U30057 ( .A(n35568), .B(n35569), .C(n35570), .Y(n35567) );
  AOI22X1 U30058 ( .A(reg_A[20]), .B(n27740), .C(reg_A[19]), .D(n27637), .Y(
        n35570) );
  OAI21X1 U30059 ( .A(n35571), .B(n35572), .C(n25044), .Y(n35569) );
  NAND2X1 U30060 ( .A(n35573), .B(n35574), .Y(n35572) );
  AOI22X1 U30061 ( .A(n25637), .B(reg_A[27]), .C(n25234), .D(reg_A[31]), .Y(
        n35574) );
  AOI22X1 U30062 ( .A(n25635), .B(reg_A[29]), .C(n25325), .D(reg_A[30]), .Y(
        n35573) );
  NAND2X1 U30063 ( .A(n35575), .B(n35576), .Y(n35571) );
  AOI22X1 U30064 ( .A(reg_A[24]), .B(n25628), .C(n25629), .D(reg_A[26]), .Y(
        n35576) );
  AOI22X1 U30065 ( .A(n25124), .B(reg_A[25]), .C(n25222), .D(reg_A[28]), .Y(
        n35575) );
  OAI21X1 U30066 ( .A(n35577), .B(n35578), .C(n25604), .Y(n35568) );
  NAND2X1 U30067 ( .A(n35579), .B(n35580), .Y(n35578) );
  AOI22X1 U30068 ( .A(n25607), .B(reg_A[27]), .C(n25608), .D(reg_A[31]), .Y(
        n35580) );
  AOI22X1 U30069 ( .A(n25609), .B(reg_A[29]), .C(n25610), .D(reg_A[30]), .Y(
        n35579) );
  NAND2X1 U30070 ( .A(n35581), .B(n35582), .Y(n35577) );
  AOI22X1 U30071 ( .A(reg_A[24]), .B(n25613), .C(n25614), .D(reg_A[26]), .Y(
        n35582) );
  AOI22X1 U30072 ( .A(n25615), .B(reg_A[25]), .C(n25616), .D(reg_A[28]), .Y(
        n35581) );
  OR2X1 U30073 ( .A(n35583), .B(n35584), .Y(n35566) );
  OAI22X1 U30074 ( .A(n25600), .B(n25230), .C(n27755), .D(n26714), .Y(n35584)
         );
  OAI21X1 U30075 ( .A(n27756), .B(n25232), .C(n35585), .Y(n35583) );
  AOI22X1 U30076 ( .A(reg_A[17]), .B(n27639), .C(reg_A[18]), .D(n25617), .Y(
        n35585) );
  AND2X1 U30077 ( .A(n35586), .B(n35587), .Y(n35404) );
  AOI22X1 U30078 ( .A(n32934), .B(n34830), .C(n34000), .D(n35019), .Y(n35587)
         );
  OAI21X1 U30079 ( .A(n33807), .B(n27953), .C(n35588), .Y(n34830) );
  AOI22X1 U30080 ( .A(n33923), .B(reg_A[1]), .C(reg_A[9]), .D(n33919), .Y(
        n35588) );
  AOI22X1 U30081 ( .A(n34015), .B(n35589), .C(n33809), .D(n35355), .Y(n35586)
         );
  OAI22X1 U30082 ( .A(n35590), .B(n30547), .C(n25230), .D(n25652), .Y(n35563)
         );
  INVX1 U30083 ( .A(n35591), .Y(n35590) );
  OR2X1 U30084 ( .A(n35592), .B(n35593), .Y(result[16]) );
  NAND3X1 U30085 ( .A(n35594), .B(n35595), .C(n35596), .Y(n35593) );
  NOR2X1 U30086 ( .A(n35597), .B(n35598), .Y(n35596) );
  OAI22X1 U30087 ( .A(n25224), .B(n25717), .C(n25220), .D(n25718), .Y(n35598)
         );
  OAI21X1 U30088 ( .A(n27953), .B(n25719), .C(n35599), .Y(n35597) );
  AOI22X1 U30089 ( .A(n34020), .B(n35600), .C(n25722), .D(reg_A[20]), .Y(
        n35599) );
  INVX1 U30090 ( .A(n30547), .Y(n34020) );
  AOI21X1 U30091 ( .A(n32020), .B(reg_A[0]), .C(n35601), .Y(n35595) );
  OAI21X1 U30092 ( .A(n35602), .B(n25726), .C(n35603), .Y(n35601) );
  OAI21X1 U30093 ( .A(n35604), .B(n35605), .C(n25382), .Y(n35603) );
  OAI21X1 U30094 ( .A(n35606), .B(n35463), .C(n35607), .Y(n35605) );
  MUX2X1 U30095 ( .B(n35608), .A(n35516), .S(reg_B[23]), .Y(n35607) );
  OAI22X1 U30096 ( .A(n25220), .B(n34822), .C(n27953), .D(n35426), .Y(n35516)
         );
  NOR2X1 U30097 ( .A(n25224), .B(n34822), .Y(n35608) );
  NAND2X1 U30098 ( .A(n35015), .B(n25589), .Y(n34822) );
  INVX1 U30099 ( .A(n34984), .Y(n35015) );
  NAND2X1 U30100 ( .A(reg_B[22]), .B(n35129), .Y(n34984) );
  NAND2X1 U30101 ( .A(reg_B[21]), .B(n25029), .Y(n35463) );
  INVX1 U30102 ( .A(n35149), .Y(n35606) );
  OAI21X1 U30103 ( .A(n30587), .B(n35468), .C(n35609), .Y(n35149) );
  MUX2X1 U30104 ( .B(n35610), .A(n35511), .S(reg_B[23]), .Y(n35609) );
  MUX2X1 U30105 ( .B(n26714), .A(n25232), .S(n34881), .Y(n35511) );
  NOR2X1 U30106 ( .A(n25230), .B(n34881), .Y(n35610) );
  NAND2X1 U30107 ( .A(n34881), .B(n35205), .Y(n35468) );
  OAI22X1 U30108 ( .A(n35391), .B(n35611), .C(n25250), .D(n34837), .Y(n35604)
         );
  NAND2X1 U30109 ( .A(n34826), .B(n35205), .Y(n34837) );
  INVX1 U30110 ( .A(n35426), .Y(n34826) );
  NAND2X1 U30111 ( .A(n34888), .B(n25029), .Y(n35426) );
  INVX1 U30112 ( .A(n35013), .Y(n34888) );
  INVX1 U30113 ( .A(n35612), .Y(n35611) );
  AND2X1 U30114 ( .A(n25052), .B(n34737), .Y(n35391) );
  NAND2X1 U30115 ( .A(n25044), .B(n31782), .Y(n34737) );
  AOI21X1 U30116 ( .A(reg_A[21]), .B(n25751), .C(n35613), .Y(n35602) );
  OAI22X1 U30117 ( .A(n25753), .B(n26714), .C(n25754), .D(n25230), .Y(n35613)
         );
  AOI22X1 U30118 ( .A(n30617), .B(n35591), .C(n25721), .D(reg_A[8]), .Y(n35594) );
  NAND2X1 U30119 ( .A(n35614), .B(n35615), .Y(n35591) );
  AOI22X1 U30120 ( .A(n32934), .B(n34928), .C(n34015), .D(n35616), .Y(n35615)
         );
  OAI21X1 U30121 ( .A(n33807), .B(n25250), .C(n35617), .Y(n34928) );
  AOI22X1 U30122 ( .A(n33923), .B(reg_A[0]), .C(n33919), .D(reg_A[8]), .Y(
        n35617) );
  AOI22X1 U30123 ( .A(n34000), .B(n35133), .C(n33809), .D(n35453), .Y(n35614)
         );
  INVX1 U30124 ( .A(n31828), .Y(n30617) );
  NAND3X1 U30125 ( .A(n35618), .B(n35619), .C(n35620), .Y(n35592) );
  NOR2X1 U30126 ( .A(n35621), .B(n35622), .Y(n35620) );
  OAI21X1 U30127 ( .A(n27839), .B(n35526), .C(n35623), .Y(n35622) );
  AND2X1 U30128 ( .A(n35624), .B(n35625), .Y(n35623) );
  OAI21X1 U30129 ( .A(n35626), .B(n35627), .C(n25310), .Y(n35625) );
  NAND3X1 U30130 ( .A(n35628), .B(n35629), .C(n35630), .Y(n35627) );
  NOR2X1 U30131 ( .A(n35631), .B(n35632), .Y(n35630) );
  OAI22X1 U30132 ( .A(n25250), .B(n25228), .C(n25239), .D(n25229), .Y(n35632)
         );
  OAI22X1 U30133 ( .A(n25244), .B(n25231), .C(n27954), .D(n25482), .Y(n35631)
         );
  AOI22X1 U30134 ( .A(reg_A[24]), .B(n25124), .C(n25222), .D(reg_A[27]), .Y(
        n35629) );
  AOI22X1 U30135 ( .A(n25637), .B(reg_A[26]), .C(n25234), .D(reg_A[30]), .Y(
        n35628) );
  NAND3X1 U30136 ( .A(n35633), .B(n35634), .C(n35635), .Y(n35626) );
  NOR2X1 U30137 ( .A(n35636), .B(n35637), .Y(n35635) );
  OAI22X1 U30138 ( .A(n25033), .B(n25230), .C(n25133), .D(n25224), .Y(n35637)
         );
  OAI22X1 U30139 ( .A(n25041), .B(n25220), .C(n25042), .D(n27953), .Y(n35636)
         );
  AOI22X1 U30140 ( .A(reg_A[23]), .B(n25628), .C(reg_A[20]), .D(n25067), .Y(
        n35634) );
  AOI22X1 U30141 ( .A(reg_A[21]), .B(n25123), .C(n25629), .D(reg_A[25]), .Y(
        n35633) );
  OAI21X1 U30142 ( .A(n27844), .B(n35528), .C(reg_A[16]), .Y(n35624) );
  OAI22X1 U30143 ( .A(n35013), .B(n34903), .C(n26147), .D(n35145), .Y(n35528)
         );
  NAND2X1 U30144 ( .A(n33890), .B(n34493), .Y(n35145) );
  NAND2X1 U30145 ( .A(n26186), .B(n35205), .Y(n34903) );
  INVX1 U30146 ( .A(reg_B[23]), .Y(n35205) );
  NAND2X1 U30147 ( .A(n35129), .B(n34881), .Y(n35013) );
  INVX1 U30148 ( .A(reg_B[22]), .Y(n34881) );
  INVX1 U30149 ( .A(reg_B[21]), .Y(n35129) );
  NAND3X1 U30150 ( .A(n25795), .B(n25032), .C(n35638), .Y(n27844) );
  AOI21X1 U30151 ( .A(n30910), .B(n26801), .C(n35639), .Y(n35638) );
  OAI21X1 U30152 ( .A(reg_B[3]), .B(n35345), .C(n35640), .Y(n35526) );
  AOI22X1 U30153 ( .A(n26530), .B(n35641), .C(n25026), .D(n33987), .Y(n35640)
         );
  MUX2X1 U30154 ( .B(reg_A[6]), .A(reg_A[14]), .S(n26596), .Y(n33987) );
  INVX1 U30155 ( .A(n35642), .Y(n35641) );
  INVX1 U30156 ( .A(n35643), .Y(n35345) );
  OAI21X1 U30157 ( .A(reg_A[16]), .B(n27857), .C(n35644), .Y(n35643) );
  AOI22X1 U30158 ( .A(n27859), .B(n26701), .C(reg_B[2]), .D(n34298), .Y(n35644) );
  NAND3X1 U30159 ( .A(n35645), .B(n35646), .C(n35647), .Y(n35621) );
  OAI21X1 U30160 ( .A(n35648), .B(n35649), .C(n25730), .Y(n35647) );
  NAND3X1 U30161 ( .A(n35650), .B(n35651), .C(n35652), .Y(n35649) );
  NOR2X1 U30162 ( .A(n35653), .B(n35654), .Y(n35652) );
  OAI22X1 U30163 ( .A(n25736), .B(n25250), .C(n25239), .D(n25737), .Y(n35654)
         );
  OAI22X1 U30164 ( .A(n25244), .B(n25738), .C(n27954), .D(n25739), .Y(n35653)
         );
  AOI22X1 U30165 ( .A(reg_A[24]), .B(n25615), .C(n25616), .D(reg_A[27]), .Y(
        n35651) );
  AOI22X1 U30166 ( .A(n25607), .B(reg_A[26]), .C(n25608), .D(reg_A[30]), .Y(
        n35650) );
  NAND3X1 U30167 ( .A(n35655), .B(n35656), .C(n35657), .Y(n35648) );
  NOR2X1 U30168 ( .A(n35658), .B(n35659), .Y(n35657) );
  OAI22X1 U30169 ( .A(n25061), .B(n25230), .C(n25746), .D(n25224), .Y(n35659)
         );
  OAI22X1 U30170 ( .A(n25747), .B(n25220), .C(n25748), .D(n27953), .Y(n35658)
         );
  AOI22X1 U30171 ( .A(reg_A[23]), .B(n25613), .C(reg_A[20]), .D(n25749), .Y(
        n35656) );
  AOI22X1 U30172 ( .A(reg_A[21]), .B(n25750), .C(n25614), .D(reg_A[25]), .Y(
        n35655) );
  OAI21X1 U30173 ( .A(n35660), .B(n35661), .C(n25840), .Y(n35645) );
  NAND3X1 U30174 ( .A(n35662), .B(n35663), .C(n35664), .Y(n35661) );
  NOR2X1 U30175 ( .A(n35665), .B(n35666), .Y(n35664) );
  OAI22X1 U30176 ( .A(n25250), .B(n25228), .C(n25130), .D(n25229), .Y(n35666)
         );
  OAI22X1 U30177 ( .A(n30569), .B(n25231), .C(n25177), .D(n25482), .Y(n35665)
         );
  AOI22X1 U30178 ( .A(n25124), .B(reg_A[8]), .C(n25222), .D(reg_A[5]), .Y(
        n35663) );
  AOI22X1 U30179 ( .A(n25637), .B(reg_A[6]), .C(n25234), .D(reg_A[2]), .Y(
        n35662) );
  NAND3X1 U30180 ( .A(n35667), .B(n35668), .C(n35669), .Y(n35660) );
  NOR2X1 U30181 ( .A(n35670), .B(n35671), .Y(n35669) );
  OAI22X1 U30182 ( .A(n25147), .B(n25131), .C(n25040), .D(n25208), .Y(n35671)
         );
  OAI21X1 U30183 ( .A(n25041), .B(n25206), .C(n35672), .Y(n35670) );
  AOI22X1 U30184 ( .A(n25247), .B(reg_A[0]), .C(reg_A[15]), .D(n25135), .Y(
        n35672) );
  AOI22X1 U30185 ( .A(n25628), .B(reg_A[9]), .C(n25069), .D(reg_A[12]), .Y(
        n35668) );
  AOI22X1 U30186 ( .A(n25123), .B(reg_A[11]), .C(n25629), .D(reg_A[7]), .Y(
        n35667) );
  AOI21X1 U30187 ( .A(n27861), .B(reg_A[1]), .C(n35673), .Y(n35619) );
  OAI22X1 U30188 ( .A(n25146), .B(n35674), .C(n35675), .D(n28058), .Y(n35673)
         );
  AOI22X1 U30189 ( .A(n35676), .B(n31782), .C(n27921), .D(n35677), .Y(n35618)
         );
  OAI21X1 U30190 ( .A(n27925), .B(n35340), .C(n35678), .Y(n35677) );
  AOI22X1 U30191 ( .A(n35679), .B(n26008), .C(n35527), .D(n25751), .Y(n35678)
         );
  INVX1 U30192 ( .A(n33800), .Y(n35340) );
  MUX2X1 U30193 ( .B(n29279), .A(n25132), .S(reg_B[1]), .Y(n33800) );
  OAI21X1 U30194 ( .A(n33964), .B(n35559), .C(n35680), .Y(n35676) );
  AOI22X1 U30195 ( .A(n35681), .B(n34217), .C(n35147), .D(n35682), .Y(n35680)
         );
  INVX1 U30196 ( .A(n35435), .Y(n35682) );
  MUX2X1 U30197 ( .B(n35326), .A(n34464), .S(reg_B[29]), .Y(n35435) );
  MUX2X1 U30198 ( .B(n27967), .A(n25130), .S(reg_B[28]), .Y(n34464) );
  MUX2X1 U30199 ( .B(n29279), .A(n25132), .S(reg_B[28]), .Y(n35326) );
  INVX1 U30200 ( .A(n35683), .Y(n35147) );
  MUX2X1 U30201 ( .B(n25206), .A(n29265), .S(reg_B[28]), .Y(n34217) );
  NOR2X1 U30202 ( .A(reg_B[29]), .B(n27943), .Y(n35681) );
  OAI21X1 U30203 ( .A(reg_B[30]), .B(n35684), .C(n35685), .Y(n35559) );
  AOI22X1 U30204 ( .A(n35686), .B(n34015), .C(n34000), .D(n33971), .Y(n35685)
         );
  MUX2X1 U30205 ( .B(reg_A[6]), .A(reg_A[14]), .S(n34493), .Y(n33971) );
  MUX2X1 U30206 ( .B(reg_A[10]), .A(reg_A[2]), .S(reg_B[28]), .Y(n35686) );
  INVX1 U30207 ( .A(n35322), .Y(n35684) );
  OAI21X1 U30208 ( .A(reg_A[16]), .B(n34230), .C(n35687), .Y(n35322) );
  AOI22X1 U30209 ( .A(reg_B[29]), .B(n35438), .C(n34180), .D(n26701), .Y(
        n35687) );
  INVX1 U30210 ( .A(n34306), .Y(n35438) );
  MUX2X1 U30211 ( .B(n25255), .A(n30569), .S(reg_B[28]), .Y(n34306) );
  OR2X1 U30212 ( .A(n35688), .B(n35689), .Y(result[15]) );
  NAND3X1 U30213 ( .A(n35690), .B(n35691), .C(n35692), .Y(n35689) );
  NOR2X1 U30214 ( .A(n35693), .B(n35694), .Y(n35692) );
  OAI21X1 U30215 ( .A(n25994), .B(n35695), .C(n35696), .Y(n35694) );
  AOI22X1 U30216 ( .A(n25948), .B(reg_A[11]), .C(n35697), .D(n32116), .Y(
        n35696) );
  INVX1 U30217 ( .A(n35698), .Y(n35697) );
  NAND2X1 U30218 ( .A(n35699), .B(n35700), .Y(n35693) );
  AOI22X1 U30219 ( .A(n30634), .B(n35701), .C(n25172), .D(n35702), .Y(n35700)
         );
  AOI22X1 U30220 ( .A(n32052), .B(reg_A[14]), .C(n25947), .D(reg_A[10]), .Y(
        n35699) );
  AOI21X1 U30221 ( .A(n25170), .B(n35703), .C(n35704), .Y(n35691) );
  OAI22X1 U30222 ( .A(n28031), .B(n30559), .C(n32135), .D(n29279), .Y(n35704)
         );
  OAI21X1 U30223 ( .A(n35705), .B(n31806), .C(n35706), .Y(n35703) );
  AOI22X1 U30224 ( .A(n35707), .B(n26733), .C(n25604), .D(n35708), .Y(n35706)
         );
  OAI21X1 U30225 ( .A(n35709), .B(n25194), .C(n35710), .Y(n35708) );
  AOI22X1 U30226 ( .A(n25172), .B(n35711), .C(n26733), .D(n35712), .Y(n35710)
         );
  NOR2X1 U30227 ( .A(n35713), .B(n26999), .Y(n35707) );
  NOR2X1 U30228 ( .A(n35714), .B(n35715), .Y(n35690) );
  OAI21X1 U30229 ( .A(n28066), .B(n26742), .C(n35716), .Y(n35715) );
  OAI21X1 U30230 ( .A(n35717), .B(n35718), .C(n25999), .Y(n35716) );
  NAND2X1 U30231 ( .A(n35719), .B(n35720), .Y(n35718) );
  AOI22X1 U30232 ( .A(n26002), .B(reg_A[8]), .C(reg_A[11]), .D(n26003), .Y(
        n35720) );
  AOI22X1 U30233 ( .A(reg_A[10]), .B(n25751), .C(reg_A[15]), .D(n26004), .Y(
        n35719) );
  NAND2X1 U30234 ( .A(n35721), .B(n35722), .Y(n35717) );
  AOI22X1 U30235 ( .A(reg_A[14]), .B(n26007), .C(reg_A[12]), .D(n26008), .Y(
        n35722) );
  AOI22X1 U30236 ( .A(reg_A[13]), .B(n26009), .C(reg_A[9]), .D(n26010), .Y(
        n35721) );
  MUX2X1 U30237 ( .B(n35723), .A(n35724), .S(reg_B[14]), .Y(n35714) );
  INVX1 U30238 ( .A(n35725), .Y(n35724) );
  NAND2X1 U30239 ( .A(n25188), .B(n35726), .Y(n35723) );
  OAI22X1 U30240 ( .A(n26723), .B(n35727), .C(n25196), .D(n35728), .Y(n35726)
         );
  INVX1 U30241 ( .A(n35729), .Y(n35727) );
  NAND3X1 U30242 ( .A(n35730), .B(n35731), .C(n35732), .Y(n35688) );
  NOR2X1 U30243 ( .A(n35733), .B(n35734), .Y(n35732) );
  OAI21X1 U30244 ( .A(n35735), .B(n26692), .C(n35736), .Y(n35734) );
  AOI21X1 U30245 ( .A(n35737), .B(n35600), .C(n35738), .Y(n35736) );
  AOI21X1 U30246 ( .A(n35739), .B(n35740), .C(n26996), .Y(n35738) );
  AOI22X1 U30247 ( .A(n33923), .B(n33806), .C(n25101), .D(n35394), .Y(n35740)
         );
  NOR2X1 U30248 ( .A(n33915), .B(n27954), .Y(n33806) );
  INVX1 U30249 ( .A(n34751), .Y(n33923) );
  AOI22X1 U30250 ( .A(n30644), .B(n34808), .C(n26772), .D(n34809), .Y(n35739)
         );
  NAND2X1 U30251 ( .A(n35741), .B(n35742), .Y(n35600) );
  AOI22X1 U30252 ( .A(n32934), .B(n35019), .C(n34015), .D(n35743), .Y(n35742)
         );
  OAI22X1 U30253 ( .A(n33807), .B(n29279), .C(n25132), .D(n34465), .Y(n35019)
         );
  AOI22X1 U30254 ( .A(n34000), .B(n35355), .C(n33809), .D(n35589), .Y(n35741)
         );
  AOI21X1 U30255 ( .A(reg_A[15]), .B(n35744), .C(n35745), .Y(n35735) );
  OAI21X1 U30256 ( .A(n35746), .B(n25697), .C(n35747), .Y(n35745) );
  NAND3X1 U30257 ( .A(reg_B[13]), .B(n35748), .C(reg_A[11]), .Y(n35747) );
  OAI21X1 U30258 ( .A(n35749), .B(n25697), .C(n25031), .Y(n35748) );
  AOI22X1 U30259 ( .A(n29245), .B(reg_A[7]), .C(n34083), .D(reg_A[3]), .Y(
        n35746) );
  INVX1 U30260 ( .A(n28026), .Y(n29245) );
  OAI21X1 U30261 ( .A(n28105), .B(n25112), .C(n35750), .Y(n35744) );
  OAI21X1 U30262 ( .A(n28052), .B(n29958), .C(n35751), .Y(n35733) );
  AOI22X1 U30263 ( .A(n35752), .B(n28138), .C(n35753), .D(n35754), .Y(n35751)
         );
  INVX1 U30264 ( .A(n28058), .Y(n35753) );
  NAND2X1 U30265 ( .A(n30634), .B(reg_B[29]), .Y(n28058) );
  NOR2X1 U30266 ( .A(n35755), .B(n35756), .Y(n35731) );
  OAI21X1 U30267 ( .A(n33977), .B(n35757), .C(n35758), .Y(n35756) );
  OAI21X1 U30268 ( .A(n35759), .B(n35760), .C(n25119), .Y(n35758) );
  NAND3X1 U30269 ( .A(n35761), .B(n35762), .C(n35763), .Y(n35760) );
  AOI21X1 U30270 ( .A(n25125), .B(reg_A[15]), .C(n35764), .Y(n35763) );
  OAI22X1 U30271 ( .A(n25128), .B(n25229), .C(n25130), .D(n25231), .Y(n35764)
         );
  AOI22X1 U30272 ( .A(n25124), .B(reg_A[7]), .C(n25222), .D(reg_A[4]), .Y(
        n35762) );
  AOI22X1 U30273 ( .A(n25637), .B(reg_A[5]), .C(n25234), .D(reg_A[1]), .Y(
        n35761) );
  NAND3X1 U30274 ( .A(n35765), .B(n35766), .C(n35767), .Y(n35759) );
  NOR2X1 U30275 ( .A(n35768), .B(n35769), .Y(n35767) );
  OAI22X1 U30276 ( .A(n25146), .B(n25131), .C(n25040), .D(n25206), .Y(n35769)
         );
  OAI22X1 U30277 ( .A(n25041), .B(n25255), .C(n25042), .D(n25208), .Y(n35768)
         );
  AOI22X1 U30278 ( .A(n25628), .B(reg_A[8]), .C(n25069), .D(reg_A[11]), .Y(
        n35766) );
  AOI22X1 U30279 ( .A(n25123), .B(reg_A[10]), .C(n25629), .D(reg_A[6]), .Y(
        n35765) );
  NAND2X1 U30280 ( .A(n25932), .B(n35133), .Y(n35757) );
  OAI21X1 U30281 ( .A(n35683), .B(n35770), .C(n35646), .Y(n35755) );
  NAND2X1 U30282 ( .A(reg_B[29]), .B(n35616), .Y(n35770) );
  NAND2X1 U30283 ( .A(n25142), .B(n25932), .Y(n35683) );
  AOI21X1 U30284 ( .A(n35771), .B(n35772), .C(n35773), .Y(n35730) );
  NAND2X1 U30285 ( .A(n35774), .B(n35775), .Y(n35773) );
  OAI21X1 U30286 ( .A(n35776), .B(n35777), .C(n25918), .Y(n35775) );
  NAND3X1 U30287 ( .A(n35778), .B(n35779), .C(n35780), .Y(n35777) );
  NOR2X1 U30288 ( .A(n35781), .B(n35782), .Y(n35780) );
  OAI22X1 U30289 ( .A(n25736), .B(n29279), .C(n25128), .D(n25737), .Y(n35782)
         );
  OAI22X1 U30290 ( .A(n25130), .B(n25738), .C(n26742), .D(n25739), .Y(n35781)
         );
  AOI22X1 U30291 ( .A(n25615), .B(reg_A[7]), .C(n25616), .D(reg_A[4]), .Y(
        n35779) );
  AOI22X1 U30292 ( .A(n25607), .B(reg_A[5]), .C(n25608), .D(reg_A[1]), .Y(
        n35778) );
  NAND3X1 U30293 ( .A(n35783), .B(n35784), .C(n35785), .Y(n35776) );
  NOR2X1 U30294 ( .A(n35786), .B(n35787), .Y(n35785) );
  OAI22X1 U30295 ( .A(n25745), .B(n25146), .C(n25746), .D(n25206), .Y(n35787)
         );
  OAI22X1 U30296 ( .A(n25747), .B(n25255), .C(n25748), .D(n25208), .Y(n35786)
         );
  AOI22X1 U30297 ( .A(n25613), .B(reg_A[8]), .C(reg_A[11]), .D(n25749), .Y(
        n35784) );
  AOI22X1 U30298 ( .A(reg_A[10]), .B(n25750), .C(n25614), .D(reg_A[6]), .Y(
        n35783) );
  OAI21X1 U30299 ( .A(n35788), .B(n35789), .C(n25310), .Y(n35774) );
  NAND3X1 U30300 ( .A(n35790), .B(n35791), .C(n35792), .Y(n35789) );
  NOR2X1 U30301 ( .A(n35793), .B(n35794), .Y(n35792) );
  OAI22X1 U30302 ( .A(n29279), .B(n25228), .C(n25244), .D(n25229), .Y(n35794)
         );
  OAI22X1 U30303 ( .A(n32918), .B(n25231), .C(n29286), .D(n25482), .Y(n35793)
         );
  AOI22X1 U30304 ( .A(reg_A[24]), .B(n25629), .C(n25222), .D(reg_A[26]), .Y(
        n35791) );
  AOI22X1 U30305 ( .A(n25637), .B(reg_A[25]), .C(n25234), .D(reg_A[29]), .Y(
        n35790) );
  NAND3X1 U30306 ( .A(n35795), .B(n35796), .C(n35797), .Y(n35788) );
  NOR2X1 U30307 ( .A(n35798), .B(n35799), .Y(n35797) );
  OAI22X1 U30308 ( .A(n25040), .B(n27953), .C(n25254), .D(n25224), .Y(n35799)
         );
  OAI21X1 U30309 ( .A(n25042), .B(n25250), .C(n35800), .Y(n35798) );
  AOI21X1 U30310 ( .A(reg_A[31]), .B(n25247), .C(n33881), .Y(n35800) );
  INVX1 U30311 ( .A(n33826), .Y(n33881) );
  NAND2X1 U30312 ( .A(reg_A[23]), .B(n25124), .Y(n33826) );
  AOI22X1 U30313 ( .A(reg_A[21]), .B(n25253), .C(reg_A[22]), .D(n25628), .Y(
        n35796) );
  AOI22X1 U30314 ( .A(reg_A[19]), .B(n25073), .C(reg_A[20]), .D(n25123), .Y(
        n35795) );
  OR2X1 U30315 ( .A(n35801), .B(n35802), .Y(result[14]) );
  NAND3X1 U30316 ( .A(n35803), .B(n35804), .C(n35805), .Y(n35802) );
  NOR2X1 U30317 ( .A(n35806), .B(n35807), .Y(n35805) );
  OAI21X1 U30318 ( .A(n35808), .B(n30547), .C(n35809), .Y(n35807) );
  AOI22X1 U30319 ( .A(n31830), .B(n34147), .C(n26045), .D(n35810), .Y(n35809)
         );
  NAND3X1 U30320 ( .A(n35811), .B(n35812), .C(n35813), .Y(n35810) );
  NOR2X1 U30321 ( .A(n35814), .B(n35815), .Y(n35813) );
  OAI21X1 U30322 ( .A(n25206), .B(n28303), .C(n35816), .Y(n35815) );
  OAI21X1 U30323 ( .A(n35817), .B(n35818), .C(n25604), .Y(n35816) );
  NAND2X1 U30324 ( .A(n35819), .B(n35820), .Y(n35818) );
  AOI22X1 U30325 ( .A(n25607), .B(reg_A[4]), .C(n25608), .D(reg_A[0]), .Y(
        n35820) );
  AOI22X1 U30326 ( .A(n25609), .B(reg_A[2]), .C(n25610), .D(reg_A[1]), .Y(
        n35819) );
  NAND2X1 U30327 ( .A(n35821), .B(n35822), .Y(n35817) );
  AOI22X1 U30328 ( .A(n25613), .B(reg_A[7]), .C(n25614), .D(reg_A[5]), .Y(
        n35822) );
  AOI22X1 U30329 ( .A(n25615), .B(reg_A[6]), .C(n25616), .D(reg_A[3]), .Y(
        n35821) );
  OAI22X1 U30330 ( .A(n26701), .B(n28311), .C(n25146), .D(n25449), .Y(n35814)
         );
  AOI22X1 U30331 ( .A(n25442), .B(reg_A[11]), .C(n27387), .D(reg_A[10]), .Y(
        n35812) );
  AOI22X1 U30332 ( .A(n28312), .B(reg_A[12]), .C(reg_A[14]), .D(n25434), .Y(
        n35811) );
  NAND2X1 U30333 ( .A(n25699), .B(reg_B[31]), .Y(n30547) );
  INVX1 U30334 ( .A(n35823), .Y(n35808) );
  OR2X1 U30335 ( .A(n35824), .B(n35825), .Y(n35806) );
  OAI21X1 U30336 ( .A(n28276), .B(n25255), .C(n35826), .Y(n35825) );
  OAI21X1 U30337 ( .A(n35827), .B(n35828), .C(n25119), .Y(n35826) );
  NAND3X1 U30338 ( .A(n35829), .B(n35830), .C(n35831), .Y(n35828) );
  AOI21X1 U30339 ( .A(n25125), .B(reg_A[14]), .C(n35832), .Y(n35831) );
  OAI22X1 U30340 ( .A(n25177), .B(n25229), .C(n25128), .D(n25231), .Y(n35832)
         );
  AOI22X1 U30341 ( .A(n25629), .B(reg_A[5]), .C(n25124), .D(reg_A[6]), .Y(
        n35830) );
  AOI22X1 U30342 ( .A(n25222), .B(reg_A[3]), .C(n25637), .D(reg_A[4]), .Y(
        n35829) );
  NAND3X1 U30343 ( .A(n35833), .B(n35834), .C(n35835), .Y(n35827) );
  AOI21X1 U30344 ( .A(n25123), .B(reg_A[9]), .C(n35836), .Y(n35835) );
  OAI22X1 U30345 ( .A(n25147), .B(n26431), .C(n25132), .D(n25129), .Y(n35836)
         );
  AOI22X1 U30346 ( .A(reg_A[13]), .B(n25135), .C(reg_A[11]), .D(n25136), .Y(
        n35834) );
  AOI22X1 U30347 ( .A(n25252), .B(reg_A[12]), .C(n25253), .D(reg_A[8]), .Y(
        n35833) );
  OAI22X1 U30348 ( .A(n32135), .B(n25208), .C(n30226), .D(n25147), .Y(n35824)
         );
  INVX1 U30349 ( .A(n26026), .Y(n30226) );
  NOR2X1 U30350 ( .A(n35837), .B(n35838), .Y(n35804) );
  OAI22X1 U30351 ( .A(n29279), .B(n25148), .C(n26421), .D(n35839), .Y(n35838)
         );
  OAI22X1 U30352 ( .A(n35840), .B(n25194), .C(n35841), .D(n25189), .Y(n35837)
         );
  NOR2X1 U30353 ( .A(n35842), .B(n35843), .Y(n35803) );
  OAI22X1 U30354 ( .A(n26041), .B(n25146), .C(n32203), .D(n26701), .Y(n35843)
         );
  OAI22X1 U30355 ( .A(n32204), .B(n26742), .C(n35705), .D(n31828), .Y(n35842)
         );
  NAND2X1 U30356 ( .A(n25699), .B(n33865), .Y(n31828) );
  AND2X1 U30357 ( .A(n35844), .B(n35845), .Y(n35705) );
  AOI22X1 U30358 ( .A(n34015), .B(n35846), .C(n34000), .D(n35453), .Y(n35845)
         );
  NAND2X1 U30359 ( .A(reg_B[30]), .B(n33955), .Y(n34167) );
  AOI22X1 U30360 ( .A(n32934), .B(n35133), .C(n33809), .D(n35616), .Y(n35844)
         );
  INVX1 U30361 ( .A(n28281), .Y(n32204) );
  NAND3X1 U30362 ( .A(n35847), .B(n35848), .C(n35849), .Y(n35801) );
  NOR2X1 U30363 ( .A(n35850), .B(n35851), .Y(n35849) );
  NAND3X1 U30364 ( .A(n35852), .B(n35853), .C(n35854), .Y(n35851) );
  AOI22X1 U30365 ( .A(n25116), .B(n35855), .C(reg_A[11]), .D(n35856), .Y(
        n35854) );
  OAI21X1 U30366 ( .A(n35857), .B(n35858), .C(n35859), .Y(n35856) );
  NAND2X1 U30367 ( .A(n26186), .B(reg_B[15]), .Y(n35858) );
  INVX1 U30368 ( .A(n35860), .Y(n35855) );
  AOI21X1 U30369 ( .A(n35711), .B(n26267), .C(n35702), .Y(n35860) );
  OAI21X1 U30370 ( .A(n35750), .B(n25208), .C(n35861), .Y(n35702) );
  NAND3X1 U30371 ( .A(reg_B[13]), .B(n26504), .C(reg_A[10]), .Y(n35861) );
  NAND2X1 U30372 ( .A(n35862), .B(n35863), .Y(n35711) );
  AOI22X1 U30373 ( .A(n35864), .B(reg_A[2]), .C(n35865), .D(reg_A[6]), .Y(
        n35863) );
  AOI22X1 U30374 ( .A(reg_A[10]), .B(n26691), .C(reg_A[14]), .D(n31796), .Y(
        n35862) );
  OR2X1 U30375 ( .A(n26731), .B(n35866), .Y(n35853) );
  AOI22X1 U30376 ( .A(n35712), .B(n26267), .C(n29315), .D(n35867), .Y(n35866)
         );
  OAI21X1 U30377 ( .A(n35868), .B(n35869), .C(n25310), .Y(n35852) );
  NAND3X1 U30378 ( .A(n35870), .B(n35871), .C(n35872), .Y(n35869) );
  NOR2X1 U30379 ( .A(n35873), .B(n35874), .Y(n35872) );
  OAI22X1 U30380 ( .A(n25244), .B(n25475), .C(n25036), .D(n27962), .Y(n35874)
         );
  OAI21X1 U30381 ( .A(n27960), .B(n25473), .C(n35875), .Y(n35873) );
  AOI22X1 U30382 ( .A(reg_A[23]), .B(n25629), .C(reg_A[22]), .D(n25124), .Y(
        n35875) );
  AOI22X1 U30383 ( .A(n25235), .B(reg_A[29]), .C(n25635), .D(reg_A[26]), .Y(
        n35871) );
  AOI22X1 U30384 ( .A(n25325), .B(reg_A[27]), .C(n25125), .D(reg_A[14]), .Y(
        n35870) );
  NAND3X1 U30385 ( .A(n35876), .B(n35877), .C(n35878), .Y(n35868) );
  NOR2X1 U30386 ( .A(n35879), .B(n35880), .Y(n35878) );
  OAI22X1 U30387 ( .A(n25040), .B(n25250), .C(n25041), .D(n27953), .Y(n35880)
         );
  OAI21X1 U30388 ( .A(n25042), .B(n29279), .C(n35881), .Y(n35879) );
  AOI22X1 U30389 ( .A(reg_A[31]), .B(n25246), .C(reg_A[30]), .D(n25247), .Y(
        n35881) );
  AOI22X1 U30390 ( .A(reg_A[20]), .B(n25253), .C(reg_A[21]), .D(n25628), .Y(
        n35877) );
  AOI22X1 U30391 ( .A(reg_A[18]), .B(n25074), .C(reg_A[19]), .D(n25123), .Y(
        n35876) );
  NAND3X1 U30392 ( .A(n35882), .B(n35646), .C(n35883), .Y(n35850) );
  AOI22X1 U30393 ( .A(n35884), .B(n26186), .C(n35885), .D(n35886), .Y(n35883)
         );
  INVX1 U30394 ( .A(n35887), .Y(n35886) );
  NOR2X1 U30395 ( .A(n25032), .B(n35728), .Y(n35885) );
  AND2X1 U30396 ( .A(n29302), .B(n35772), .Y(n35884) );
  OAI21X1 U30397 ( .A(n25208), .B(n35888), .C(n35889), .Y(n35772) );
  MUX2X1 U30398 ( .B(n35890), .A(n35891), .S(reg_B[14]), .Y(n35889) );
  NOR2X1 U30399 ( .A(n26723), .B(n25147), .Y(n35890) );
  NOR2X1 U30400 ( .A(n35892), .B(n35893), .Y(n35848) );
  INVX1 U30401 ( .A(n35894), .Y(n35893) );
  AOI22X1 U30402 ( .A(n35701), .B(n29316), .C(n29246), .D(n35895), .Y(n35894)
         );
  OAI21X1 U30403 ( .A(reg_B[29]), .B(n35896), .C(n35897), .Y(n35701) );
  OAI21X1 U30404 ( .A(n26145), .B(n35898), .C(n35899), .Y(n35892) );
  OAI21X1 U30405 ( .A(n30650), .B(n28332), .C(reg_A[13]), .Y(n35899) );
  NOR2X1 U30406 ( .A(n26727), .B(n26731), .Y(n30650) );
  INVX1 U30407 ( .A(n35900), .Y(n35898) );
  AOI21X1 U30408 ( .A(n25932), .B(n35901), .C(n35902), .Y(n35847) );
  OAI21X1 U30409 ( .A(n28057), .B(n35903), .C(n35904), .Y(n35902) );
  OAI21X1 U30410 ( .A(n35905), .B(n35906), .C(n26480), .Y(n35904) );
  OAI22X1 U30411 ( .A(n29239), .B(n28033), .C(n34906), .D(n25099), .Y(n35906)
         );
  OAI22X1 U30412 ( .A(n34494), .B(n25106), .C(n34016), .D(n35907), .Y(n35905)
         );
  INVX1 U30413 ( .A(n34908), .Y(n34016) );
  INVX1 U30414 ( .A(n34909), .Y(n34494) );
  NAND2X1 U30415 ( .A(n25188), .B(reg_B[13]), .Y(n28057) );
  NAND2X1 U30416 ( .A(n35908), .B(n35909), .Y(n35901) );
  AOI22X1 U30417 ( .A(n34015), .B(n35754), .C(n33890), .D(n35133), .Y(n35909)
         );
  OAI22X1 U30418 ( .A(n33807), .B(n25208), .C(n26677), .D(n34465), .Y(n35133)
         );
  INVX1 U30419 ( .A(n29255), .Y(n34015) );
  NAND2X1 U30420 ( .A(reg_B[30]), .B(reg_B[29]), .Y(n29255) );
  AOI22X1 U30421 ( .A(reg_B[31]), .B(n35823), .C(n35910), .D(n35616), .Y(
        n35908) );
  NAND3X1 U30422 ( .A(n35911), .B(n35912), .C(n35913), .Y(result[13]) );
  NOR2X1 U30423 ( .A(n35914), .B(n35915), .Y(n35913) );
  NAND2X1 U30424 ( .A(n35916), .B(n35917), .Y(n35915) );
  AOI21X1 U30425 ( .A(n31830), .B(n25102), .C(n35918), .Y(n35917) );
  OAI22X1 U30426 ( .A(n25994), .B(n35919), .C(n35920), .D(n27943), .Y(n35918)
         );
  NAND2X1 U30427 ( .A(n35921), .B(n35922), .Y(n25102) );
  AOI22X1 U30428 ( .A(reg_A[13]), .B(n25156), .C(n25142), .D(reg_A[14]), .Y(
        n35922) );
  AOI22X1 U30429 ( .A(reg_A[15]), .B(n25258), .C(reg_A[16]), .D(n26761), .Y(
        n35921) );
  INVX1 U30430 ( .A(n30559), .Y(n31830) );
  AOI21X1 U30431 ( .A(n28343), .B(reg_A[13]), .C(n35923), .Y(n35916) );
  OAI21X1 U30432 ( .A(n35924), .B(n25835), .C(n35925), .Y(n35923) );
  OAI21X1 U30433 ( .A(n35926), .B(n35927), .C(n26045), .Y(n35925) );
  NAND3X1 U30434 ( .A(n35928), .B(n35929), .C(n35930), .Y(n35927) );
  AOI21X1 U30435 ( .A(reg_A[13]), .B(n25434), .C(n35931), .Y(n35930) );
  OAI22X1 U30436 ( .A(n28353), .B(n27967), .C(n25205), .D(n25146), .Y(n35931)
         );
  AOI22X1 U30437 ( .A(n25097), .B(n35932), .C(reg_A[8]), .D(n28355), .Y(n35929) );
  AOI22X1 U30438 ( .A(reg_A[12]), .B(n25441), .C(reg_A[10]), .D(n27241), .Y(
        n35928) );
  NAND3X1 U30439 ( .A(n35933), .B(n35934), .C(n35935), .Y(n35926) );
  NOR2X1 U30440 ( .A(n35936), .B(n35937), .Y(n35935) );
  OAI22X1 U30441 ( .A(n28361), .B(n26742), .C(n25132), .D(n28311), .Y(n35937)
         );
  OAI22X1 U30442 ( .A(n25130), .B(n28362), .C(n25128), .D(n28363), .Y(n35936)
         );
  AOI22X1 U30443 ( .A(n28364), .B(reg_A[1]), .C(n25500), .D(reg_A[4]), .Y(
        n35934) );
  AOI22X1 U30444 ( .A(n25501), .B(reg_A[5]), .C(n25502), .D(reg_A[6]), .Y(
        n35933) );
  INVX1 U30445 ( .A(n35932), .Y(n35924) );
  NAND3X1 U30446 ( .A(n35938), .B(n35939), .C(n35940), .Y(n35932) );
  NOR2X1 U30447 ( .A(n35941), .B(n35942), .Y(n35940) );
  OAI21X1 U30448 ( .A(n25206), .B(n25043), .C(n35943), .Y(n35942) );
  AOI22X1 U30449 ( .A(n25637), .B(reg_A[3]), .C(n25635), .D(reg_A[1]), .Y(
        n35943) );
  OAI21X1 U30450 ( .A(n25128), .B(n25473), .C(n35944), .Y(n35941) );
  AOI22X1 U30451 ( .A(n25629), .B(reg_A[4]), .C(n25124), .D(reg_A[5]), .Y(
        n35944) );
  NOR2X1 U30452 ( .A(n35945), .B(n35946), .Y(n35939) );
  OAI22X1 U30453 ( .A(n25132), .B(n25131), .C(n25040), .D(n27967), .Y(n35946)
         );
  OAI22X1 U30454 ( .A(n25147), .B(n25254), .C(n25784), .D(n25255), .Y(n35945)
         );
  AOI21X1 U30455 ( .A(n25123), .B(reg_A[8]), .C(n35947), .Y(n35938) );
  OAI22X1 U30456 ( .A(n25146), .B(n26431), .C(n26677), .D(n25129), .Y(n35947)
         );
  NAND3X1 U30457 ( .A(n35948), .B(n35949), .C(n35950), .Y(n35914) );
  AOI21X1 U30458 ( .A(n28280), .B(reg_A[14]), .C(n35951), .Y(n35950) );
  OAI22X1 U30459 ( .A(n29279), .B(n28569), .C(n26854), .D(n35695), .Y(n35951)
         );
  OAI21X1 U30460 ( .A(n35952), .B(n26452), .C(n35953), .Y(n35695) );
  AOI22X1 U30461 ( .A(n26293), .B(n34207), .C(n26295), .D(n34298), .Y(n35953)
         );
  INVX1 U30462 ( .A(n35445), .Y(n34298) );
  MUX2X1 U30463 ( .B(n25255), .A(n30569), .S(reg_B[1]), .Y(n35445) );
  INVX1 U30464 ( .A(n35679), .Y(n34207) );
  MUX2X1 U30465 ( .B(n25206), .A(n29265), .S(reg_B[1]), .Y(n35679) );
  INVX1 U30466 ( .A(n35954), .Y(n35952) );
  AOI22X1 U30467 ( .A(n35823), .B(n35737), .C(n32356), .D(reg_A[10]), .Y(
        n35949) );
  OAI21X1 U30468 ( .A(n25697), .B(n32935), .C(n33964), .Y(n35737) );
  NAND2X1 U30469 ( .A(n25932), .B(n33865), .Y(n33964) );
  OAI21X1 U30470 ( .A(n35955), .B(n34176), .C(n35956), .Y(n35823) );
  AOI22X1 U30471 ( .A(n32934), .B(n35355), .C(n33809), .D(n35743), .Y(n35956)
         );
  OAI22X1 U30472 ( .A(n33807), .B(n25206), .C(n29265), .D(n34465), .Y(n35355)
         );
  AOI22X1 U30473 ( .A(n35725), .B(n29256), .C(n26734), .D(n35957), .Y(n35948)
         );
  OAI22X1 U30474 ( .A(n35958), .B(n35959), .C(n25342), .D(n35960), .Y(n35725)
         );
  MUX2X1 U30475 ( .B(n35867), .A(n35891), .S(reg_B[15]), .Y(n35960) );
  OAI21X1 U30476 ( .A(n35961), .B(n26723), .C(n25188), .Y(n35959) );
  OAI22X1 U30477 ( .A(n35962), .B(n35728), .C(n29304), .D(n35963), .Y(n35958)
         );
  MUX2X1 U30478 ( .B(n25206), .A(n25255), .S(reg_B[15]), .Y(n35963) );
  NOR2X1 U30479 ( .A(n35964), .B(n35965), .Y(n35912) );
  OAI21X1 U30480 ( .A(n26278), .B(n35698), .C(n35966), .Y(n35965) );
  AOI22X1 U30481 ( .A(n35771), .B(n35967), .C(n35968), .D(n35969), .Y(n35966)
         );
  INVX1 U30482 ( .A(n35970), .Y(n35967) );
  NAND2X1 U30483 ( .A(n35971), .B(n35972), .Y(n35698) );
  AOI22X1 U30484 ( .A(n26292), .B(n25146), .C(n26293), .D(n25206), .Y(n35972)
         );
  AOI22X1 U30485 ( .A(n26294), .B(n26701), .C(n26295), .D(n25255), .Y(n35971)
         );
  NAND3X1 U30486 ( .A(n35973), .B(n35974), .C(n35975), .Y(n35964) );
  AND2X1 U30487 ( .A(n35646), .B(n35882), .Y(n35975) );
  NAND3X1 U30488 ( .A(reg_B[13]), .B(n25114), .C(reg_B[14]), .Y(n35882) );
  OAI21X1 U30489 ( .A(n35976), .B(n35977), .C(n25310), .Y(n35974) );
  NAND3X1 U30490 ( .A(n35978), .B(n35979), .C(n35980), .Y(n35977) );
  NOR2X1 U30491 ( .A(n35981), .B(n35982), .Y(n35980) );
  OAI22X1 U30492 ( .A(n32918), .B(n25475), .C(n25036), .D(n26714), .Y(n35982)
         );
  OAI21X1 U30493 ( .A(n25027), .B(n27962), .C(n35983), .Y(n35981) );
  AOI22X1 U30494 ( .A(reg_A[22]), .B(n25629), .C(reg_A[21]), .D(n25124), .Y(
        n35983) );
  AOI22X1 U30495 ( .A(n25235), .B(reg_A[28]), .C(n25635), .D(reg_A[25]), .Y(
        n35979) );
  AOI22X1 U30496 ( .A(n25325), .B(reg_A[26]), .C(n25125), .D(reg_A[13]), .Y(
        n35978) );
  NAND3X1 U30497 ( .A(n35984), .B(n35985), .C(n35986), .Y(n35976) );
  NOR2X1 U30498 ( .A(n35987), .B(n35988), .Y(n35986) );
  OAI22X1 U30499 ( .A(n25041), .B(n25250), .C(n25784), .D(n25208), .Y(n35988)
         );
  OAI21X1 U30500 ( .A(n25051), .B(n27954), .C(n35989), .Y(n35987) );
  AOI22X1 U30501 ( .A(reg_A[30]), .B(n25246), .C(reg_A[29]), .D(n25247), .Y(
        n35989) );
  AOI21X1 U30502 ( .A(reg_A[20]), .B(n25628), .C(n35990), .Y(n35985) );
  OAI22X1 U30503 ( .A(n25033), .B(n25220), .C(n25040), .D(n29279), .Y(n35990)
         );
  AOI22X1 U30504 ( .A(reg_A[17]), .B(n25073), .C(reg_A[18]), .D(n25123), .Y(
        n35984) );
  NAND2X1 U30505 ( .A(reg_A[11]), .B(n35991), .Y(n35973) );
  OAI21X1 U30506 ( .A(n25189), .B(n35992), .C(n28415), .Y(n35991) );
  NOR2X1 U30507 ( .A(n35993), .B(n35994), .Y(n35911) );
  OAI21X1 U30508 ( .A(n26701), .B(n28434), .C(n35995), .Y(n35994) );
  AOI22X1 U30509 ( .A(n26267), .B(n35996), .C(n25170), .D(n35997), .Y(n35995)
         );
  OAI22X1 U30510 ( .A(n35998), .B(n31806), .C(n35999), .D(n36000), .Y(n35997)
         );
  AOI22X1 U30511 ( .A(n35867), .B(n29256), .C(n36001), .D(reg_A[11]), .Y(
        n35999) );
  INVX1 U30512 ( .A(n35713), .Y(n35867) );
  MUX2X1 U30513 ( .B(reg_A[13]), .A(reg_A[9]), .S(reg_B[13]), .Y(n35713) );
  NAND2X1 U30514 ( .A(reg_B[31]), .B(n25044), .Y(n31806) );
  OAI21X1 U30515 ( .A(n36002), .B(n25189), .C(n36003), .Y(n35996) );
  AOI22X1 U30516 ( .A(n25116), .B(n35712), .C(n25172), .D(n36004), .Y(n36003)
         );
  NAND2X1 U30517 ( .A(n36005), .B(n36006), .Y(n35712) );
  AOI22X1 U30518 ( .A(n35865), .B(reg_A[5]), .C(reg_A[13]), .D(n31796), .Y(
        n36006) );
  AOI22X1 U30519 ( .A(n35864), .B(reg_A[1]), .C(reg_A[9]), .D(n26691), .Y(
        n36005) );
  NAND3X1 U30520 ( .A(n36007), .B(n36008), .C(n36009), .Y(n35993) );
  AOI22X1 U30521 ( .A(n35895), .B(n35288), .C(n28453), .D(reg_A[0]), .Y(n36009) );
  OAI21X1 U30522 ( .A(n25206), .B(n26692), .C(n36010), .Y(n35288) );
  AOI22X1 U30523 ( .A(reg_A[15]), .B(n26733), .C(reg_A[14]), .D(n25172), .Y(
        n36010) );
  OAI21X1 U30524 ( .A(n36011), .B(n36012), .C(n26480), .Y(n36008) );
  OAI22X1 U30525 ( .A(n25098), .B(n28033), .C(n35020), .D(n35907), .Y(n36012)
         );
  INVX1 U30526 ( .A(n25109), .Y(n35020) );
  OAI21X1 U30527 ( .A(n29305), .B(n27954), .C(n36013), .Y(n25109) );
  AOI22X1 U30528 ( .A(reg_A[29]), .B(n25156), .C(n25142), .D(reg_A[30]), .Y(
        n36013) );
  INVX1 U30529 ( .A(n30643), .Y(n25098) );
  NAND2X1 U30530 ( .A(n36014), .B(n36015), .Y(n30643) );
  AOI22X1 U30531 ( .A(reg_A[17]), .B(n25156), .C(n25142), .D(reg_A[18]), .Y(
        n36015) );
  AOI22X1 U30532 ( .A(reg_A[19]), .B(n25258), .C(reg_A[20]), .D(n26761), .Y(
        n36014) );
  OAI22X1 U30533 ( .A(n36016), .B(n25106), .C(n25105), .D(n25099), .Y(n36011)
         );
  INVX1 U30534 ( .A(n35022), .Y(n25105) );
  NAND2X1 U30535 ( .A(n36017), .B(n36018), .Y(n35022) );
  AOI22X1 U30536 ( .A(reg_A[21]), .B(n25156), .C(n25142), .D(reg_A[22]), .Y(
        n36018) );
  AOI22X1 U30537 ( .A(reg_A[23]), .B(n25258), .C(reg_A[24]), .D(n26761), .Y(
        n36017) );
  INVX1 U30538 ( .A(n25104), .Y(n36016) );
  NAND2X1 U30539 ( .A(n36019), .B(n36020), .Y(n25104) );
  AOI22X1 U30540 ( .A(reg_A[25]), .B(n25156), .C(n25142), .D(reg_A[26]), .Y(
        n36020) );
  AOI22X1 U30541 ( .A(reg_A[27]), .B(n25258), .C(reg_A[28]), .D(n26761), .Y(
        n36019) );
  OAI21X1 U30542 ( .A(n36021), .B(n36022), .C(n25932), .Y(n36007) );
  OAI22X1 U30543 ( .A(n36023), .B(n30648), .C(n26758), .D(n35897), .Y(n36022)
         );
  NAND2X1 U30544 ( .A(reg_B[29]), .B(n25262), .Y(n30648) );
  NOR2X1 U30545 ( .A(n35896), .B(n33977), .Y(n36021) );
  INVX1 U30546 ( .A(n35453), .Y(n35896) );
  NAND2X1 U30547 ( .A(n36024), .B(n36025), .Y(result[12]) );
  NOR2X1 U30548 ( .A(n36026), .B(n36027), .Y(n36025) );
  NAND3X1 U30549 ( .A(n36028), .B(n36029), .C(n36030), .Y(n36027) );
  NOR2X1 U30550 ( .A(n36031), .B(n36032), .Y(n36030) );
  OAI21X1 U30551 ( .A(n36033), .B(n25697), .C(n36034), .Y(n36032) );
  OAI21X1 U30552 ( .A(n36035), .B(n36036), .C(n26480), .Y(n36034) );
  OAI22X1 U30553 ( .A(n35126), .B(n25099), .C(n34726), .D(n25106), .Y(n36036)
         );
  INVX1 U30554 ( .A(n26778), .Y(n34726) );
  INVX1 U30555 ( .A(n26773), .Y(n35126) );
  OAI22X1 U30556 ( .A(n26769), .B(n28033), .C(n34284), .D(n35907), .Y(n36035)
         );
  INVX1 U30557 ( .A(n26777), .Y(n34284) );
  INVX1 U30558 ( .A(n36037), .Y(n26769) );
  AOI21X1 U30559 ( .A(n36038), .B(n36039), .C(n36040), .Y(n36033) );
  OAI22X1 U30560 ( .A(n35998), .B(n32935), .C(n35970), .D(n36000), .Y(n36040)
         );
  AOI22X1 U30561 ( .A(reg_A[10]), .B(n36001), .C(n29256), .D(n35891), .Y(
        n35970) );
  MUX2X1 U30562 ( .B(n25255), .A(n26701), .S(reg_B[13]), .Y(n35891) );
  INVX1 U30563 ( .A(n35857), .Y(n36001) );
  NAND2X1 U30564 ( .A(n25044), .B(n33865), .Y(n32935) );
  INVX1 U30565 ( .A(n36041), .Y(n35998) );
  OAI21X1 U30566 ( .A(n35920), .B(n34176), .C(n36042), .Y(n36041) );
  AOI22X1 U30567 ( .A(n33809), .B(n35846), .C(n32934), .D(n35453), .Y(n36042)
         );
  NAND2X1 U30568 ( .A(reg_B[29]), .B(n34176), .Y(n33966) );
  INVX1 U30569 ( .A(n36043), .Y(n36031) );
  AOI22X1 U30570 ( .A(n36044), .B(n25159), .C(n36045), .D(n25168), .Y(n36043)
         );
  AOI22X1 U30571 ( .A(n25932), .B(n36046), .C(n25188), .D(n36047), .Y(n36029)
         );
  OAI21X1 U30572 ( .A(n35728), .B(n26686), .C(n36048), .Y(n36047) );
  INVX1 U30573 ( .A(n36049), .Y(n36048) );
  OAI21X1 U30574 ( .A(n26726), .B(n30552), .C(n36050), .Y(n36049) );
  NAND2X1 U30575 ( .A(n36051), .B(n36052), .Y(n26726) );
  AOI22X1 U30576 ( .A(n26733), .B(n26677), .C(n25172), .D(n25132), .Y(n36052)
         );
  AOI22X1 U30577 ( .A(n26734), .B(n29265), .C(n25116), .D(n26701), .Y(n36051)
         );
  NAND2X1 U30578 ( .A(n36053), .B(n36054), .Y(n26686) );
  AOI22X1 U30579 ( .A(n26733), .B(n25128), .C(n25172), .D(n25130), .Y(n36054)
         );
  AOI22X1 U30580 ( .A(n26734), .B(n25177), .C(n25116), .D(n30569), .Y(n36053)
         );
  OAI21X1 U30581 ( .A(n35920), .B(n29305), .C(n36055), .Y(n36046) );
  AOI22X1 U30582 ( .A(n36056), .B(n25156), .C(n33890), .D(n35453), .Y(n36055)
         );
  OAI22X1 U30583 ( .A(n33807), .B(n25255), .C(n30569), .D(n34465), .Y(n35453)
         );
  INVX1 U30584 ( .A(n35897), .Y(n36056) );
  NAND2X1 U30585 ( .A(n25101), .B(reg_A[8]), .Y(n35897) );
  INVX1 U30586 ( .A(n36057), .Y(n36028) );
  OAI22X1 U30587 ( .A(n26692), .B(n35841), .C(n26731), .D(n35840), .Y(n36057)
         );
  AOI22X1 U30588 ( .A(n36058), .B(n26267), .C(n36059), .D(reg_A[11]), .Y(
        n35840) );
  AOI22X1 U30589 ( .A(n36004), .B(n26267), .C(n36059), .D(reg_A[12]), .Y(
        n35841) );
  INVX1 U30590 ( .A(n35709), .Y(n36004) );
  NOR2X1 U30591 ( .A(n36060), .B(n36061), .Y(n35709) );
  OAI22X1 U30592 ( .A(n26701), .B(n30552), .C(n29304), .D(n25255), .Y(n36061)
         );
  OAI21X1 U30593 ( .A(n30569), .B(n35728), .C(n36050), .Y(n36060) );
  NAND3X1 U30594 ( .A(n36062), .B(n36063), .C(n36064), .Y(n36026) );
  NOR2X1 U30595 ( .A(n36065), .B(n36066), .Y(n36064) );
  OAI21X1 U30596 ( .A(n36067), .B(n25147), .C(n36068), .Y(n36066) );
  OAI21X1 U30597 ( .A(n36069), .B(n36070), .C(n25310), .Y(n36068) );
  NAND3X1 U30598 ( .A(n36071), .B(n36072), .C(n36073), .Y(n36070) );
  NOR2X1 U30599 ( .A(n36074), .B(n36075), .Y(n36073) );
  OAI22X1 U30600 ( .A(n25255), .B(n25228), .C(n27960), .D(n25229), .Y(n36075)
         );
  OAI21X1 U30601 ( .A(n27962), .B(n25231), .C(n36076), .Y(n36074) );
  AOI22X1 U30602 ( .A(n25234), .B(reg_A[26]), .C(n25235), .D(reg_A[27]), .Y(
        n36076) );
  AOI21X1 U30603 ( .A(reg_A[20]), .B(n25124), .C(n36077), .Y(n36072) );
  OAI22X1 U30604 ( .A(n25037), .B(n25232), .C(n25028), .D(n27953), .Y(n36077)
         );
  AOI22X1 U30605 ( .A(reg_A[23]), .B(n25222), .C(reg_A[22]), .D(n25637), .Y(
        n36071) );
  NAND3X1 U30606 ( .A(n36078), .B(n36079), .C(n36080), .Y(n36069) );
  NOR2X1 U30607 ( .A(n36081), .B(n36082), .Y(n36080) );
  OAI22X1 U30608 ( .A(n25042), .B(n25206), .C(n25331), .D(n29286), .Y(n36082)
         );
  OAI21X1 U30609 ( .A(n25038), .B(n27954), .C(n36083), .Y(n36081) );
  AOI22X1 U30610 ( .A(reg_A[29]), .B(n25246), .C(reg_A[28]), .D(n25247), .Y(
        n36083) );
  AOI21X1 U30611 ( .A(reg_A[18]), .B(n25253), .C(n36084), .Y(n36079) );
  OAI22X1 U30612 ( .A(n25040), .B(n25208), .C(n25041), .D(n29279), .Y(n36084)
         );
  AOI22X1 U30613 ( .A(reg_A[19]), .B(n25628), .C(n25070), .D(reg_A[16]), .Y(
        n36078) );
  AOI21X1 U30614 ( .A(n26733), .B(n36059), .C(n28496), .Y(n36067) );
  OAI21X1 U30615 ( .A(n25198), .B(n36085), .C(n36086), .Y(n36065) );
  OAI21X1 U30616 ( .A(n36087), .B(n36088), .C(n25119), .Y(n36086) );
  OR2X1 U30617 ( .A(n36089), .B(n36090), .Y(n36088) );
  OAI21X1 U30618 ( .A(n30569), .B(n25467), .C(n36091), .Y(n36090) );
  AOI22X1 U30619 ( .A(n25253), .B(reg_A[6]), .C(n25628), .D(reg_A[5]), .Y(
        n36091) );
  OAI21X1 U30620 ( .A(n25128), .B(n25219), .C(n36092), .Y(n36089) );
  AOI22X1 U30621 ( .A(n25629), .B(reg_A[3]), .C(n25222), .D(reg_A[1]), .Y(
        n36092) );
  OR2X1 U30622 ( .A(n36093), .B(n36094), .Y(n36087) );
  OAI21X1 U30623 ( .A(n25255), .B(n25043), .C(n36095), .Y(n36094) );
  AOI22X1 U30624 ( .A(reg_A[11]), .B(n25135), .C(n25252), .D(reg_A[10]), .Y(
        n36095) );
  OAI21X1 U30625 ( .A(n25132), .B(n26703), .C(n36096), .Y(n36093) );
  AOI22X1 U30626 ( .A(n25136), .B(reg_A[9]), .C(n25069), .D(reg_A[8]), .Y(
        n36096) );
  AOI22X1 U30627 ( .A(n25142), .B(n36097), .C(n26761), .D(n36098), .Y(n36085)
         );
  AOI22X1 U30628 ( .A(reg_A[9]), .B(n36099), .C(n35895), .D(n26779), .Y(n36063) );
  OAI21X1 U30629 ( .A(n35750), .B(n25194), .C(n32433), .Y(n36099) );
  INVX1 U30630 ( .A(n36059), .Y(n35750) );
  NAND2X1 U30631 ( .A(n26727), .B(n35992), .Y(n36059) );
  NAND2X1 U30632 ( .A(n25188), .B(n31796), .Y(n26727) );
  AOI22X1 U30633 ( .A(n28549), .B(reg_A[1]), .C(n28649), .D(reg_A[2]), .Y(
        n36062) );
  NOR2X1 U30634 ( .A(n36100), .B(n36101), .Y(n36024) );
  NAND3X1 U30635 ( .A(n36102), .B(n36103), .C(n36104), .Y(n36101) );
  NOR2X1 U30636 ( .A(n36105), .B(n36106), .Y(n36104) );
  OAI21X1 U30637 ( .A(n29265), .B(n28562), .C(n25088), .Y(n36106) );
  OAI22X1 U30638 ( .A(n31780), .B(n30559), .C(n32494), .D(n26701), .Y(n36105)
         );
  INVX1 U30639 ( .A(n26771), .Y(n31780) );
  AOI22X1 U30640 ( .A(n25153), .B(reg_A[14]), .C(n28280), .D(reg_A[13]), .Y(
        n36103) );
  AOI22X1 U30641 ( .A(reg_A[11]), .B(n26358), .C(reg_A[12]), .D(n28563), .Y(
        n36102) );
  NAND3X1 U30642 ( .A(n36107), .B(n36108), .C(n36109), .Y(n36100) );
  NOR2X1 U30643 ( .A(n36110), .B(n36111), .Y(n36109) );
  OAI22X1 U30644 ( .A(n29279), .B(n28570), .C(n25132), .D(n28571), .Y(n36111)
         );
  OAI22X1 U30645 ( .A(n30569), .B(n25178), .C(n26677), .D(n28714), .Y(n36110)
         );
  AOI22X1 U30646 ( .A(reg_A[0]), .B(n28494), .C(n28572), .D(reg_A[3]), .Y(
        n36108) );
  INVX1 U30647 ( .A(n36112), .Y(n36107) );
  OAI22X1 U30648 ( .A(n26741), .B(n26421), .C(n26728), .D(n26420), .Y(n36112)
         );
  NAND2X1 U30649 ( .A(n36113), .B(n36114), .Y(n26728) );
  AOI22X1 U30650 ( .A(n26601), .B(n26677), .C(n26602), .D(n29265), .Y(n36114)
         );
  AOI22X1 U30651 ( .A(n27012), .B(n26701), .C(n26597), .D(n25132), .Y(n36113)
         );
  NAND2X1 U30652 ( .A(n36115), .B(n36116), .Y(n26741) );
  AOI22X1 U30653 ( .A(n26601), .B(n25128), .C(n26602), .D(n25177), .Y(n36116)
         );
  AOI22X1 U30654 ( .A(n27012), .B(n30569), .C(n26597), .D(n25130), .Y(n36115)
         );
  NAND3X1 U30655 ( .A(n36117), .B(n36118), .C(n36119), .Y(result[127]) );
  NOR2X1 U30656 ( .A(n36120), .B(n36121), .Y(n36119) );
  NAND3X1 U30657 ( .A(n36122), .B(n36123), .C(n36124), .Y(n36121) );
  AOI21X1 U30658 ( .A(n25999), .B(n36125), .C(n36126), .Y(n36124) );
  OAI21X1 U30659 ( .A(n25994), .B(n36127), .C(n36128), .Y(n36126) );
  OAI21X1 U30660 ( .A(n36129), .B(n36130), .C(n25170), .Y(n36128) );
  OAI21X1 U30661 ( .A(n36131), .B(n36132), .C(n36133), .Y(n36130) );
  NAND2X1 U30662 ( .A(n25044), .B(n36134), .Y(n36133) );
  OAI21X1 U30663 ( .A(n36135), .B(n36136), .C(n36137), .Y(n36134) );
  OAI21X1 U30664 ( .A(n36138), .B(n36139), .C(n25793), .Y(n36137) );
  OAI22X1 U30665 ( .A(n36140), .B(n25549), .C(n25452), .D(n36141), .Y(n36139)
         );
  INVX1 U30666 ( .A(n36142), .Y(n36138) );
  AOI22X1 U30667 ( .A(n36143), .B(reg_B[125]), .C(reg_A[103]), .D(n36144), .Y(
        n36142) );
  OAI21X1 U30668 ( .A(n36136), .B(n36145), .C(n36146), .Y(n36129) );
  OAI21X1 U30669 ( .A(n36147), .B(n25393), .C(n36148), .Y(n36146) );
  INVX1 U30670 ( .A(n36149), .Y(n36147) );
  OR2X1 U30671 ( .A(n26999), .B(n36150), .Y(n36145) );
  NAND3X1 U30672 ( .A(n36151), .B(n36152), .C(n36153), .Y(n36125) );
  NOR2X1 U30673 ( .A(n36154), .B(n36155), .Y(n36153) );
  OAI22X1 U30674 ( .A(n26943), .B(n25497), .C(n26944), .D(n25494), .Y(n36155)
         );
  OAI22X1 U30675 ( .A(n26945), .B(n25321), .C(n25753), .D(n25493), .Y(n36154)
         );
  AOI22X1 U30676 ( .A(reg_A[126]), .B(n26007), .C(reg_A[124]), .D(n26008), .Y(
        n36152) );
  AOI22X1 U30677 ( .A(reg_A[125]), .B(n26009), .C(reg_A[121]), .D(n26010), .Y(
        n36151) );
  AOI22X1 U30678 ( .A(n25948), .B(reg_A[123]), .C(reg_A[127]), .D(n29972), .Y(
        n36123) );
  OAI21X1 U30679 ( .A(n25063), .B(n36156), .C(n36157), .Y(n29972) );
  NOR2X1 U30680 ( .A(n26179), .B(n36158), .Y(n36157) );
  NAND2X1 U30681 ( .A(n27676), .B(n26004), .Y(n36156) );
  AOI22X1 U30682 ( .A(n36159), .B(n32116), .C(n36160), .D(n26260), .Y(n36122)
         );
  NAND3X1 U30683 ( .A(n36161), .B(n36162), .C(n36163), .Y(n36120) );
  AOI21X1 U30684 ( .A(reg_B[127]), .B(n36164), .C(n36165), .Y(n36163) );
  OAI21X1 U30685 ( .A(n36166), .B(n26147), .C(n36167), .Y(n36165) );
  OAI21X1 U30686 ( .A(n36168), .B(n36169), .C(n25932), .Y(n36167) );
  OAI22X1 U30687 ( .A(n25356), .B(n36170), .C(n36136), .D(n36171), .Y(n36169)
         );
  OAI21X1 U30688 ( .A(n36172), .B(n36173), .C(n36174), .Y(n36168) );
  OAI21X1 U30689 ( .A(n36175), .B(n36176), .C(n25793), .Y(n36174) );
  OAI22X1 U30690 ( .A(n36177), .B(n36178), .C(n36179), .D(n36180), .Y(n36176)
         );
  NOR2X1 U30691 ( .A(n36140), .B(n25549), .Y(n36175) );
  AOI22X1 U30692 ( .A(reg_A[126]), .B(n36181), .C(n25840), .D(n36182), .Y(
        n36162) );
  NAND2X1 U30693 ( .A(n36183), .B(n36184), .Y(n36182) );
  NOR2X1 U30694 ( .A(n36185), .B(n36186), .Y(n36184) );
  NAND3X1 U30695 ( .A(n36187), .B(n36188), .C(n36189), .Y(n36186) );
  NOR2X1 U30696 ( .A(n36190), .B(n36191), .Y(n36189) );
  OAI22X1 U30697 ( .A(n25059), .B(n25670), .C(n25318), .D(n25436), .Y(n36191)
         );
  OAI22X1 U30698 ( .A(n25320), .B(n25448), .C(n25322), .D(n25361), .Y(n36190)
         );
  AOI22X1 U30699 ( .A(n25631), .B(reg_A[97]), .C(n25764), .D(reg_A[96]), .Y(
        n36188) );
  AOI22X1 U30700 ( .A(n25324), .B(reg_A[99]), .C(n25765), .D(reg_A[98]), .Y(
        n36187) );
  NAND3X1 U30701 ( .A(n36192), .B(n36193), .C(n36194), .Y(n36185) );
  NOR2X1 U30702 ( .A(n36195), .B(n36196), .Y(n36194) );
  OAI22X1 U30703 ( .A(n25051), .B(n25474), .C(n25038), .D(n25469), .Y(n36196)
         );
  OAI22X1 U30704 ( .A(n25048), .B(n25452), .C(n25336), .D(n25450), .Y(n36195)
         );
  AOI22X1 U30705 ( .A(reg_A[105]), .B(n25242), .C(reg_A[104]), .D(n25338), .Y(
        n36193) );
  AOI22X1 U30706 ( .A(reg_A[107]), .B(n25339), .C(reg_A[106]), .D(n25257), .Y(
        n36192) );
  NOR2X1 U30707 ( .A(n36197), .B(n36198), .Y(n36183) );
  NAND3X1 U30708 ( .A(n36199), .B(n36200), .C(n36201), .Y(n36198) );
  NOR2X1 U30709 ( .A(n36202), .B(n36203), .Y(n36201) );
  OAI22X1 U30710 ( .A(n25043), .B(n25497), .C(n25039), .D(n25771), .Y(n36203)
         );
  OAI22X1 U30711 ( .A(n25064), .B(n25335), .C(n25482), .D(n25476), .Y(n36202)
         );
  AOI22X1 U30712 ( .A(reg_A[119]), .B(n25124), .C(reg_A[116]), .D(n25222), .Y(
        n36200) );
  AOI22X1 U30713 ( .A(reg_A[117]), .B(n25637), .C(reg_A[113]), .D(n25234), .Y(
        n36199) );
  NAND3X1 U30714 ( .A(n36204), .B(n36205), .C(n36206), .Y(n36197) );
  NOR2X1 U30715 ( .A(n36207), .B(n36208), .Y(n36206) );
  OAI22X1 U30716 ( .A(n25033), .B(n25490), .C(n25040), .D(n25317), .Y(n36208)
         );
  OAI22X1 U30717 ( .A(n25041), .B(n25323), .C(n25042), .D(n25319), .Y(n36207)
         );
  AOI22X1 U30718 ( .A(reg_A[120]), .B(n25628), .C(reg_A[123]), .D(n25068), .Y(
        n36205) );
  AOI22X1 U30719 ( .A(reg_A[122]), .B(n25123), .C(reg_A[118]), .D(n25629), .Y(
        n36204) );
  AOI22X1 U30720 ( .A(n25275), .B(n36209), .C(n36210), .D(reg_A[119]), .Y(
        n36161) );
  INVX1 U30721 ( .A(n30044), .Y(n36210) );
  NAND3X1 U30722 ( .A(n27676), .B(n26004), .C(n26038), .Y(n30044) );
  NOR2X1 U30723 ( .A(n36211), .B(n36212), .Y(n36118) );
  NAND3X1 U30724 ( .A(n36213), .B(n36214), .C(n36215), .Y(n36212) );
  OAI21X1 U30725 ( .A(n36216), .B(n25947), .C(reg_A[122]), .Y(n36215) );
  INVX1 U30726 ( .A(n32117), .Y(n25947) );
  INVX1 U30727 ( .A(n36217), .Y(n36216) );
  OAI21X1 U30728 ( .A(n36218), .B(n36219), .C(n25918), .Y(n36214) );
  NAND3X1 U30729 ( .A(n36220), .B(n36221), .C(n36222), .Y(n36219) );
  NOR2X1 U30730 ( .A(n36223), .B(n36224), .Y(n36222) );
  OAI22X1 U30731 ( .A(n25736), .B(n25497), .C(n25737), .D(n25771), .Y(n36224)
         );
  OAI22X1 U30732 ( .A(n25738), .B(n25335), .C(n25739), .D(n25476), .Y(n36223)
         );
  AOI22X1 U30733 ( .A(reg_A[119]), .B(n25615), .C(reg_A[116]), .D(n25616), .Y(
        n36221) );
  AOI22X1 U30734 ( .A(reg_A[117]), .B(n25607), .C(reg_A[113]), .D(n25608), .Y(
        n36220) );
  NAND3X1 U30735 ( .A(n36225), .B(n36226), .C(n36227), .Y(n36218) );
  NOR2X1 U30736 ( .A(n36228), .B(n36229), .Y(n36227) );
  OAI22X1 U30737 ( .A(n25745), .B(n25490), .C(n25746), .D(n25317), .Y(n36229)
         );
  OAI22X1 U30738 ( .A(n25747), .B(n25323), .C(n25748), .D(n25319), .Y(n36228)
         );
  AOI22X1 U30739 ( .A(reg_A[120]), .B(n25613), .C(reg_A[123]), .D(n25749), .Y(
        n36226) );
  AOI22X1 U30740 ( .A(reg_A[122]), .B(n25750), .C(reg_A[118]), .D(n25614), .Y(
        n36225) );
  NAND2X1 U30741 ( .A(n25188), .B(n36230), .Y(n36213) );
  OAI21X1 U30742 ( .A(n25493), .B(n36231), .C(n36232), .Y(n36230) );
  OAI21X1 U30743 ( .A(n36233), .B(n36234), .C(n36235), .Y(n36232) );
  OAI21X1 U30744 ( .A(n36236), .B(n36170), .C(n36166), .Y(n36234) );
  INVX1 U30745 ( .A(n36237), .Y(n36166) );
  OAI22X1 U30746 ( .A(n36238), .B(n36136), .C(n36239), .D(n25397), .Y(n36237)
         );
  AOI22X1 U30747 ( .A(n36240), .B(reg_A[115]), .C(n36241), .D(reg_A[119]), .Y(
        n36239) );
  INVX1 U30748 ( .A(n36242), .Y(n36233) );
  AOI21X1 U30749 ( .A(n36243), .B(n25700), .C(n36244), .Y(n36242) );
  OAI22X1 U30750 ( .A(n36245), .B(n36246), .C(n36131), .D(n36247), .Y(n36244)
         );
  NAND3X1 U30751 ( .A(n36248), .B(n36249), .C(n36250), .Y(n36211) );
  AOI22X1 U30752 ( .A(n36251), .B(n36252), .C(n36253), .D(n25700), .Y(n36250)
         );
  NOR2X1 U30753 ( .A(n36254), .B(n26610), .Y(n36253) );
  NOR2X1 U30754 ( .A(n36246), .B(n36177), .Y(n36251) );
  NAND3X1 U30755 ( .A(reg_B[126]), .B(n26504), .C(n36255), .Y(n36249) );
  OAI21X1 U30756 ( .A(n36256), .B(n36257), .C(n36148), .Y(n36248) );
  NOR2X1 U30757 ( .A(n36258), .B(n36259), .Y(n36117) );
  OAI21X1 U30758 ( .A(n25323), .B(n36260), .C(n36261), .Y(n36259) );
  AOI22X1 U30759 ( .A(n36262), .B(n25900), .C(n36263), .D(n36264), .Y(n36261)
         );
  INVX1 U30760 ( .A(n36131), .Y(n36264) );
  NOR2X1 U30761 ( .A(n31636), .B(n26943), .Y(n25900) );
  NAND2X1 U30762 ( .A(n36265), .B(n36266), .Y(n36258) );
  AOI22X1 U30763 ( .A(n36267), .B(n25910), .C(n36268), .D(n28138), .Y(n36266)
         );
  INVX1 U30764 ( .A(n29964), .Y(n25910) );
  NAND2X1 U30765 ( .A(n27676), .B(n26003), .Y(n29964) );
  INVX1 U30766 ( .A(n36269), .Y(n36267) );
  AOI22X1 U30767 ( .A(n36270), .B(n29963), .C(n36271), .D(n25935), .Y(n36265)
         );
  INVX1 U30768 ( .A(n29958), .Y(n25935) );
  INVX1 U30769 ( .A(n25939), .Y(n29963) );
  NAND3X1 U30770 ( .A(n36272), .B(n36273), .C(n36274), .Y(result[126]) );
  NOR2X1 U30771 ( .A(n36275), .B(n36276), .Y(n36274) );
  NAND3X1 U30772 ( .A(n36277), .B(n36278), .C(n36279), .Y(n36276) );
  AOI21X1 U30773 ( .A(n36280), .B(n36252), .C(n36281), .Y(n36279) );
  OAI21X1 U30774 ( .A(n25031), .B(n36282), .C(n36283), .Y(n36281) );
  OAI21X1 U30775 ( .A(n36284), .B(n36285), .C(n36286), .Y(n36283) );
  OAI22X1 U30776 ( .A(n36287), .B(n25397), .C(n36136), .D(n36245), .Y(n36285)
         );
  OAI21X1 U30777 ( .A(n36288), .B(n36289), .C(n36290), .Y(n36284) );
  NAND3X1 U30778 ( .A(n36291), .B(n36172), .C(n36292), .Y(n36290) );
  INVX1 U30779 ( .A(n36293), .Y(n36292) );
  NAND2X1 U30780 ( .A(n25355), .B(reg_A[115]), .Y(n36289) );
  AOI22X1 U30781 ( .A(n36294), .B(n36295), .C(n36296), .D(n36263), .Y(n36278)
         );
  AOI22X1 U30782 ( .A(n36297), .B(reg_A[119]), .C(reg_A[125]), .D(n36181), .Y(
        n36277) );
  OR2X1 U30783 ( .A(n32052), .B(n36298), .Y(n36181) );
  NAND3X1 U30784 ( .A(n36299), .B(n36300), .C(n36301), .Y(n36275) );
  AOI21X1 U30785 ( .A(n36302), .B(n36303), .C(n36304), .Y(n36301) );
  OAI21X1 U30786 ( .A(n26145), .B(n36305), .C(n36306), .Y(n36304) );
  OAI21X1 U30787 ( .A(n36158), .B(n26179), .C(reg_A[126]), .Y(n36306) );
  INVX1 U30788 ( .A(n30282), .Y(n26179) );
  INVX1 U30789 ( .A(n36307), .Y(n36158) );
  AOI22X1 U30790 ( .A(n36308), .B(n25700), .C(n25277), .D(n36309), .Y(n36300)
         );
  OAI21X1 U30791 ( .A(reg_B[126]), .B(n36254), .C(n36310), .Y(n36309) );
  INVX1 U30792 ( .A(n36209), .Y(n36310) );
  OAI21X1 U30793 ( .A(n36311), .B(n36312), .C(n36313), .Y(n36209) );
  AOI22X1 U30794 ( .A(n36314), .B(n36315), .C(reg_B[126]), .D(n36316), .Y(
        n36313) );
  INVX1 U30795 ( .A(n36317), .Y(n36316) );
  NOR2X1 U30796 ( .A(n25333), .B(n36318), .Y(n36314) );
  INVX1 U30797 ( .A(n36319), .Y(n36254) );
  OAI21X1 U30798 ( .A(n25356), .B(n25319), .C(n36320), .Y(n36319) );
  AOI22X1 U30799 ( .A(n36144), .B(reg_A[102]), .C(n36321), .D(reg_A[110]), .Y(
        n36320) );
  NOR2X1 U30800 ( .A(n36238), .B(n36322), .Y(n36308) );
  AOI22X1 U30801 ( .A(reg_A[121]), .B(n36323), .C(reg_A[124]), .D(n36324), .Y(
        n36299) );
  OAI21X1 U30802 ( .A(n36136), .B(n36325), .C(n28276), .Y(n36324) );
  NAND2X1 U30803 ( .A(n26041), .B(n36217), .Y(n36323) );
  NAND2X1 U30804 ( .A(n36263), .B(n25700), .Y(n36217) );
  NOR2X1 U30805 ( .A(n36326), .B(n36327), .Y(n36273) );
  OAI21X1 U30806 ( .A(n32203), .B(n25493), .C(n36328), .Y(n36327) );
  AOI22X1 U30807 ( .A(n36329), .B(n36330), .C(n36331), .D(n36256), .Y(n36328)
         );
  INVX1 U30808 ( .A(n36173), .Y(n36330) );
  OAI21X1 U30809 ( .A(n36332), .B(n36312), .C(n36333), .Y(n36173) );
  AOI22X1 U30810 ( .A(n36315), .B(n36334), .C(reg_B[126]), .D(n36335), .Y(
        n36333) );
  OAI21X1 U30811 ( .A(reg_A[118]), .B(n36318), .C(n36336), .Y(n36334) );
  AOI22X1 U30812 ( .A(reg_B[123]), .B(n36337), .C(n36338), .D(n25319), .Y(
        n36336) );
  INVX1 U30813 ( .A(n36339), .Y(n36332) );
  NAND2X1 U30814 ( .A(n36340), .B(n36341), .Y(n36326) );
  AOI22X1 U30815 ( .A(reg_A[123]), .B(n36342), .C(n25275), .D(n36343), .Y(
        n36341) );
  AOI22X1 U30816 ( .A(n36344), .B(n26139), .C(n26408), .D(reg_A[127]), .Y(
        n36340) );
  INVX1 U30817 ( .A(n36345), .Y(n36344) );
  NOR2X1 U30818 ( .A(n36346), .B(n36347), .Y(n36272) );
  NAND2X1 U30819 ( .A(n36348), .B(n36349), .Y(n36347) );
  MUX2X1 U30820 ( .B(n36164), .A(n36350), .S(reg_B[127]), .Y(n36349) );
  AND2X1 U30821 ( .A(n36351), .B(n26186), .Y(n36350) );
  OAI22X1 U30822 ( .A(n36293), .B(n26151), .C(n26147), .D(n36352), .Y(n36164)
         );
  MUX2X1 U30823 ( .B(n36243), .A(n36353), .S(reg_B[126]), .Y(n36352) );
  NAND2X1 U30824 ( .A(n36354), .B(n36287), .Y(n36243) );
  AOI22X1 U30825 ( .A(reg_A[118]), .B(n36241), .C(reg_A[114]), .D(n36240), .Y(
        n36287) );
  AOI22X1 U30826 ( .A(n36355), .B(reg_A[122]), .C(reg_A[126]), .D(n36356), .Y(
        n36354) );
  NOR2X1 U30827 ( .A(n36357), .B(n36358), .Y(n36293) );
  OAI22X1 U30828 ( .A(n25494), .B(n36312), .C(n25319), .D(n36359), .Y(n36358)
         );
  OAI21X1 U30829 ( .A(n25323), .B(n36360), .C(n36282), .Y(n36357) );
  AOI22X1 U30830 ( .A(n26045), .B(n36361), .C(n36257), .D(n36362), .Y(n36348)
         );
  NAND3X1 U30831 ( .A(n36363), .B(n36364), .C(n36365), .Y(n36361) );
  NOR2X1 U30832 ( .A(n36366), .B(n36367), .Y(n36365) );
  OAI22X1 U30833 ( .A(n25598), .B(n25323), .C(n25599), .D(n25321), .Y(n36367)
         );
  OAI21X1 U30834 ( .A(n25600), .B(n25490), .C(n36368), .Y(n36366) );
  OAI21X1 U30835 ( .A(n36369), .B(n36370), .C(n25604), .Y(n36368) );
  NAND2X1 U30836 ( .A(n36371), .B(n36372), .Y(n36370) );
  AOI22X1 U30837 ( .A(reg_A[116]), .B(n25607), .C(reg_A[112]), .D(n25608), .Y(
        n36372) );
  AOI22X1 U30838 ( .A(reg_A[114]), .B(n25609), .C(reg_A[113]), .D(n25610), .Y(
        n36371) );
  NAND2X1 U30839 ( .A(n36373), .B(n36374), .Y(n36369) );
  AOI22X1 U30840 ( .A(reg_A[119]), .B(n25613), .C(reg_A[117]), .D(n25614), .Y(
        n36374) );
  AOI22X1 U30841 ( .A(reg_A[118]), .B(n25615), .C(reg_A[115]), .D(n25616), .Y(
        n36373) );
  AOI21X1 U30842 ( .A(reg_A[125]), .B(n25617), .C(n36375), .Y(n36364) );
  OAI21X1 U30843 ( .A(n25619), .B(n25319), .C(n36376), .Y(n36375) );
  OAI21X1 U30844 ( .A(n36377), .B(n36378), .C(n25044), .Y(n36376) );
  NAND2X1 U30845 ( .A(n36379), .B(n36380), .Y(n36378) );
  NOR2X1 U30846 ( .A(n36381), .B(n36382), .Y(n36380) );
  OAI21X1 U30847 ( .A(n25034), .B(n25333), .C(n36383), .Y(n36382) );
  AOI22X1 U30848 ( .A(reg_A[119]), .B(n25628), .C(reg_A[117]), .D(n25629), .Y(
        n36383) );
  OAI21X1 U30849 ( .A(n25287), .B(n25498), .C(n36384), .Y(n36381) );
  AOI22X1 U30850 ( .A(n25631), .B(reg_A[96]), .C(n25324), .D(reg_A[98]), .Y(
        n36384) );
  NOR2X1 U30851 ( .A(n36385), .B(n36386), .Y(n36379) );
  OAI21X1 U30852 ( .A(n25039), .B(n25483), .C(n36387), .Y(n36386) );
  AOI22X1 U30853 ( .A(reg_A[111]), .B(n25235), .C(reg_A[114]), .D(n25635), .Y(
        n36387) );
  OAI21X1 U30854 ( .A(n25035), .B(n25476), .C(n36388), .Y(n36385) );
  AOI22X1 U30855 ( .A(reg_A[115]), .B(n25222), .C(reg_A[116]), .D(n25637), .Y(
        n36388) );
  NAND2X1 U30856 ( .A(n36389), .B(n36390), .Y(n36377) );
  NOR2X1 U30857 ( .A(n36391), .B(n36392), .Y(n36390) );
  OAI21X1 U30858 ( .A(n25491), .B(n25448), .C(n36393), .Y(n36392) );
  AOI22X1 U30859 ( .A(reg_A[108]), .B(n25241), .C(reg_A[104]), .D(n25242), .Y(
        n36393) );
  OAI21X1 U30860 ( .A(n25038), .B(n25470), .C(n36394), .Y(n36391) );
  AOI22X1 U30861 ( .A(reg_A[109]), .B(n25246), .C(reg_A[110]), .D(n25247), .Y(
        n36394) );
  NOR2X1 U30862 ( .A(n36395), .B(n36396), .Y(n36389) );
  OAI21X1 U30863 ( .A(n25059), .B(n25436), .C(n36397), .Y(n36396) );
  AOI22X1 U30864 ( .A(reg_A[102]), .B(n25647), .C(n25648), .D(reg_A[99]), .Y(
        n36397) );
  OAI21X1 U30865 ( .A(n25322), .B(n25670), .C(n36398), .Y(n36395) );
  AOI22X1 U30866 ( .A(reg_A[106]), .B(n25339), .C(reg_A[105]), .D(n25257), .Y(
        n36398) );
  AOI22X1 U30867 ( .A(reg_A[122]), .B(n25650), .C(reg_A[120]), .D(n25651), .Y(
        n36363) );
  OAI21X1 U30868 ( .A(n26012), .B(n36399), .C(n36400), .Y(n36346) );
  AOI22X1 U30869 ( .A(reg_A[122]), .B(n26026), .C(n36160), .D(n26028), .Y(
        n36400) );
  INVX1 U30870 ( .A(n36401), .Y(n36160) );
  OAI21X1 U30871 ( .A(n36402), .B(n26030), .C(n36403), .Y(n36401) );
  AOI22X1 U30872 ( .A(n26032), .B(n36404), .C(n25025), .D(n36405), .Y(n36403)
         );
  OAI21X1 U30873 ( .A(reg_A[126]), .B(n25063), .C(n36406), .Y(n36404) );
  AOI22X1 U30874 ( .A(n26038), .B(n25333), .C(reg_B[0]), .D(n36407), .Y(n36406) );
  NAND3X1 U30875 ( .A(n36408), .B(n36409), .C(n36410), .Y(result[125]) );
  AND2X1 U30876 ( .A(n36411), .B(n36412), .Y(n36410) );
  NOR2X1 U30877 ( .A(n36413), .B(n36414), .Y(n36412) );
  OAI21X1 U30878 ( .A(n36238), .B(n36415), .C(n36416), .Y(n36414) );
  AOI22X1 U30879 ( .A(n36159), .B(n32319), .C(n36417), .D(n36303), .Y(n36416)
         );
  AND2X1 U30880 ( .A(n36418), .B(n36419), .Y(n36159) );
  AOI22X1 U30881 ( .A(n26292), .B(n25490), .C(n26293), .D(n25317), .Y(n36419)
         );
  AOI22X1 U30882 ( .A(n26294), .B(n25493), .C(n26295), .D(n25323), .Y(n36418)
         );
  AND2X1 U30883 ( .A(n36420), .B(n36421), .Y(n36238) );
  AOI22X1 U30884 ( .A(n36240), .B(reg_A[113]), .C(n36241), .D(reg_A[117]), .Y(
        n36421) );
  AOI22X1 U30885 ( .A(n36355), .B(reg_A[121]), .C(reg_A[125]), .D(n36356), .Y(
        n36420) );
  NAND3X1 U30886 ( .A(n36422), .B(n36423), .C(n36424), .Y(n36413) );
  AOI22X1 U30887 ( .A(n26504), .B(n36425), .C(reg_A[123]), .D(n36426), .Y(
        n36424) );
  OAI21X1 U30888 ( .A(n36136), .B(n36325), .C(n26206), .Y(n36426) );
  INVX1 U30889 ( .A(n33943), .Y(n26206) );
  NAND2X1 U30890 ( .A(n28415), .B(n30486), .Y(n33943) );
  OAI21X1 U30891 ( .A(reg_B[126]), .B(n36427), .C(n36282), .Y(n36425) );
  NAND2X1 U30892 ( .A(n36280), .B(reg_A[120]), .Y(n36282) );
  INVX1 U30893 ( .A(n36255), .Y(n36427) );
  MUX2X1 U30894 ( .B(n36150), .A(n36428), .S(reg_B[127]), .Y(n36255) );
  MUX2X1 U30895 ( .B(reg_A[124]), .A(reg_A[120]), .S(reg_B[125]), .Y(n36428)
         );
  MUX2X1 U30896 ( .B(reg_A[125]), .A(reg_A[121]), .S(reg_B[125]), .Y(n36150)
         );
  NAND3X1 U30897 ( .A(n36241), .B(n36429), .C(n36286), .Y(n36423) );
  NAND3X1 U30898 ( .A(n26267), .B(n36353), .C(n25700), .Y(n36422) );
  NOR2X1 U30899 ( .A(n36430), .B(n36431), .Y(n36411) );
  OAI21X1 U30900 ( .A(n26265), .B(n25493), .C(n36432), .Y(n36431) );
  AOI22X1 U30901 ( .A(n26269), .B(reg_A[121]), .C(n25355), .D(n36433), .Y(
        n36432) );
  INVX1 U30902 ( .A(n34156), .Y(n26265) );
  OAI21X1 U30903 ( .A(n27523), .B(n30355), .C(n28434), .Y(n34156) );
  OAI21X1 U30904 ( .A(n25333), .B(n36434), .C(n36435), .Y(n36430) );
  AOI22X1 U30905 ( .A(n36436), .B(n36343), .C(n36437), .D(n36252), .Y(n36435)
         );
  OAI21X1 U30906 ( .A(n36438), .B(n36439), .C(n36440), .Y(n36343) );
  AOI22X1 U30907 ( .A(n36441), .B(n25428), .C(n36442), .D(n36143), .Y(n36440)
         );
  INVX1 U30908 ( .A(n36135), .Y(n36441) );
  NOR2X1 U30909 ( .A(n36443), .B(n36444), .Y(n36135) );
  OAI22X1 U30910 ( .A(n25356), .B(n25317), .C(n25332), .D(n25549), .Y(n36444)
         );
  OAI21X1 U30911 ( .A(n25474), .B(n36141), .C(n36445), .Y(n36443) );
  AOI22X1 U30912 ( .A(n36144), .B(reg_A[101]), .C(reg_B[125]), .D(n36446), .Y(
        n36445) );
  INVX1 U30913 ( .A(n36447), .Y(n36438) );
  NOR2X1 U30914 ( .A(n36448), .B(n36449), .Y(n36409) );
  OAI21X1 U30915 ( .A(n26525), .B(n36399), .C(n36450), .Y(n36449) );
  AOI22X1 U30916 ( .A(n36329), .B(n36295), .C(reg_A[122]), .D(n30287), .Y(
        n36450) );
  OAI21X1 U30917 ( .A(n27523), .B(n36451), .C(n28379), .Y(n30287) );
  INVX1 U30918 ( .A(n36452), .Y(n36295) );
  OAI21X1 U30919 ( .A(n36453), .B(n36439), .C(n36454), .Y(n36452) );
  AOI22X1 U30920 ( .A(n36171), .B(n25428), .C(n36442), .D(n36178), .Y(n36454)
         );
  NAND2X1 U30921 ( .A(n36455), .B(n36456), .Y(n36171) );
  AOI22X1 U30922 ( .A(n36457), .B(n36458), .C(reg_B[125]), .D(n36459), .Y(
        n36456) );
  AOI22X1 U30923 ( .A(n25409), .B(n25332), .C(n25427), .D(n25317), .Y(n36455)
         );
  OAI21X1 U30924 ( .A(n36460), .B(n26208), .C(n36461), .Y(n36399) );
  AOI22X1 U30925 ( .A(n25026), .B(n36269), .C(n36462), .D(n26030), .Y(n36461)
         );
  INVX1 U30926 ( .A(n36270), .Y(n36462) );
  MUX2X1 U30927 ( .B(n36463), .A(n36464), .S(reg_B[2]), .Y(n36270) );
  OAI21X1 U30928 ( .A(reg_A[125]), .B(n25063), .C(n36465), .Y(n36463) );
  AOI22X1 U30929 ( .A(n26038), .B(n25332), .C(reg_B[0]), .D(n36466), .Y(n36465) );
  OAI21X1 U30930 ( .A(n25319), .B(n26136), .C(n36467), .Y(n36448) );
  AOI22X1 U30931 ( .A(n36468), .B(n25150), .C(n26310), .D(reg_A[127]), .Y(
        n36467) );
  INVX1 U30932 ( .A(n36127), .Y(n36468) );
  NAND2X1 U30933 ( .A(n36469), .B(n36470), .Y(n36127) );
  AOI22X1 U30934 ( .A(n26313), .B(n25323), .C(n26314), .D(n25317), .Y(n36470)
         );
  NOR2X1 U30935 ( .A(n27857), .B(reg_B[4]), .Y(n26314) );
  NOR2X1 U30936 ( .A(n27857), .B(n26863), .Y(n26313) );
  AOI22X1 U30937 ( .A(reg_B[1]), .B(n36471), .C(reg_B[2]), .D(n36472), .Y(
        n36469) );
  INVX1 U30938 ( .A(n36473), .Y(n36471) );
  NOR2X1 U30939 ( .A(n36474), .B(n36475), .Y(n36408) );
  OR2X1 U30940 ( .A(n36476), .B(n36477), .Y(n36475) );
  OAI21X1 U30941 ( .A(n36478), .B(n36479), .C(n36480), .Y(n36477) );
  OAI21X1 U30942 ( .A(n36481), .B(n36482), .C(n26045), .Y(n36480) );
  NAND3X1 U30943 ( .A(n36483), .B(n36484), .C(n36485), .Y(n36482) );
  AOI21X1 U30944 ( .A(reg_A[125]), .B(n25434), .C(n36486), .Y(n36485) );
  OAI22X1 U30945 ( .A(n25321), .B(n25437), .C(n25490), .D(n25438), .Y(n36486)
         );
  AOI22X1 U30946 ( .A(n25439), .B(reg_A[115]), .C(n25440), .D(reg_A[119]), .Y(
        n36484) );
  INVX1 U30947 ( .A(n28311), .Y(n25440) );
  AOI22X1 U30948 ( .A(reg_A[124]), .B(n25441), .C(n25442), .D(reg_A[122]), .Y(
        n36483) );
  NAND3X1 U30949 ( .A(n36487), .B(n36488), .C(n36489), .Y(n36481) );
  NOR2X1 U30950 ( .A(n36490), .B(n36491), .Y(n36489) );
  OAI22X1 U30951 ( .A(n25493), .B(n25449), .C(n25483), .D(n25451), .Y(n36491)
         );
  OAI21X1 U30952 ( .A(n25476), .B(n25453), .C(n36492), .Y(n36490) );
  OAI21X1 U30953 ( .A(n36493), .B(n36494), .C(n25044), .Y(n36492) );
  NAND3X1 U30954 ( .A(n36495), .B(n36496), .C(n36497), .Y(n36494) );
  NOR2X1 U30955 ( .A(n36498), .B(n36499), .Y(n36497) );
  OAI21X1 U30956 ( .A(n25043), .B(n25317), .C(n36500), .Y(n36499) );
  AOI22X1 U30957 ( .A(reg_A[124]), .B(n25135), .C(reg_A[123]), .D(n25252), .Y(
        n36500) );
  NAND2X1 U30958 ( .A(n36501), .B(n36502), .Y(n36498) );
  AOI22X1 U30959 ( .A(reg_A[122]), .B(n25136), .C(reg_A[119]), .D(n25253), .Y(
        n36502) );
  AOI22X1 U30960 ( .A(reg_A[121]), .B(n25074), .C(reg_A[120]), .D(n25123), .Y(
        n36501) );
  NOR2X1 U30961 ( .A(n36503), .B(n36504), .Y(n36496) );
  OAI22X1 U30962 ( .A(n25034), .B(n25332), .C(n25129), .D(n25333), .Y(n36504)
         );
  OAI22X1 U30963 ( .A(n25036), .B(n25335), .C(n25223), .D(n25337), .Y(n36503)
         );
  NOR2X1 U30964 ( .A(n36505), .B(n36506), .Y(n36495) );
  OAI22X1 U30965 ( .A(n25064), .B(n25483), .C(n25473), .D(n25771), .Y(n36506)
         );
  OAI22X1 U30966 ( .A(n25039), .B(n25476), .C(n25475), .D(n25452), .Y(n36505)
         );
  NAND3X1 U30967 ( .A(n36507), .B(n36508), .C(n36509), .Y(n36493) );
  NOR2X1 U30968 ( .A(n36510), .B(n36511), .Y(n36509) );
  OAI21X1 U30969 ( .A(n25065), .B(n25450), .C(n36512), .Y(n36511) );
  AOI22X1 U30970 ( .A(reg_A[108]), .B(n25246), .C(reg_A[109]), .D(n25247), .Y(
        n36512) );
  NAND2X1 U30971 ( .A(n36513), .B(n36514), .Y(n36510) );
  AOI22X1 U30972 ( .A(reg_A[106]), .B(n25487), .C(reg_A[107]), .D(n25241), .Y(
        n36514) );
  AOI22X1 U30973 ( .A(reg_A[105]), .B(n25339), .C(reg_A[104]), .D(n25257), .Y(
        n36513) );
  NOR2X1 U30974 ( .A(n36515), .B(n36516), .Y(n36508) );
  OAI22X1 U30975 ( .A(n25491), .B(n25361), .C(n25492), .D(n25448), .Y(n36516)
         );
  OAI22X1 U30976 ( .A(n25320), .B(n25670), .C(n25322), .D(n25436), .Y(n36515)
         );
  NOR2X1 U30977 ( .A(n36517), .B(n36518), .Y(n36507) );
  OAI22X1 U30978 ( .A(n25396), .B(n25316), .C(n25289), .D(n25318), .Y(n36518)
         );
  OAI22X1 U30979 ( .A(n25424), .B(n25498), .C(n25287), .D(n25499), .Y(n36517)
         );
  AOI22X1 U30980 ( .A(n25500), .B(reg_A[116]), .C(n25501), .D(reg_A[117]), .Y(
        n36488) );
  AOI22X1 U30981 ( .A(n25502), .B(reg_A[118]), .C(n25503), .D(reg_A[114]), .Y(
        n36487) );
  INVX1 U30982 ( .A(n28363), .Y(n25503) );
  MUX2X1 U30983 ( .B(n36519), .A(n36520), .S(reg_B[127]), .Y(n36476) );
  AOI21X1 U30984 ( .A(n36521), .B(n25932), .C(n36522), .Y(n36520) );
  OAI21X1 U30985 ( .A(n36523), .B(n25697), .C(n36524), .Y(n36522) );
  NAND3X1 U30986 ( .A(n36525), .B(n36291), .C(n36286), .Y(n36524) );
  INVX1 U30987 ( .A(n36526), .Y(n36523) );
  NAND2X1 U30988 ( .A(n26186), .B(n36351), .Y(n36519) );
  OAI21X1 U30989 ( .A(n25490), .B(n36312), .C(n36527), .Y(n36351) );
  AOI22X1 U30990 ( .A(n36442), .B(reg_A[123]), .C(n36315), .D(reg_A[125]), .Y(
        n36527) );
  OAI21X1 U30991 ( .A(n25317), .B(n30282), .C(n36528), .Y(n36474) );
  AOI22X1 U30992 ( .A(n36529), .B(n26260), .C(n36530), .D(n26262), .Y(n36528)
         );
  NAND3X1 U30993 ( .A(n36531), .B(n36532), .C(n36533), .Y(result[124]) );
  NOR2X1 U30994 ( .A(n36534), .B(n36535), .Y(n36533) );
  NAND3X1 U30995 ( .A(n36536), .B(n36537), .C(n36538), .Y(n36535) );
  NOR2X1 U30996 ( .A(n36539), .B(n36540), .Y(n36538) );
  OAI21X1 U30997 ( .A(n26393), .B(n25494), .C(n36541), .Y(n36540) );
  OAI21X1 U30998 ( .A(n36542), .B(n36543), .C(n25840), .Y(n36541) );
  NAND3X1 U30999 ( .A(n36544), .B(n36545), .C(n36546), .Y(n36543) );
  NOR2X1 U31000 ( .A(n36547), .B(n36548), .Y(n36546) );
  OAI22X1 U31001 ( .A(n25039), .B(n25452), .C(n25475), .D(n25450), .Y(n36548)
         );
  OAI22X1 U31002 ( .A(n26431), .B(n25493), .C(n25042), .D(n25321), .Y(n36547)
         );
  AOI22X1 U31003 ( .A(reg_A[100]), .B(n25647), .C(n25648), .D(reg_A[97]), .Y(
        n36545) );
  AOI22X1 U31004 ( .A(n26432), .B(reg_A[98]), .C(n25324), .D(reg_A[96]), .Y(
        n36544) );
  NAND3X1 U31005 ( .A(n36549), .B(n36550), .C(n36551), .Y(n36542) );
  NOR2X1 U31006 ( .A(n36552), .B(n36553), .Y(n36551) );
  OAI22X1 U31007 ( .A(n25492), .B(n25361), .C(n25331), .D(n25468), .Y(n36553)
         );
  OAI21X1 U31008 ( .A(n25038), .B(n25296), .C(n36554), .Y(n36552) );
  AOI22X1 U31009 ( .A(reg_A[107]), .B(n25246), .C(reg_A[108]), .D(n25247), .Y(
        n36554) );
  AOI22X1 U31010 ( .A(reg_A[101]), .B(n25338), .C(reg_A[104]), .D(n25339), .Y(
        n36550) );
  AOI22X1 U31011 ( .A(reg_A[103]), .B(n25257), .C(n25857), .D(reg_A[99]), .Y(
        n36549) );
  NOR2X1 U31012 ( .A(n34633), .B(n36555), .Y(n26393) );
  OAI22X1 U31013 ( .A(n26370), .B(n25476), .C(n36556), .D(n36136), .Y(n36539)
         );
  INVX1 U31014 ( .A(n36433), .Y(n36556) );
  OAI22X1 U31015 ( .A(n36557), .B(n26147), .C(n25494), .D(n36325), .Y(n36433)
         );
  NOR2X1 U31016 ( .A(n36558), .B(n26519), .Y(n26370) );
  AOI22X1 U31017 ( .A(n36559), .B(n26139), .C(n36560), .D(n28575), .Y(n36537)
         );
  AOI22X1 U31018 ( .A(n26451), .B(reg_A[127]), .C(n26310), .D(reg_A[126]), .Y(
        n36536) );
  NAND3X1 U31019 ( .A(n36561), .B(n36562), .C(n36563), .Y(n36534) );
  NOR2X1 U31020 ( .A(n36564), .B(n36565), .Y(n36563) );
  OAI21X1 U31021 ( .A(n36566), .B(n25490), .C(n36567), .Y(n36565) );
  OAI21X1 U31022 ( .A(n36298), .B(n26358), .C(reg_A[123]), .Y(n36567) );
  INVX1 U31023 ( .A(n32496), .Y(n26358) );
  NOR2X1 U31024 ( .A(n26472), .B(n36342), .Y(n36566) );
  OR2X1 U31025 ( .A(n28206), .B(n36568), .Y(n36342) );
  OAI21X1 U31026 ( .A(n36246), .B(n36325), .C(n36260), .Y(n36568) );
  OAI21X1 U31027 ( .A(n36172), .B(n36569), .C(n36570), .Y(n36564) );
  NAND2X1 U31028 ( .A(n25170), .B(n36571), .Y(n36569) );
  AOI22X1 U31029 ( .A(reg_A[124]), .B(n36572), .C(n36573), .D(n36526), .Y(
        n36562) );
  OAI21X1 U31030 ( .A(n36574), .B(n26999), .C(n36575), .Y(n36526) );
  OAI21X1 U31031 ( .A(n36576), .B(n36577), .C(n25044), .Y(n36575) );
  OAI22X1 U31032 ( .A(n36311), .B(n36360), .C(reg_B[126]), .D(n36317), .Y(
        n36577) );
  NOR2X1 U31033 ( .A(n36578), .B(n36579), .Y(n36317) );
  OAI22X1 U31034 ( .A(n25356), .B(n25323), .C(n25337), .D(n25549), .Y(n36579)
         );
  OAI21X1 U31035 ( .A(n25469), .B(n36141), .C(n36580), .Y(n36578) );
  AOI22X1 U31036 ( .A(n36144), .B(reg_A[100]), .C(reg_B[125]), .D(n36581), .Y(
        n36580) );
  NOR2X1 U31037 ( .A(n36288), .B(n25551), .Y(n36144) );
  AND2X1 U31038 ( .A(n36582), .B(n36280), .Y(n36576) );
  INVX1 U31039 ( .A(n36525), .Y(n36574) );
  OAI21X1 U31040 ( .A(n25397), .B(n36325), .C(n36583), .Y(n36572) );
  INVX1 U31041 ( .A(n26398), .Y(n36583) );
  NAND3X1 U31042 ( .A(n36307), .B(n30908), .C(n36584), .Y(n26398) );
  AOI22X1 U31043 ( .A(n36585), .B(n36294), .C(n26267), .D(n36586), .Y(n36561)
         );
  OAI21X1 U31044 ( .A(n36587), .B(n36246), .C(n36588), .Y(n36586) );
  AOI22X1 U31045 ( .A(n25793), .B(n36353), .C(n25700), .D(n36303), .Y(n36588)
         );
  OR2X1 U31046 ( .A(n36589), .B(n36590), .Y(n36353) );
  OAI21X1 U31047 ( .A(n36236), .B(n25323), .C(n36245), .Y(n36590) );
  NAND2X1 U31048 ( .A(n36241), .B(reg_A[116]), .Y(n36245) );
  OAI21X1 U31049 ( .A(n25493), .B(n36247), .C(n36591), .Y(n36589) );
  NOR2X1 U31050 ( .A(n36592), .B(n36593), .Y(n36532) );
  NAND2X1 U31051 ( .A(n36594), .B(n36595), .Y(n36593) );
  AOI22X1 U31052 ( .A(n36529), .B(n26028), .C(n36596), .D(n26260), .Y(n36595)
         );
  INVX1 U31053 ( .A(n36597), .Y(n36529) );
  OAI21X1 U31054 ( .A(n36598), .B(n26208), .C(n36599), .Y(n36597) );
  AOI22X1 U31055 ( .A(n25026), .B(n36405), .C(n36600), .D(n26030), .Y(n36599)
         );
  INVX1 U31056 ( .A(n36402), .Y(n36600) );
  MUX2X1 U31057 ( .B(n36601), .A(n36602), .S(reg_B[2]), .Y(n36402) );
  OAI21X1 U31058 ( .A(reg_A[124]), .B(n25063), .C(n36603), .Y(n36601) );
  AOI22X1 U31059 ( .A(n26038), .B(n25337), .C(reg_B[0]), .D(n36604), .Y(n36603) );
  AOI22X1 U31060 ( .A(reg_A[116]), .B(n26551), .C(reg_A[119]), .D(n26353), .Y(
        n36594) );
  NAND2X1 U31061 ( .A(n36605), .B(n36606), .Y(n36592) );
  AOI22X1 U31062 ( .A(n26408), .B(reg_A[125]), .C(n36521), .D(n36329), .Y(
        n36606) );
  INVX1 U31063 ( .A(n36607), .Y(n36521) );
  OAI21X1 U31064 ( .A(n36608), .B(n36439), .C(n36609), .Y(n36607) );
  AOI22X1 U31065 ( .A(n36335), .B(n25428), .C(n36442), .D(n36339), .Y(n36609)
         );
  NAND2X1 U31066 ( .A(n36610), .B(n36611), .Y(n36335) );
  AOI22X1 U31067 ( .A(n36457), .B(n36612), .C(reg_B[125]), .D(n36613), .Y(
        n36611) );
  INVX1 U31068 ( .A(n36180), .Y(n36457) );
  NAND2X1 U31069 ( .A(reg_B[123]), .B(n36177), .Y(n36180) );
  AOI22X1 U31070 ( .A(n25409), .B(n25337), .C(n25427), .D(n25323), .Y(n36610)
         );
  AOI22X1 U31071 ( .A(reg_A[113]), .B(n26357), .C(reg_A[114]), .D(n26359), .Y(
        n36605) );
  INVX1 U31072 ( .A(n36614), .Y(n26357) );
  NOR2X1 U31073 ( .A(n36615), .B(n36616), .Y(n36531) );
  OAI21X1 U31074 ( .A(n26328), .B(n25332), .C(n36617), .Y(n36616) );
  AOI22X1 U31075 ( .A(n25188), .B(n36618), .C(n36619), .D(n36257), .Y(n36617)
         );
  OAI21X1 U31076 ( .A(n25332), .B(n36231), .C(n36620), .Y(n36618) );
  OAI21X1 U31077 ( .A(n36621), .B(n36622), .C(n36235), .Y(n36620) );
  OAI21X1 U31078 ( .A(n36623), .B(n25568), .C(n36624), .Y(n36622) );
  NAND2X1 U31079 ( .A(n36241), .B(n36625), .Y(n36624) );
  OAI21X1 U31080 ( .A(n25483), .B(n36246), .C(n36626), .Y(n36625) );
  INVX1 U31081 ( .A(n36303), .Y(n36623) );
  OAI21X1 U31082 ( .A(n36247), .B(n36627), .C(n36628), .Y(n36621) );
  AOI21X1 U31083 ( .A(n36629), .B(n36525), .C(n36630), .Y(n36628) );
  OAI21X1 U31084 ( .A(n25493), .B(n36312), .C(n36631), .Y(n36525) );
  AOI22X1 U31085 ( .A(n36442), .B(reg_A[122]), .C(n36315), .D(reg_A[124]), .Y(
        n36631) );
  NOR2X1 U31086 ( .A(reg_B[127]), .B(reg_B[124]), .Y(n36629) );
  NAND2X1 U31087 ( .A(n25399), .B(reg_A[118]), .Y(n36627) );
  NAND2X1 U31088 ( .A(n36632), .B(n36633), .Y(n36615) );
  AOI22X1 U31089 ( .A(reg_A[115]), .B(n26346), .C(reg_A[118]), .D(n26347), .Y(
        n36633) );
  AOI22X1 U31090 ( .A(reg_A[120]), .B(n26348), .C(n26349), .D(reg_A[109]), .Y(
        n36632) );
  NAND2X1 U31091 ( .A(n36634), .B(n36635), .Y(result[123]) );
  NOR2X1 U31092 ( .A(n36636), .B(n36637), .Y(n36635) );
  NAND3X1 U31093 ( .A(n36638), .B(n36639), .C(n36640), .Y(n36637) );
  NOR2X1 U31094 ( .A(n36641), .B(n36642), .Y(n36640) );
  INVX1 U31095 ( .A(n36643), .Y(n36642) );
  AOI22X1 U31096 ( .A(n36329), .B(n36585), .C(n36286), .D(n36630), .Y(n36643)
         );
  INVX1 U31097 ( .A(n36591), .Y(n36630) );
  NAND2X1 U31098 ( .A(n36240), .B(reg_A[112]), .Y(n36591) );
  AND2X1 U31099 ( .A(n36644), .B(n36645), .Y(n36585) );
  AOI22X1 U31100 ( .A(n36315), .B(n36178), .C(n36442), .D(n36459), .Y(n36645)
         );
  OAI21X1 U31101 ( .A(reg_A[115]), .B(n36318), .C(n36646), .Y(n36178) );
  AOI22X1 U31102 ( .A(reg_B[123]), .B(n36647), .C(n36338), .D(n25321), .Y(
        n36646) );
  INVX1 U31103 ( .A(n36648), .Y(n36647) );
  AOI22X1 U31104 ( .A(n36649), .B(n36650), .C(n36280), .D(n36651), .Y(n36644)
         );
  OAI22X1 U31105 ( .A(n25323), .B(n26136), .C(n25317), .D(n26812), .Y(n36641)
         );
  AOI22X1 U31106 ( .A(reg_A[116]), .B(n36652), .C(reg_A[123]), .D(n26450), .Y(
        n36639) );
  AOI22X1 U31107 ( .A(n26451), .B(reg_A[126]), .C(n36530), .D(n25150), .Y(
        n36638) );
  INVX1 U31108 ( .A(n36653), .Y(n36530) );
  OAI21X1 U31109 ( .A(reg_B[2]), .B(n36268), .C(n36654), .Y(n36653) );
  AOI22X1 U31110 ( .A(n26455), .B(n25476), .C(n26456), .D(n36655), .Y(n36654)
         );
  INVX1 U31111 ( .A(n36271), .Y(n36655) );
  AND2X1 U31112 ( .A(n36656), .B(n36657), .Y(n36268) );
  AOI22X1 U31113 ( .A(n26460), .B(n25335), .C(n26461), .D(n25321), .Y(n36657)
         );
  NOR2X1 U31114 ( .A(reg_B[1]), .B(reg_B[4]), .Y(n26461) );
  NOR2X1 U31115 ( .A(n26596), .B(reg_B[4]), .Y(n26460) );
  AOI22X1 U31116 ( .A(n26462), .B(n25494), .C(n26463), .D(n25771), .Y(n36656)
         );
  INVX1 U31117 ( .A(n26418), .Y(n26451) );
  NAND3X1 U31118 ( .A(n36658), .B(n36659), .C(n36660), .Y(n36636) );
  NOR2X1 U31119 ( .A(n36661), .B(n36662), .Y(n36660) );
  OAI21X1 U31120 ( .A(n26490), .B(n25490), .C(n36663), .Y(n36662) );
  OAI21X1 U31121 ( .A(n36664), .B(n36665), .C(n36666), .Y(n36663) );
  OAI21X1 U31122 ( .A(n25087), .B(n36667), .C(n25523), .Y(n36665) );
  NOR2X1 U31123 ( .A(n26996), .B(n36668), .Y(n36664) );
  NOR2X1 U31124 ( .A(n34633), .B(n36669), .Y(n26490) );
  OAI21X1 U31125 ( .A(n36670), .B(n36671), .C(n36672), .Y(n36661) );
  OAI21X1 U31126 ( .A(n36673), .B(n36674), .C(reg_A[120]), .Y(n36672) );
  OAI21X1 U31127 ( .A(n25031), .B(n36246), .C(n26473), .Y(n36674) );
  AND2X1 U31128 ( .A(n36675), .B(n36570), .Y(n36659) );
  OAI21X1 U31129 ( .A(n36298), .B(n26626), .C(reg_A[122]), .Y(n36675) );
  NOR2X1 U31130 ( .A(n36325), .B(n25568), .Y(n36298) );
  AOI22X1 U31131 ( .A(n36573), .B(n36571), .C(n26482), .D(reg_A[127]), .Y(
        n36658) );
  OAI21X1 U31132 ( .A(n36676), .B(n26999), .C(n36677), .Y(n36571) );
  INVX1 U31133 ( .A(n36678), .Y(n36677) );
  AOI21X1 U31134 ( .A(n36679), .B(n36680), .C(n25403), .Y(n36678) );
  AOI22X1 U31135 ( .A(n36681), .B(n36280), .C(n36447), .D(n36649), .Y(n36680)
         );
  AOI22X1 U31136 ( .A(n36446), .B(n36442), .C(n36143), .D(n36315), .Y(n36679)
         );
  NAND2X1 U31137 ( .A(n36682), .B(n36683), .Y(n36143) );
  AOI22X1 U31138 ( .A(n36684), .B(reg_A[99]), .C(n36685), .D(reg_A[107]), .Y(
        n36683) );
  AOI22X1 U31139 ( .A(n36338), .B(reg_A[123]), .C(n36686), .D(reg_A[115]), .Y(
        n36682) );
  INVX1 U31140 ( .A(n36687), .Y(n36573) );
  NOR2X1 U31141 ( .A(n36688), .B(n36689), .Y(n36634) );
  NAND3X1 U31142 ( .A(n36690), .B(n36691), .C(n36692), .Y(n36689) );
  NOR2X1 U31143 ( .A(n36693), .B(n36694), .Y(n36692) );
  OAI22X1 U31144 ( .A(n25469), .B(n26625), .C(n25452), .D(n26917), .Y(n36694)
         );
  MUX2X1 U31145 ( .B(n36695), .A(n36696), .S(reg_B[127]), .Y(n36693) );
  AOI21X1 U31146 ( .A(n25170), .B(n36697), .C(n36698), .Y(n36696) );
  OAI21X1 U31147 ( .A(n27438), .B(n36699), .C(n36700), .Y(n36698) );
  OR2X1 U31148 ( .A(n25031), .B(n36676), .Y(n36695) );
  AOI22X1 U31149 ( .A(reg_A[123]), .B(n36315), .C(reg_A[121]), .D(n36442), .Y(
        n36676) );
  AOI22X1 U31150 ( .A(reg_A[118]), .B(n26353), .C(reg_A[114]), .D(n26346), .Y(
        n36691) );
  AOI22X1 U31151 ( .A(reg_A[117]), .B(n26347), .C(n36701), .D(n36702), .Y(
        n36690) );
  OAI21X1 U31152 ( .A(n36587), .B(n36136), .C(n36703), .Y(n36701) );
  AOI22X1 U31153 ( .A(n25793), .B(n36303), .C(n25700), .D(n36704), .Y(n36703)
         );
  OAI21X1 U31154 ( .A(n36236), .B(n25321), .C(n36705), .Y(n36303) );
  AOI22X1 U31155 ( .A(n36241), .B(reg_A[115]), .C(n36355), .D(reg_A[119]), .Y(
        n36705) );
  INVX1 U31156 ( .A(n36706), .Y(n36587) );
  NAND3X1 U31157 ( .A(n36707), .B(n36708), .C(n36709), .Y(n36688) );
  NOR2X1 U31158 ( .A(n36710), .B(n36711), .Y(n36709) );
  OAI22X1 U31159 ( .A(n26526), .B(n25483), .C(n26534), .D(n36140), .Y(n36711)
         );
  OAI21X1 U31160 ( .A(n36614), .B(n25476), .C(n36712), .Y(n36710) );
  OAI21X1 U31161 ( .A(n36713), .B(n36714), .C(n25840), .Y(n36712) );
  NAND3X1 U31162 ( .A(n36715), .B(n36716), .C(n36717), .Y(n36714) );
  AOI21X1 U31163 ( .A(reg_A[110]), .B(n25325), .C(n36718), .Y(n36717) );
  OAI22X1 U31164 ( .A(n25035), .B(n25474), .C(n25784), .D(n25494), .Y(n36718)
         );
  AOI22X1 U31165 ( .A(n25857), .B(reg_A[98]), .C(n25647), .D(reg_A[99]), .Y(
        n36716) );
  AOI22X1 U31166 ( .A(n25648), .B(reg_A[96]), .C(n26432), .D(reg_A[97]), .Y(
        n36715) );
  NAND3X1 U31167 ( .A(n36719), .B(n36720), .C(n36721), .Y(n36713) );
  NOR2X1 U31168 ( .A(n36722), .B(n36723), .Y(n36721) );
  OAI22X1 U31169 ( .A(n25051), .B(n25296), .C(n25038), .D(n25298), .Y(n36723)
         );
  OAI22X1 U31170 ( .A(n25334), .B(n25470), .C(n25336), .D(n25468), .Y(n36722)
         );
  AOI22X1 U31171 ( .A(reg_A[101]), .B(n25242), .C(reg_A[100]), .D(n25338), .Y(
        n36720) );
  AOI22X1 U31172 ( .A(reg_A[103]), .B(n25339), .C(reg_A[102]), .D(n25257), .Y(
        n36719) );
  AOI22X1 U31173 ( .A(n36596), .B(n26028), .C(n36724), .D(n26260), .Y(n36708)
         );
  INVX1 U31174 ( .A(n36725), .Y(n36724) );
  AND2X1 U31175 ( .A(n36726), .B(n36727), .Y(n36596) );
  AOI22X1 U31176 ( .A(n25025), .B(n36728), .C(n25026), .D(n36464), .Y(n36727)
         );
  AOI22X1 U31177 ( .A(n26032), .B(n36269), .C(n26530), .D(n36729), .Y(n36726)
         );
  OAI21X1 U31178 ( .A(reg_A[123]), .B(n25063), .C(n36730), .Y(n36269) );
  AOI22X1 U31179 ( .A(n26038), .B(n25335), .C(reg_B[0]), .D(n36731), .Y(n36730) );
  AOI22X1 U31180 ( .A(n36732), .B(n26262), .C(reg_A[115]), .D(n26551), .Y(
        n36707) );
  INVX1 U31181 ( .A(n36733), .Y(n36732) );
  NAND2X1 U31182 ( .A(n36734), .B(n36735), .Y(result[122]) );
  NOR2X1 U31183 ( .A(n36736), .B(n36737), .Y(n36735) );
  NAND3X1 U31184 ( .A(n36738), .B(n36739), .C(n36740), .Y(n36737) );
  AND2X1 U31185 ( .A(n36741), .B(n36742), .Y(n36740) );
  AOI22X1 U31186 ( .A(n36652), .B(reg_A[115]), .C(n36256), .D(n36296), .Y(
        n36742) );
  INVX1 U31187 ( .A(n36743), .Y(n36296) );
  NAND2X1 U31188 ( .A(n26328), .B(n36434), .Y(n36652) );
  INVX1 U31189 ( .A(n36297), .Y(n36434) );
  INVX1 U31190 ( .A(n34282), .Y(n26328) );
  AOI21X1 U31191 ( .A(n36362), .B(n36744), .C(n36745), .Y(n36741) );
  OAI22X1 U31192 ( .A(n36746), .B(n36747), .C(n36136), .D(n36748), .Y(n36745)
         );
  AOI22X1 U31193 ( .A(reg_A[119]), .B(n36673), .C(reg_A[112]), .D(n26572), .Y(
        n36739) );
  NAND2X1 U31194 ( .A(n26526), .B(n30827), .Y(n26572) );
  INVX1 U31195 ( .A(n26359), .Y(n26526) );
  OAI21X1 U31196 ( .A(n25036), .B(n30951), .C(n28512), .Y(n26359) );
  NAND2X1 U31197 ( .A(n26634), .B(n36260), .Y(n36673) );
  INVX1 U31198 ( .A(n26472), .Y(n26634) );
  OAI21X1 U31199 ( .A(n25041), .B(n30951), .C(n28715), .Y(n26472) );
  AOI22X1 U31200 ( .A(n25700), .B(n36749), .C(reg_A[122]), .D(n26450), .Y(
        n36738) );
  NAND2X1 U31201 ( .A(n36584), .B(n36750), .Y(n26450) );
  INVX1 U31202 ( .A(n36751), .Y(n36584) );
  OAI21X1 U31203 ( .A(n25043), .B(n30951), .C(n36752), .Y(n36751) );
  AND2X1 U31204 ( .A(n30282), .B(n32827), .Y(n36752) );
  NAND3X1 U31205 ( .A(n36753), .B(n36754), .C(n36755), .Y(n36736) );
  NOR2X1 U31206 ( .A(n36756), .B(n36757), .Y(n36755) );
  OAI22X1 U31207 ( .A(n36557), .B(n36415), .C(n26584), .D(n36305), .Y(n36757)
         );
  NAND2X1 U31208 ( .A(n36758), .B(n36759), .Y(n36305) );
  AOI22X1 U31209 ( .A(n26593), .B(n25771), .C(n26594), .D(n25476), .Y(n36759)
         );
  INVX1 U31210 ( .A(n28739), .Y(n26594) );
  NOR2X1 U31211 ( .A(n26599), .B(n26596), .Y(n26593) );
  AOI22X1 U31212 ( .A(n36760), .B(n26596), .C(n26597), .D(n36761), .Y(n36758)
         );
  OAI21X1 U31213 ( .A(reg_A[122]), .B(n26599), .C(n36762), .Y(n36760) );
  AOI22X1 U31214 ( .A(n26601), .B(n25493), .C(n26602), .D(n36140), .Y(n36762)
         );
  INVX1 U31215 ( .A(n36704), .Y(n36557) );
  OAI21X1 U31216 ( .A(n36236), .B(n25494), .C(n36763), .Y(n36704) );
  AOI22X1 U31217 ( .A(n36241), .B(reg_A[114]), .C(n36355), .D(reg_A[118]), .Y(
        n36763) );
  OAI21X1 U31218 ( .A(n36764), .B(n36687), .C(n36765), .Y(n36756) );
  AOI21X1 U31219 ( .A(reg_A[120]), .B(n36766), .C(n36767), .Y(n36765) );
  INVX1 U31220 ( .A(n36700), .Y(n36767) );
  OAI21X1 U31221 ( .A(n36315), .B(n25342), .C(n26573), .Y(n36766) );
  NOR2X1 U31222 ( .A(n34633), .B(n36768), .Y(n26573) );
  OAI21X1 U31223 ( .A(n25040), .B(n30951), .C(n32817), .Y(n34633) );
  NAND2X1 U31224 ( .A(n25170), .B(n36172), .Y(n36687) );
  INVX1 U31225 ( .A(n36697), .Y(n36764) );
  OAI21X1 U31226 ( .A(n36769), .B(n26999), .C(n36770), .Y(n36697) );
  OAI21X1 U31227 ( .A(n36771), .B(n36772), .C(n25044), .Y(n36770) );
  INVX1 U31228 ( .A(n36773), .Y(n36772) );
  AOI22X1 U31229 ( .A(n36774), .B(n36280), .C(n36582), .D(n36649), .Y(n36773)
         );
  OAI22X1 U31230 ( .A(n36775), .B(n36360), .C(n36311), .D(n36359), .Y(n36771)
         );
  AND2X1 U31231 ( .A(n36776), .B(n36777), .Y(n36311) );
  AOI22X1 U31232 ( .A(n36338), .B(reg_A[122]), .C(n36686), .D(reg_A[114]), .Y(
        n36777) );
  AOI22X1 U31233 ( .A(n36685), .B(reg_A[106]), .C(n36684), .D(reg_A[98]), .Y(
        n36776) );
  INVX1 U31234 ( .A(n36581), .Y(n36775) );
  AOI22X1 U31235 ( .A(n36442), .B(reg_A[120]), .C(n36315), .D(reg_A[122]), .Y(
        n36769) );
  AOI22X1 U31236 ( .A(n36778), .B(n36779), .C(n30865), .D(reg_A[127]), .Y(
        n36754) );
  INVX1 U31237 ( .A(n26581), .Y(n30865) );
  NAND2X1 U31238 ( .A(n25203), .B(n34599), .Y(n26581) );
  AOI22X1 U31239 ( .A(n26482), .B(reg_A[126]), .C(n36302), .D(n36780), .Y(
        n36753) );
  NOR2X1 U31240 ( .A(n30931), .B(n26895), .Y(n26482) );
  NOR2X1 U31241 ( .A(n36781), .B(n36782), .Y(n36734) );
  NAND3X1 U31242 ( .A(n36783), .B(n36784), .C(n36785), .Y(n36782) );
  NOR2X1 U31243 ( .A(n36786), .B(n36787), .Y(n36785) );
  OAI22X1 U31244 ( .A(n26483), .B(n25490), .C(n34625), .D(n25337), .Y(n36787)
         );
  INVX1 U31245 ( .A(n26347), .Y(n34625) );
  OAI21X1 U31246 ( .A(n25033), .B(n30951), .C(n28714), .Y(n26347) );
  OAI21X1 U31247 ( .A(n26633), .B(n25483), .C(n36788), .Y(n36786) );
  AOI22X1 U31248 ( .A(reg_A[114]), .B(n26551), .C(reg_A[117]), .D(n26353), .Y(
        n36788) );
  OAI21X1 U31249 ( .A(n25028), .B(n30951), .C(n28571), .Y(n26353) );
  OAI21X1 U31250 ( .A(n25034), .B(n30951), .C(n25178), .Y(n26551) );
  INVX1 U31251 ( .A(n26346), .Y(n26633) );
  OAI21X1 U31252 ( .A(n25037), .B(n30951), .C(n36789), .Y(n26346) );
  AOI22X1 U31253 ( .A(n26627), .B(reg_A[111]), .C(n26519), .D(reg_A[110]), .Y(
        n36784) );
  INVX1 U31254 ( .A(n26917), .Y(n26519) );
  AOI22X1 U31255 ( .A(n26349), .B(reg_A[107]), .C(n36790), .D(n36257), .Y(
        n36783) );
  NAND3X1 U31256 ( .A(n36791), .B(n36792), .C(n36793), .Y(n36781) );
  NOR2X1 U31257 ( .A(n36794), .B(n36795), .Y(n36793) );
  OAI22X1 U31258 ( .A(n26012), .B(n36796), .C(n26525), .D(n36725), .Y(n36795)
         );
  NAND2X1 U31259 ( .A(n36797), .B(n36798), .Y(n36725) );
  AOI22X1 U31260 ( .A(n25025), .B(n36799), .C(n25026), .D(n36602), .Y(n36798)
         );
  AOI22X1 U31261 ( .A(n26032), .B(n36405), .C(n26530), .D(n36800), .Y(n36797)
         );
  NAND2X1 U31262 ( .A(n36801), .B(n36802), .Y(n36405) );
  AOI22X1 U31263 ( .A(n26662), .B(n25289), .C(n26663), .D(n25468), .Y(n36802)
         );
  AOI22X1 U31264 ( .A(n26038), .B(n25771), .C(n26664), .D(n25494), .Y(n36801)
         );
  OAI21X1 U31265 ( .A(n26534), .B(n25333), .C(n36803), .Y(n36794) );
  OAI21X1 U31266 ( .A(n36804), .B(n36805), .C(n25840), .Y(n36803) );
  NAND3X1 U31267 ( .A(n36806), .B(n36807), .C(n36808), .Y(n36805) );
  AOI21X1 U31268 ( .A(reg_A[109]), .B(n25325), .C(n36809), .Y(n36808) );
  OAI22X1 U31269 ( .A(n25035), .B(n25469), .C(n25042), .D(n25490), .Y(n36809)
         );
  AOI22X1 U31270 ( .A(reg_A[101]), .B(n25257), .C(n25857), .D(reg_A[97]), .Y(
        n36807) );
  AOI22X1 U31271 ( .A(n25647), .B(reg_A[98]), .C(n26432), .D(reg_A[96]), .Y(
        n36806) );
  INVX1 U31272 ( .A(n25316), .Y(n26432) );
  NAND3X1 U31273 ( .A(n36810), .B(n36811), .C(n36812), .Y(n36804) );
  AOI21X1 U31274 ( .A(reg_A[102]), .B(n25339), .C(n36813), .Y(n36812) );
  OAI22X1 U31275 ( .A(n25396), .B(n25491), .C(n25492), .D(n25436), .Y(n36813)
         );
  AOI22X1 U31276 ( .A(reg_A[105]), .B(n25246), .C(reg_A[106]), .D(n25247), .Y(
        n36811) );
  AOI22X1 U31277 ( .A(reg_A[103]), .B(n25487), .C(reg_A[104]), .D(n25241), .Y(
        n36810) );
  INVX1 U31278 ( .A(n26636), .Y(n26534) );
  OAI21X1 U31279 ( .A(n25056), .B(n30951), .C(n28679), .Y(n26636) );
  AOI21X1 U31280 ( .A(n26310), .B(reg_A[124]), .C(n36814), .Y(n36792) );
  OAI22X1 U31281 ( .A(n25317), .B(n26418), .C(n26420), .D(n36345), .Y(n36814)
         );
  INVX1 U31282 ( .A(n26812), .Y(n26310) );
  AOI22X1 U31283 ( .A(n26408), .B(reg_A[123]), .C(n36815), .D(n36329), .Y(
        n36791) );
  INVX1 U31284 ( .A(n36699), .Y(n36815) );
  NAND2X1 U31285 ( .A(n36816), .B(n36817), .Y(n36699) );
  AOI22X1 U31286 ( .A(n36315), .B(n36339), .C(n36442), .D(n36613), .Y(n36817)
         );
  NAND2X1 U31287 ( .A(n36818), .B(n36819), .Y(n36339) );
  AOI22X1 U31288 ( .A(n36684), .B(n25289), .C(n36685), .D(n25468), .Y(n36819)
         );
  AOI22X1 U31289 ( .A(n36338), .B(n25494), .C(n36686), .D(n25771), .Y(n36818)
         );
  AOI22X1 U31290 ( .A(n36649), .B(n36820), .C(n36280), .D(n36821), .Y(n36816)
         );
  INVX1 U31291 ( .A(n26136), .Y(n26408) );
  NAND3X1 U31292 ( .A(n36822), .B(n36823), .C(n36824), .Y(result[121]) );
  NOR2X1 U31293 ( .A(n36825), .B(n36826), .Y(n36824) );
  NAND3X1 U31294 ( .A(n36827), .B(n36828), .C(n36829), .Y(n36826) );
  NOR2X1 U31295 ( .A(n36830), .B(n36831), .Y(n36829) );
  OAI22X1 U31296 ( .A(n26012), .B(n36832), .C(n26525), .D(n36796), .Y(n36831)
         );
  NAND2X1 U31297 ( .A(n36833), .B(n36834), .Y(n36796) );
  AOI22X1 U31298 ( .A(n25025), .B(n36729), .C(n25026), .D(n36728), .Y(n36834)
         );
  AOI22X1 U31299 ( .A(n26032), .B(n36464), .C(n26530), .D(n36835), .Y(n36833)
         );
  NAND2X1 U31300 ( .A(n36836), .B(n36837), .Y(n36464) );
  AOI22X1 U31301 ( .A(n26662), .B(n25287), .C(n26663), .D(n25296), .Y(n36837)
         );
  INVX1 U31302 ( .A(n26982), .Y(n26663) );
  AOI22X1 U31303 ( .A(n26038), .B(n25483), .C(n26664), .D(n25490), .Y(n36836)
         );
  OAI21X1 U31304 ( .A(n36838), .B(n36746), .C(n36839), .Y(n36830) );
  OAI21X1 U31305 ( .A(n36840), .B(n36841), .C(n25840), .Y(n36839) );
  NAND2X1 U31306 ( .A(n36842), .B(n36843), .Y(n36841) );
  NOR2X1 U31307 ( .A(n36844), .B(n36845), .Y(n36843) );
  OAI21X1 U31308 ( .A(n25034), .B(n25483), .C(n36846), .Y(n36845) );
  AOI22X1 U31309 ( .A(reg_A[116]), .B(n25123), .C(reg_A[112]), .D(n25629), .Y(
        n36846) );
  OAI21X1 U31310 ( .A(n25056), .B(n25332), .C(n36847), .Y(n36844) );
  AOI22X1 U31311 ( .A(reg_A[115]), .B(n25253), .C(reg_A[114]), .D(n25628), .Y(
        n36847) );
  NOR2X1 U31312 ( .A(n36848), .B(n36849), .Y(n36842) );
  OAI21X1 U31313 ( .A(n25043), .B(n25490), .C(n36850), .Y(n36849) );
  AOI22X1 U31314 ( .A(reg_A[109]), .B(n25635), .C(reg_A[108]), .D(n25325), .Y(
        n36850) );
  OAI21X1 U31315 ( .A(n25035), .B(n25470), .C(n36851), .Y(n36848) );
  AOI22X1 U31316 ( .A(reg_A[110]), .B(n25222), .C(reg_A[111]), .D(n25637), .Y(
        n36851) );
  NAND3X1 U31317 ( .A(n36852), .B(n36853), .C(n36854), .Y(n36840) );
  NOR2X1 U31318 ( .A(n36855), .B(n36856), .Y(n36854) );
  OAI21X1 U31319 ( .A(n25040), .B(n36140), .C(n36857), .Y(n36856) );
  AOI22X1 U31320 ( .A(reg_A[120]), .B(n25135), .C(reg_A[118]), .D(n25136), .Y(
        n36857) );
  OAI21X1 U31321 ( .A(n25287), .B(n25320), .C(n36858), .Y(n36855) );
  AOI22X1 U31322 ( .A(reg_A[100]), .B(n25257), .C(n25857), .D(reg_A[96]), .Y(
        n36858) );
  NOR2X1 U31323 ( .A(n36859), .B(n36860), .Y(n36853) );
  OAI22X1 U31324 ( .A(n25051), .B(n25448), .C(n25038), .D(n25361), .Y(n36860)
         );
  OAI22X1 U31325 ( .A(n25334), .B(n25296), .C(n25336), .D(n25298), .Y(n36859)
         );
  AOI21X1 U31326 ( .A(reg_A[101]), .B(n25339), .C(n36861), .Y(n36852) );
  OAI22X1 U31327 ( .A(n25289), .B(n25491), .C(n25492), .D(n25396), .Y(n36861)
         );
  NAND2X1 U31328 ( .A(n36862), .B(n36863), .Y(n36746) );
  AOI22X1 U31329 ( .A(n36315), .B(n36459), .C(n36442), .D(n36650), .Y(n36863)
         );
  INVX1 U31330 ( .A(n36453), .Y(n36650) );
  NAND2X1 U31331 ( .A(n36864), .B(n36865), .Y(n36459) );
  AOI22X1 U31332 ( .A(n36684), .B(n25287), .C(n36685), .D(n25296), .Y(n36865)
         );
  AOI22X1 U31333 ( .A(n36338), .B(n25490), .C(n36686), .D(n25483), .Y(n36864)
         );
  AOI22X1 U31334 ( .A(n36649), .B(n36651), .C(n36280), .D(n36866), .Y(n36862)
         );
  INVX1 U31335 ( .A(n36867), .Y(n36866) );
  OAI21X1 U31336 ( .A(n36868), .B(n36869), .C(n25918), .Y(n36828) );
  OR2X1 U31337 ( .A(n36870), .B(n36871), .Y(n36869) );
  OAI21X1 U31338 ( .A(n25736), .B(n25490), .C(n36872), .Y(n36871) );
  INVX1 U31339 ( .A(n36873), .Y(n36872) );
  OAI22X1 U31340 ( .A(n27252), .B(n25483), .C(n27253), .D(n25476), .Y(n36870)
         );
  OR2X1 U31341 ( .A(n36874), .B(n36875), .Y(n36868) );
  OAI22X1 U31342 ( .A(n26800), .B(n25337), .C(n26801), .D(n25332), .Y(n36875)
         );
  OAI21X1 U31343 ( .A(n25062), .B(n36140), .C(n36876), .Y(n36874) );
  AOI22X1 U31344 ( .A(reg_A[120]), .B(n26803), .C(reg_A[118]), .D(n26804), .Y(
        n36876) );
  AOI22X1 U31345 ( .A(n26349), .B(reg_A[106]), .C(n36877), .D(n36257), .Y(
        n36827) );
  INVX1 U31346 ( .A(n26625), .Y(n26349) );
  NAND3X1 U31347 ( .A(n36878), .B(n36879), .C(n36880), .Y(n36825) );
  NOR2X1 U31348 ( .A(n36881), .B(n36882), .Y(n36880) );
  OAI22X1 U31349 ( .A(n25494), .B(n26136), .C(n25321), .D(n26812), .Y(n36882)
         );
  NAND2X1 U31350 ( .A(n25203), .B(n29569), .Y(n26812) );
  NAND2X1 U31351 ( .A(n25203), .B(n29568), .Y(n26136) );
  OAI22X1 U31352 ( .A(n26854), .B(n36733), .C(n25323), .D(n26418), .Y(n36881)
         );
  NAND2X1 U31353 ( .A(n25203), .B(n36883), .Y(n26418) );
  NAND2X1 U31354 ( .A(n36884), .B(n36885), .Y(n36733) );
  AOI22X1 U31355 ( .A(n26859), .B(n25337), .C(n26860), .D(n25332), .Y(n36885)
         );
  AOI22X1 U31356 ( .A(n26455), .B(n25476), .C(n36472), .D(n26452), .Y(n36884)
         );
  OAI21X1 U31357 ( .A(reg_A[112]), .B(n26861), .C(n36886), .Y(n36472) );
  AOI22X1 U31358 ( .A(n36761), .B(n26863), .C(n26462), .D(n25493), .Y(n36886)
         );
  MUX2X1 U31359 ( .B(reg_A[113]), .A(reg_A[121]), .S(n26596), .Y(n36761) );
  AOI22X1 U31360 ( .A(n30910), .B(n36873), .C(n36252), .D(reg_B[127]), .Y(
        n36879) );
  INVX1 U31361 ( .A(n36887), .Y(n36252) );
  OAI22X1 U31362 ( .A(n26936), .B(n25771), .C(n25745), .D(n25335), .Y(n36873)
         );
  AOI22X1 U31363 ( .A(n25793), .B(n36749), .C(n25700), .D(n36888), .Y(n36878)
         );
  OAI21X1 U31364 ( .A(n36889), .B(n25490), .C(n36890), .Y(n36749) );
  OAI21X1 U31365 ( .A(n26267), .B(n36286), .C(n36706), .Y(n36890) );
  OAI21X1 U31366 ( .A(n36236), .B(n25490), .C(n36891), .Y(n36706) );
  AOI22X1 U31367 ( .A(n36241), .B(reg_A[113]), .C(n36355), .D(reg_A[117]), .Y(
        n36891) );
  AOI21X1 U31368 ( .A(n26186), .B(n36177), .C(n36256), .Y(n36889) );
  INVX1 U31369 ( .A(n36325), .Y(n36256) );
  NAND2X1 U31370 ( .A(n26504), .B(n36177), .Y(n36325) );
  NOR2X1 U31371 ( .A(n36892), .B(n36893), .Y(n36823) );
  NAND2X1 U31372 ( .A(n36894), .B(n36895), .Y(n36893) );
  AOI22X1 U31373 ( .A(n36778), .B(n36896), .C(n36436), .D(n36779), .Y(n36895)
         );
  NAND2X1 U31374 ( .A(n36897), .B(n36898), .Y(n36779) );
  AOI22X1 U31375 ( .A(n36315), .B(n36446), .C(n36442), .D(n36447), .Y(n36898)
         );
  NAND2X1 U31376 ( .A(n36899), .B(n36900), .Y(n36446) );
  AOI22X1 U31377 ( .A(n36684), .B(reg_A[97]), .C(n36685), .D(reg_A[105]), .Y(
        n36900) );
  AOI22X1 U31378 ( .A(n36338), .B(reg_A[121]), .C(n36686), .D(reg_A[113]), .Y(
        n36899) );
  AOI22X1 U31379 ( .A(n36649), .B(n36681), .C(n36280), .D(n36901), .Y(n36897)
         );
  AOI22X1 U31380 ( .A(n36271), .B(n25166), .C(n36302), .D(n36902), .Y(n36894)
         );
  INVX1 U31381 ( .A(n26881), .Y(n25166) );
  NAND3X1 U31382 ( .A(n36700), .B(n36570), .C(n36903), .Y(n36892) );
  AOI22X1 U31383 ( .A(reg_A[120]), .B(n36904), .C(n36417), .D(n36780), .Y(
        n36903) );
  INVX1 U31384 ( .A(n36905), .Y(n36417) );
  OAI21X1 U31385 ( .A(n25793), .B(n25342), .C(n26791), .Y(n36904) );
  INVX1 U31386 ( .A(n34606), .Y(n26791) );
  NAND2X1 U31387 ( .A(n36263), .B(reg_A[120]), .Y(n36570) );
  NOR2X1 U31388 ( .A(n36177), .B(n25031), .Y(n36263) );
  NAND3X1 U31389 ( .A(reg_B[124]), .B(n25188), .C(n36906), .Y(n36700) );
  NOR2X1 U31390 ( .A(n36907), .B(n36908), .Y(n36822) );
  OAI21X1 U31391 ( .A(n36909), .B(n25490), .C(n36910), .Y(n36908) );
  AOI22X1 U31392 ( .A(n36744), .B(n36911), .C(n26866), .D(reg_A[112]), .Y(
        n36910) );
  INVX1 U31393 ( .A(n30913), .Y(n26866) );
  INVX1 U31394 ( .A(n26883), .Y(n36909) );
  NAND2X1 U31395 ( .A(n36750), .B(n30282), .Y(n26883) );
  NAND2X1 U31396 ( .A(n25203), .B(n25284), .Y(n30282) );
  NAND2X1 U31397 ( .A(n36912), .B(n36913), .Y(n36907) );
  AOI22X1 U31398 ( .A(n36914), .B(n36294), .C(n36297), .D(reg_A[114]), .Y(
        n36913) );
  INVX1 U31399 ( .A(n36915), .Y(n36914) );
  AOI22X1 U31400 ( .A(n36916), .B(reg_A[118]), .C(n25203), .D(n36917), .Y(
        n36912) );
  OAI21X1 U31401 ( .A(n26895), .B(n25317), .C(n36918), .Y(n36917) );
  AOI22X1 U31402 ( .A(reg_A[127]), .B(n34598), .C(reg_A[126]), .D(n34599), .Y(
        n36918) );
  NAND2X1 U31403 ( .A(n36919), .B(n36920), .Y(result[120]) );
  NOR2X1 U31404 ( .A(n36921), .B(n36922), .Y(n36920) );
  NAND3X1 U31405 ( .A(n36923), .B(n36924), .C(n36925), .Y(n36922) );
  NOR2X1 U31406 ( .A(n36926), .B(n36927), .Y(n36925) );
  OAI21X1 U31407 ( .A(n26525), .B(n36832), .C(n36928), .Y(n36927) );
  OAI21X1 U31408 ( .A(n36929), .B(n36930), .C(n25840), .Y(n36928) );
  NAND3X1 U31409 ( .A(n36931), .B(n36932), .C(n36933), .Y(n36930) );
  NOR2X1 U31410 ( .A(n36934), .B(n36935), .Y(n36933) );
  OAI21X1 U31411 ( .A(n25037), .B(n25452), .C(n36936), .Y(n36935) );
  AOI22X1 U31412 ( .A(reg_A[116]), .B(n25073), .C(reg_A[115]), .D(n25123), .Y(
        n36936) );
  OAI21X1 U31413 ( .A(n25030), .B(n25483), .C(n36937), .Y(n36934) );
  AOI22X1 U31414 ( .A(reg_A[118]), .B(n25252), .C(reg_A[114]), .D(n25253), .Y(
        n36937) );
  AOI21X1 U31415 ( .A(reg_A[106]), .B(n25234), .C(n36938), .Y(n36932) );
  OAI22X1 U31416 ( .A(n25036), .B(n25450), .C(n25467), .D(n25476), .Y(n36938)
         );
  AOI22X1 U31417 ( .A(reg_A[107]), .B(n25325), .C(reg_A[120]), .D(n25125), .Y(
        n36931) );
  NAND3X1 U31418 ( .A(n36939), .B(n36940), .C(n36941), .Y(n36929) );
  NOR2X1 U31419 ( .A(n36942), .B(n36943), .Y(n36941) );
  OAI21X1 U31420 ( .A(n25287), .B(n25491), .C(n36944), .Y(n36943) );
  AOI22X1 U31421 ( .A(reg_A[102]), .B(n25241), .C(reg_A[98]), .D(n25242), .Y(
        n36944) );
  OAI21X1 U31422 ( .A(n25038), .B(n25670), .C(n36945), .Y(n36942) );
  AOI22X1 U31423 ( .A(reg_A[103]), .B(n25246), .C(reg_A[104]), .D(n25247), .Y(
        n36945) );
  AOI21X1 U31424 ( .A(n25647), .B(reg_A[96]), .C(n36946), .Y(n36940) );
  OAI22X1 U31425 ( .A(n26719), .B(n25396), .C(n25238), .D(n25436), .Y(n36946)
         );
  AOI22X1 U31426 ( .A(reg_A[119]), .B(n25135), .C(reg_A[117]), .D(n25136), .Y(
        n36939) );
  NAND2X1 U31427 ( .A(n36947), .B(n36948), .Y(n36832) );
  AOI22X1 U31428 ( .A(n25025), .B(n36800), .C(n25026), .D(n36799), .Y(n36948)
         );
  AOI22X1 U31429 ( .A(n26032), .B(n36602), .C(n26530), .D(n36949), .Y(n36947)
         );
  OR2X1 U31430 ( .A(n36950), .B(n36951), .Y(n36602) );
  OAI22X1 U31431 ( .A(reg_A[120]), .B(n25063), .C(reg_A[112]), .D(n26981), .Y(
        n36951) );
  OAI21X1 U31432 ( .A(reg_A[104]), .B(n26982), .C(n36952), .Y(n36950) );
  OAI22X1 U31433 ( .A(n29036), .B(n25490), .C(n36838), .D(n36915), .Y(n36926)
         );
  NAND2X1 U31434 ( .A(n36953), .B(n36954), .Y(n36915) );
  AOI22X1 U31435 ( .A(n36315), .B(n36613), .C(n36442), .D(n36820), .Y(n36954)
         );
  OR2X1 U31436 ( .A(n36955), .B(n36956), .Y(n36613) );
  OAI22X1 U31437 ( .A(reg_A[112]), .B(n36318), .C(reg_A[120]), .D(n36668), .Y(
        n36956) );
  OAI21X1 U31438 ( .A(reg_A[104]), .B(n36957), .C(n36958), .Y(n36955) );
  AOI22X1 U31439 ( .A(n36649), .B(n36821), .C(n36280), .D(n36959), .Y(n36953)
         );
  AOI22X1 U31440 ( .A(n36916), .B(reg_A[117]), .C(n36744), .D(n36619), .Y(
        n36924) );
  OAI21X1 U31441 ( .A(n25087), .B(n36132), .C(n36960), .Y(n36744) );
  OAI21X1 U31442 ( .A(n25589), .B(n36961), .C(reg_B[125]), .Y(n36132) );
  AOI22X1 U31443 ( .A(n25793), .B(n36888), .C(n36559), .D(n28575), .Y(n36923)
         );
  INVX1 U31444 ( .A(n36962), .Y(n36559) );
  OAI21X1 U31445 ( .A(n25493), .B(n36963), .C(n36748), .Y(n36888) );
  AOI22X1 U31446 ( .A(n36964), .B(n26267), .C(n36965), .D(n36286), .Y(n36748)
         );
  INVX1 U31447 ( .A(n36670), .Y(n36964) );
  AOI21X1 U31448 ( .A(reg_A[112]), .B(n36241), .C(n36965), .Y(n36670) );
  OAI22X1 U31449 ( .A(n36236), .B(n25493), .C(n25337), .D(n36247), .Y(n36965)
         );
  NAND2X1 U31450 ( .A(n26186), .B(n36177), .Y(n36963) );
  NAND3X1 U31451 ( .A(n36966), .B(n36967), .C(n36968), .Y(n36921) );
  NOR2X1 U31452 ( .A(n36969), .B(n36970), .Y(n36968) );
  OAI21X1 U31453 ( .A(n36971), .B(n36905), .C(n36972), .Y(n36970) );
  OAI21X1 U31454 ( .A(n36973), .B(n27032), .C(reg_A[120]), .Y(n36972) );
  OAI21X1 U31455 ( .A(n25043), .B(n26990), .C(n32826), .Y(n27032) );
  NAND2X1 U31456 ( .A(n25399), .B(n36702), .Y(n36905) );
  OAI21X1 U31457 ( .A(n25568), .B(n36974), .C(n36887), .Y(n36969) );
  NAND2X1 U31458 ( .A(n36702), .B(n36780), .Y(n36974) );
  AOI22X1 U31459 ( .A(n36302), .B(n36975), .C(n36976), .D(n36294), .Y(n36967)
         );
  INVX1 U31460 ( .A(n36671), .Y(n36302) );
  NAND2X1 U31461 ( .A(n25355), .B(n26267), .Y(n36671) );
  AOI22X1 U31462 ( .A(n36560), .B(n27008), .C(n36297), .D(reg_A[113]), .Y(
        n36966) );
  AND2X1 U31463 ( .A(n36977), .B(n36978), .Y(n36560) );
  AOI22X1 U31464 ( .A(n26601), .B(n25333), .C(n26602), .D(n25332), .Y(n36978)
         );
  AOI22X1 U31465 ( .A(n27012), .B(n25493), .C(n26597), .D(n36140), .Y(n36977)
         );
  NOR2X1 U31466 ( .A(n36979), .B(n36980), .Y(n36919) );
  NAND3X1 U31467 ( .A(n36981), .B(n36982), .C(n36983), .Y(n36980) );
  NOR2X1 U31468 ( .A(n36984), .B(n36985), .Y(n36983) );
  OAI22X1 U31469 ( .A(n36478), .B(n36986), .C(n25296), .D(n26625), .Y(n36985)
         );
  INVX1 U31470 ( .A(n36257), .Y(n36478) );
  OAI21X1 U31471 ( .A(n25087), .B(n36149), .C(n36987), .Y(n36257) );
  OAI21X1 U31472 ( .A(n36961), .B(n25589), .C(n36177), .Y(n36149) );
  OAI22X1 U31473 ( .A(n25469), .B(n26917), .C(n25474), .D(n31000), .Y(n36984)
         );
  AOI22X1 U31474 ( .A(n26928), .B(n36988), .C(n25918), .D(n36989), .Y(n36982)
         );
  NAND3X1 U31475 ( .A(n36990), .B(n36991), .C(n36992), .Y(n36989) );
  NOR2X1 U31476 ( .A(n36993), .B(n36994), .Y(n36992) );
  OAI22X1 U31477 ( .A(n26936), .B(n25483), .C(n25745), .D(n25771), .Y(n36994)
         );
  OAI21X1 U31478 ( .A(n25062), .B(n25333), .C(n36995), .Y(n36993) );
  AOI22X1 U31479 ( .A(reg_A[119]), .B(n26803), .C(reg_A[117]), .D(n26804), .Y(
        n36995) );
  AOI22X1 U31480 ( .A(reg_A[116]), .B(n25749), .C(reg_A[115]), .D(n25750), .Y(
        n36991) );
  AOI22X1 U31481 ( .A(reg_A[112]), .B(n25615), .C(reg_A[120]), .D(n26924), .Y(
        n36990) );
  NAND3X1 U31482 ( .A(n36996), .B(n36997), .C(n36998), .Y(n36988) );
  NOR2X1 U31483 ( .A(n36999), .B(n37000), .Y(n36998) );
  OAI22X1 U31484 ( .A(n26943), .B(n25493), .C(n26944), .D(n25317), .Y(n37000)
         );
  OAI22X1 U31485 ( .A(n26945), .B(n25323), .C(n25753), .D(n25497), .Y(n36999)
         );
  AOI22X1 U31486 ( .A(reg_A[121]), .B(n26007), .C(reg_A[123]), .D(n26008), .Y(
        n36997) );
  AOI22X1 U31487 ( .A(reg_A[122]), .B(n26009), .C(reg_A[126]), .D(n26010), .Y(
        n36996) );
  AOI22X1 U31488 ( .A(n25277), .B(n36896), .C(n25275), .D(n37001), .Y(n36981)
         );
  NAND2X1 U31489 ( .A(n37002), .B(n37003), .Y(n36896) );
  AOI22X1 U31490 ( .A(n36315), .B(n36581), .C(n36442), .D(n36582), .Y(n37003)
         );
  NAND2X1 U31491 ( .A(n37004), .B(n37005), .Y(n36581) );
  AOI22X1 U31492 ( .A(n36685), .B(reg_A[104]), .C(n37006), .D(reg_B[124]), .Y(
        n37005) );
  AOI22X1 U31493 ( .A(n36338), .B(reg_A[120]), .C(n36686), .D(reg_A[112]), .Y(
        n37004) );
  AOI22X1 U31494 ( .A(n36649), .B(n36774), .C(n36280), .D(n37007), .Y(n37002)
         );
  NAND3X1 U31495 ( .A(n37008), .B(n37009), .C(n37010), .Y(n36979) );
  NOR2X1 U31496 ( .A(n37011), .B(n37012), .Y(n37010) );
  OAI22X1 U31497 ( .A(n27971), .B(n25497), .C(n25295), .D(n25319), .Y(n37012)
         );
  OAI22X1 U31498 ( .A(n25297), .B(n25317), .C(n27511), .D(n25323), .Y(n37011)
         );
  AOI22X1 U31499 ( .A(n37013), .B(n26260), .C(reg_A[112]), .D(n37014), .Y(
        n37009) );
  AOI22X1 U31500 ( .A(reg_A[122]), .B(n37015), .C(reg_A[123]), .D(n29051), .Y(
        n37008) );
  NAND2X1 U31501 ( .A(n37016), .B(n37017), .Y(result[11]) );
  NOR2X1 U31502 ( .A(n37018), .B(n37019), .Y(n37017) );
  NAND3X1 U31503 ( .A(n37020), .B(n37021), .C(n37022), .Y(n37019) );
  NOR2X1 U31504 ( .A(n37023), .B(n37024), .Y(n37022) );
  OAI21X1 U31505 ( .A(n28586), .B(n25146), .C(n37025), .Y(n37024) );
  OAI21X1 U31506 ( .A(n37026), .B(n37027), .C(n26267), .Y(n37025) );
  OAI22X1 U31507 ( .A(n37028), .B(n25189), .C(n36002), .D(n26692), .Y(n37027)
         );
  INVX1 U31508 ( .A(n36058), .Y(n36002) );
  OAI21X1 U31509 ( .A(n29304), .B(n27967), .C(n37029), .Y(n36058) );
  AOI22X1 U31510 ( .A(n35865), .B(reg_A[3]), .C(reg_A[7]), .D(n26691), .Y(
        n37029) );
  NOR2X1 U31511 ( .A(n26721), .B(n25194), .Y(n37026) );
  INVX1 U31512 ( .A(n37030), .Y(n26721) );
  OAI21X1 U31513 ( .A(n32522), .B(n26742), .C(n37031), .Y(n37023) );
  OAI21X1 U31514 ( .A(n37032), .B(n37033), .C(n26480), .Y(n37031) );
  OAI22X1 U31515 ( .A(n34403), .B(n34751), .C(n37034), .D(n25106), .Y(n37033)
         );
  INVX1 U31516 ( .A(n34808), .Y(n37034) );
  NAND2X1 U31517 ( .A(n37035), .B(n37036), .Y(n34808) );
  AOI22X1 U31518 ( .A(reg_A[23]), .B(n25156), .C(n25142), .D(reg_A[24]), .Y(
        n37036) );
  AOI22X1 U31519 ( .A(reg_A[25]), .B(n25258), .C(reg_A[26]), .D(n26761), .Y(
        n37035) );
  NAND2X1 U31520 ( .A(reg_B[27]), .B(n34493), .Y(n34751) );
  AOI22X1 U31521 ( .A(n34809), .B(n33955), .C(reg_A[31]), .D(n35910), .Y(
        n34403) );
  INVX1 U31522 ( .A(n33872), .Y(n35910) );
  NAND2X1 U31523 ( .A(n25156), .B(reg_B[29]), .Y(n33872) );
  NAND2X1 U31524 ( .A(n37037), .B(n37038), .Y(n34809) );
  AOI22X1 U31525 ( .A(reg_A[27]), .B(n25156), .C(n25142), .D(reg_A[28]), .Y(
        n37038) );
  AOI22X1 U31526 ( .A(reg_A[29]), .B(n25258), .C(reg_A[30]), .D(n26761), .Y(
        n37037) );
  OAI22X1 U31527 ( .A(n28031), .B(n28033), .C(n28034), .D(n25099), .Y(n37032)
         );
  INVX1 U31528 ( .A(n35394), .Y(n28034) );
  NAND2X1 U31529 ( .A(n37039), .B(n37040), .Y(n35394) );
  AOI22X1 U31530 ( .A(reg_A[19]), .B(n25156), .C(n25142), .D(reg_A[20]), .Y(
        n37040) );
  AOI22X1 U31531 ( .A(reg_A[21]), .B(n25258), .C(reg_A[22]), .D(n26761), .Y(
        n37039) );
  INVX1 U31532 ( .A(n32983), .Y(n28031) );
  NAND2X1 U31533 ( .A(n37041), .B(n37042), .Y(n32983) );
  AOI22X1 U31534 ( .A(reg_A[15]), .B(n25156), .C(n25142), .D(reg_A[16]), .Y(
        n37042) );
  AOI22X1 U31535 ( .A(reg_A[17]), .B(n25258), .C(reg_A[18]), .D(n26761), .Y(
        n37041) );
  INVX1 U31536 ( .A(n28590), .Y(n32522) );
  AOI22X1 U31537 ( .A(n25172), .B(n35957), .C(n28572), .D(reg_A[2]), .Y(n37021) );
  AOI22X1 U31538 ( .A(n28576), .B(reg_A[5]), .C(n25181), .D(reg_A[7]), .Y(
        n37020) );
  NAND3X1 U31539 ( .A(n37043), .B(n37044), .C(n37045), .Y(n37018) );
  NOR2X1 U31540 ( .A(n37046), .B(n37047), .Y(n37045) );
  OAI21X1 U31541 ( .A(n37048), .B(n26701), .C(n37049), .Y(n37047) );
  OAI21X1 U31542 ( .A(n37050), .B(n37051), .C(n25310), .Y(n37049) );
  NAND3X1 U31543 ( .A(n37052), .B(n37053), .C(n37054), .Y(n37051) );
  NOR2X1 U31544 ( .A(n37055), .B(n37056), .Y(n37054) );
  OAI22X1 U31545 ( .A(n27967), .B(n25228), .C(n27962), .D(n25229), .Y(n37056)
         );
  OAI21X1 U31546 ( .A(n26714), .B(n25231), .C(n37057), .Y(n37055) );
  AOI22X1 U31547 ( .A(n25234), .B(reg_A[25]), .C(n25235), .D(reg_A[26]), .Y(
        n37057) );
  INVX1 U31548 ( .A(reg_A[23]), .Y(n26714) );
  AOI21X1 U31549 ( .A(reg_A[19]), .B(n25124), .C(n37058), .Y(n37053) );
  OAI22X1 U31550 ( .A(n25037), .B(n30587), .C(n25250), .D(n26703), .Y(n37058)
         );
  AOI22X1 U31551 ( .A(reg_A[22]), .B(n25222), .C(reg_A[21]), .D(n25637), .Y(
        n37052) );
  NAND3X1 U31552 ( .A(n37059), .B(n37060), .C(n37061), .Y(n37050) );
  NOR2X1 U31553 ( .A(n37062), .B(n37063), .Y(n37061) );
  OAI21X1 U31554 ( .A(n25042), .B(n25255), .C(n37064), .Y(n37063) );
  AOI22X1 U31555 ( .A(reg_A[29]), .B(n25241), .C(n25339), .D(reg_A[31]), .Y(
        n37064) );
  OAI21X1 U31556 ( .A(n25038), .B(n29286), .C(n37065), .Y(n37062) );
  AOI22X1 U31557 ( .A(reg_A[28]), .B(n25246), .C(reg_A[27]), .D(n25247), .Y(
        n37065) );
  AOI21X1 U31558 ( .A(reg_A[17]), .B(n25253), .C(n37066), .Y(n37060) );
  OAI22X1 U31559 ( .A(n25040), .B(n25206), .C(n25254), .D(n25208), .Y(n37066)
         );
  AOI22X1 U31560 ( .A(reg_A[18]), .B(n25628), .C(n25069), .D(reg_A[15]), .Y(
        n37059) );
  AOI21X1 U31561 ( .A(n30634), .B(n25110), .C(n32603), .Y(n37048) );
  OAI21X1 U31562 ( .A(n37067), .B(n37068), .C(n37069), .Y(n37046) );
  AOI22X1 U31563 ( .A(n37070), .B(n35969), .C(n37071), .D(n25382), .Y(n37069)
         );
  NOR2X1 U31564 ( .A(n35749), .B(n32996), .Y(n37071) );
  MUX2X1 U31565 ( .B(n28039), .A(n37072), .S(reg_B[13]), .Y(n32996) );
  NOR2X1 U31566 ( .A(n29279), .B(n26692), .Y(n37072) );
  NAND2X1 U31567 ( .A(n37073), .B(n37074), .Y(n28039) );
  AOI22X1 U31568 ( .A(reg_A[13]), .B(n26733), .C(reg_A[12]), .D(n25172), .Y(
        n37074) );
  AOI22X1 U31569 ( .A(reg_A[14]), .B(n26734), .C(n25116), .D(reg_A[11]), .Y(
        n37073) );
  INVX1 U31570 ( .A(n37075), .Y(n35749) );
  INVX1 U31571 ( .A(n37076), .Y(n35969) );
  OAI21X1 U31572 ( .A(reg_B[13]), .B(n35729), .C(n37077), .Y(n37076) );
  AOI21X1 U31573 ( .A(n26691), .B(n25196), .C(n37078), .Y(n37077) );
  MUX2X1 U31574 ( .B(reg_A[6]), .A(reg_A[7]), .S(n29302), .Y(n25196) );
  MUX2X1 U31575 ( .B(n37079), .A(n37080), .S(reg_B[15]), .Y(n35729) );
  MUX2X1 U31576 ( .B(reg_A[11]), .A(reg_A[3]), .S(reg_B[12]), .Y(n37079) );
  NOR2X1 U31577 ( .A(reg_B[14]), .B(n25032), .Y(n37070) );
  AOI22X1 U31578 ( .A(n37081), .B(n25170), .C(n26504), .D(n29302), .Y(n37068)
         );
  INVX1 U31579 ( .A(n36000), .Y(n37081) );
  INVX1 U31580 ( .A(n36039), .Y(n37067) );
  OAI22X1 U31581 ( .A(n25146), .B(n35857), .C(n27967), .D(n35888), .Y(n36039)
         );
  AOI22X1 U31582 ( .A(n35771), .B(n37082), .C(n35968), .D(n25192), .Y(n37044)
         );
  INVX1 U31583 ( .A(n37083), .Y(n25192) );
  OAI21X1 U31584 ( .A(reg_B[13]), .B(n35961), .C(n37084), .Y(n37083) );
  AOI21X1 U31585 ( .A(n26691), .B(n37085), .C(n37078), .Y(n37084) );
  AND2X1 U31586 ( .A(n35864), .B(n26742), .Y(n37078) );
  INVX1 U31587 ( .A(n35962), .Y(n37085) );
  MUX2X1 U31588 ( .B(n29265), .A(n30569), .S(reg_B[15]), .Y(n35962) );
  MUX2X1 U31589 ( .B(n37086), .A(n37087), .S(reg_B[15]), .Y(n35961) );
  MUX2X1 U31590 ( .B(reg_A[8]), .A(reg_A[0]), .S(reg_B[12]), .Y(n37087) );
  INVX1 U31591 ( .A(n34071), .Y(n35968) );
  NAND2X1 U31592 ( .A(n25188), .B(reg_B[14]), .Y(n34071) );
  AND2X1 U31593 ( .A(n36038), .B(n25170), .Y(n35771) );
  NOR2X1 U31594 ( .A(n29302), .B(n26999), .Y(n36038) );
  AOI22X1 U31595 ( .A(n28649), .B(reg_A[1]), .C(n28802), .D(reg_A[15]), .Y(
        n37043) );
  NOR2X1 U31596 ( .A(n37088), .B(n37089), .Y(n37016) );
  NAND3X1 U31597 ( .A(n37090), .B(n37091), .C(n37092), .Y(n37089) );
  NOR2X1 U31598 ( .A(n37093), .B(n37094), .Y(n37092) );
  OAI21X1 U31599 ( .A(n37095), .B(n25194), .C(n25088), .Y(n37094) );
  AOI21X1 U31600 ( .A(n25114), .B(reg_B[13]), .C(n37096), .Y(n25088) );
  OAI21X1 U31601 ( .A(n33955), .B(n25157), .C(n35646), .Y(n37096) );
  INVX1 U31602 ( .A(n37095), .Y(n25114) );
  OAI22X1 U31603 ( .A(n30569), .B(n28562), .C(n28032), .D(n30559), .Y(n37093)
         );
  INVX1 U31604 ( .A(n32982), .Y(n28032) );
  NAND2X1 U31605 ( .A(n37097), .B(n37098), .Y(n32982) );
  AOI22X1 U31606 ( .A(reg_A[11]), .B(n25156), .C(n25142), .D(reg_A[12]), .Y(
        n37098) );
  AOI22X1 U31607 ( .A(reg_A[13]), .B(n25258), .C(reg_A[14]), .D(n26761), .Y(
        n37097) );
  AOI22X1 U31608 ( .A(reg_A[11]), .B(n28661), .C(reg_A[10]), .D(n26626), .Y(
        n37091) );
  AOI22X1 U31609 ( .A(n37099), .B(n26756), .C(n37100), .D(n25119), .Y(n37090)
         );
  NAND3X1 U31610 ( .A(n37101), .B(n37102), .C(n37103), .Y(n37100) );
  NOR2X1 U31611 ( .A(n37104), .B(n37105), .Y(n37103) );
  OAI21X1 U31612 ( .A(n25132), .B(n26431), .C(n37106), .Y(n37105) );
  AOI22X1 U31613 ( .A(n25253), .B(reg_A[5]), .C(n25628), .D(reg_A[4]), .Y(
        n37106) );
  OAI21X1 U31614 ( .A(n25146), .B(n25133), .C(n37107), .Y(n37104) );
  AOI22X1 U31615 ( .A(reg_A[10]), .B(n25135), .C(n25136), .D(reg_A[8]), .Y(
        n37107) );
  AOI21X1 U31616 ( .A(n25124), .B(reg_A[3]), .C(n37108), .Y(n37102) );
  OAI22X1 U31617 ( .A(n25128), .B(n25223), .C(n26677), .D(n26703), .Y(n37108)
         );
  AOI22X1 U31618 ( .A(n25637), .B(reg_A[1]), .C(n25125), .D(reg_A[11]), .Y(
        n37101) );
  OAI21X1 U31619 ( .A(n25261), .B(n29305), .C(n37109), .Y(n37099) );
  AOI22X1 U31620 ( .A(n25156), .B(n36097), .C(n25142), .D(n37110), .Y(n37109)
         );
  INVX1 U31621 ( .A(n35955), .Y(n36097) );
  AOI22X1 U31622 ( .A(n35589), .B(n33955), .C(reg_A[7]), .D(n25101), .Y(n35955) );
  OAI22X1 U31623 ( .A(n33807), .B(n27967), .C(n25130), .D(n34465), .Y(n35589)
         );
  INVX1 U31624 ( .A(n36098), .Y(n25261) );
  NAND3X1 U31625 ( .A(n37111), .B(n37112), .C(n37113), .Y(n37088) );
  NOR2X1 U31626 ( .A(n37114), .B(n37115), .Y(n37113) );
  OAI22X1 U31627 ( .A(n25206), .B(n28569), .C(n25208), .D(n28570), .Y(n37115)
         );
  OAI21X1 U31628 ( .A(n26854), .B(n35919), .C(n37116), .Y(n37114) );
  AOI22X1 U31629 ( .A(n28717), .B(reg_A[3]), .C(n25149), .D(reg_A[6]), .Y(
        n37116) );
  INVX1 U31630 ( .A(n25178), .Y(n28717) );
  OAI21X1 U31631 ( .A(reg_B[2]), .B(n35752), .C(n37117), .Y(n35919) );
  AOI22X1 U31632 ( .A(n26455), .B(n26742), .C(n26456), .D(n28052), .Y(n37117)
         );
  INVX1 U31633 ( .A(n25167), .Y(n28052) );
  MUX2X1 U31634 ( .B(n25132), .A(n26677), .S(reg_B[4]), .Y(n25167) );
  INVX1 U31635 ( .A(n37118), .Y(n35752) );
  OAI21X1 U31636 ( .A(reg_B[4]), .B(n35527), .C(n37119), .Y(n37118) );
  AOI22X1 U31637 ( .A(n26462), .B(n25147), .C(n26463), .D(n25128), .Y(n37119)
         );
  MUX2X1 U31638 ( .B(n27967), .A(n25130), .S(reg_B[1]), .Y(n35527) );
  AOI22X1 U31639 ( .A(n28280), .B(reg_A[12]), .C(n30634), .D(n35754), .Y(
        n37112) );
  INVX1 U31640 ( .A(n27943), .Y(n30634) );
  NAND2X1 U31641 ( .A(n26761), .B(n25932), .Y(n27943) );
  AOI22X1 U31642 ( .A(n26761), .B(n25143), .C(n25151), .D(n26262), .Y(n37111)
         );
  AND2X1 U31643 ( .A(n37120), .B(n37121), .Y(n25151) );
  AOI22X1 U31644 ( .A(n26859), .B(n30569), .C(n26860), .D(n29265), .Y(n37121)
         );
  AOI22X1 U31645 ( .A(n26455), .B(n26742), .C(n35954), .D(n26452), .Y(n37120)
         );
  OAI21X1 U31646 ( .A(reg_A[0]), .B(n26861), .C(n37122), .Y(n35954) );
  AOI22X1 U31647 ( .A(n37123), .B(n26863), .C(n26462), .D(n26701), .Y(n37122)
         );
  INVX1 U31648 ( .A(n37124), .Y(n37123) );
  NAND3X1 U31649 ( .A(n37125), .B(n37126), .C(n37127), .Y(result[119]) );
  NOR2X1 U31650 ( .A(n37128), .B(n37129), .Y(n37127) );
  NAND3X1 U31651 ( .A(n37130), .B(n37131), .C(n37132), .Y(n37129) );
  AOI22X1 U31652 ( .A(n25310), .B(n37133), .C(n37134), .D(n37135), .Y(n37132)
         );
  NAND3X1 U31653 ( .A(n37136), .B(n37137), .C(n37138), .Y(n37133) );
  NOR2X1 U31654 ( .A(n37139), .B(n37140), .Y(n37138) );
  OAI22X1 U31655 ( .A(n25030), .B(n25319), .C(n25131), .D(n25317), .Y(n37140)
         );
  OAI21X1 U31656 ( .A(n25040), .B(n25490), .C(n37141), .Y(n37139) );
  AOI22X1 U31657 ( .A(reg_A[120]), .B(n25135), .C(reg_A[122]), .D(n25136), .Y(
        n37141) );
  AOI22X1 U31658 ( .A(reg_A[123]), .B(n25074), .C(reg_A[124]), .D(n25123), .Y(
        n37137) );
  AOI22X1 U31659 ( .A(reg_A[127]), .B(n25124), .C(reg_A[119]), .D(n25125), .Y(
        n37136) );
  OAI21X1 U31660 ( .A(n37142), .B(n37143), .C(n25730), .Y(n37131) );
  NAND2X1 U31661 ( .A(n37144), .B(n37145), .Y(n37143) );
  AOI22X1 U31662 ( .A(reg_A[123]), .B(n25749), .C(reg_A[124]), .D(n25750), .Y(
        n37145) );
  AOI22X1 U31663 ( .A(reg_A[127]), .B(n25615), .C(reg_A[119]), .D(n26924), .Y(
        n37144) );
  OR2X1 U31664 ( .A(n37146), .B(n37147), .Y(n37142) );
  OAI22X1 U31665 ( .A(n26936), .B(n25319), .C(n25745), .D(n25317), .Y(n37147)
         );
  OAI21X1 U31666 ( .A(n25062), .B(n25490), .C(n37148), .Y(n37146) );
  AOI22X1 U31667 ( .A(reg_A[120]), .B(n26803), .C(reg_A[122]), .D(n26804), .Y(
        n37148) );
  AOI22X1 U31668 ( .A(n37013), .B(n26028), .C(n37149), .D(n26260), .Y(n37130)
         );
  AND2X1 U31669 ( .A(n37150), .B(n37151), .Y(n37013) );
  AOI22X1 U31670 ( .A(n25025), .B(n36835), .C(n25026), .D(n36729), .Y(n37151)
         );
  INVX1 U31671 ( .A(n37152), .Y(n36835) );
  AOI22X1 U31672 ( .A(n26032), .B(n36728), .C(n26530), .D(n37153), .Y(n37150)
         );
  INVX1 U31673 ( .A(n36460), .Y(n36728) );
  NOR2X1 U31674 ( .A(n37154), .B(n37155), .Y(n36460) );
  OAI22X1 U31675 ( .A(reg_A[119]), .B(n26036), .C(reg_A[111]), .D(n26981), .Y(
        n37155) );
  OAI21X1 U31676 ( .A(reg_A[103]), .B(n26982), .C(n36952), .Y(n37154) );
  NAND2X1 U31677 ( .A(n37156), .B(n37157), .Y(n37128) );
  AOI21X1 U31678 ( .A(n36286), .B(n37158), .C(n37159), .Y(n37157) );
  OAI21X1 U31679 ( .A(n25335), .B(n27995), .C(n37160), .Y(n37159) );
  OAI21X1 U31680 ( .A(n37161), .B(n37162), .C(n26504), .Y(n37160) );
  OAI21X1 U31681 ( .A(n37163), .B(n37164), .C(n37165), .Y(n37162) );
  NAND3X1 U31682 ( .A(reg_B[117]), .B(reg_A[115]), .C(n37166), .Y(n37165) );
  MUX2X1 U31683 ( .B(n37167), .A(n37168), .S(reg_B[119]), .Y(n37161) );
  NAND2X1 U31684 ( .A(n37169), .B(reg_A[119]), .Y(n37167) );
  AOI22X1 U31685 ( .A(n37170), .B(n32116), .C(n36976), .D(n36329), .Y(n37156)
         );
  NOR2X1 U31686 ( .A(n37171), .B(n37172), .Y(n36976) );
  OAI22X1 U31687 ( .A(n36359), .B(n36453), .C(n36360), .D(n37173), .Y(n37172)
         );
  NOR2X1 U31688 ( .A(n37174), .B(n37175), .Y(n36453) );
  OAI22X1 U31689 ( .A(reg_A[111]), .B(n36318), .C(reg_A[119]), .D(n36668), .Y(
        n37175) );
  OAI21X1 U31690 ( .A(reg_A[103]), .B(n36957), .C(n36958), .Y(n37174) );
  OAI22X1 U31691 ( .A(n36312), .B(n36867), .C(n36439), .D(n37176), .Y(n37171)
         );
  NOR2X1 U31692 ( .A(n37177), .B(n37178), .Y(n37126) );
  NAND3X1 U31693 ( .A(n37179), .B(n37180), .C(n37181), .Y(n37178) );
  NAND2X1 U31694 ( .A(reg_A[119]), .B(n37182), .Y(n37181) );
  OAI21X1 U31695 ( .A(n28105), .B(n37183), .C(n34838), .Y(n37182) );
  INVX1 U31696 ( .A(n27046), .Y(n34838) );
  OAI21X1 U31697 ( .A(n26943), .B(n37184), .C(n25795), .Y(n27046) );
  NOR2X1 U31698 ( .A(n25170), .B(n25382), .Y(n28105) );
  OAI21X1 U31699 ( .A(n36297), .B(n27051), .C(reg_A[112]), .Y(n37180) );
  OAI21X1 U31700 ( .A(n25753), .B(n37184), .C(n37185), .Y(n27051) );
  NOR2X1 U31701 ( .A(n32498), .B(n37186), .Y(n37185) );
  NOR2X1 U31702 ( .A(n36231), .B(n25032), .Y(n36297) );
  NAND3X1 U31703 ( .A(n36355), .B(n25355), .C(n36235), .Y(n36231) );
  OAI21X1 U31704 ( .A(n36916), .B(n28004), .C(reg_A[116]), .Y(n37179) );
  INVX1 U31705 ( .A(n27095), .Y(n28004) );
  INVX1 U31706 ( .A(n36260), .Y(n36916) );
  NAND3X1 U31707 ( .A(n36356), .B(n25188), .C(n37187), .Y(n36260) );
  NOR2X1 U31708 ( .A(n36246), .B(n37188), .Y(n37187) );
  NAND3X1 U31709 ( .A(n37189), .B(n36887), .C(n37190), .Y(n37177) );
  OAI21X1 U31710 ( .A(n37191), .B(n37192), .C(n27067), .Y(n37190) );
  OAI21X1 U31711 ( .A(n25736), .B(n36140), .C(n37193), .Y(n37192) );
  AOI22X1 U31712 ( .A(reg_A[115]), .B(n25749), .C(reg_A[114]), .D(n25750), .Y(
        n37193) );
  NAND2X1 U31713 ( .A(n37194), .B(n37195), .Y(n37191) );
  AOI22X1 U31714 ( .A(reg_A[118]), .B(n26803), .C(reg_A[116]), .D(n26804), .Y(
        n37195) );
  AOI22X1 U31715 ( .A(reg_A[117]), .B(n26927), .C(reg_A[113]), .D(n26878), .Y(
        n37194) );
  OAI21X1 U31716 ( .A(n37196), .B(n37197), .C(n25840), .Y(n37189) );
  NAND2X1 U31717 ( .A(n37198), .B(n37199), .Y(n37197) );
  NOR2X1 U31718 ( .A(n37200), .B(n37201), .Y(n37199) );
  OAI21X1 U31719 ( .A(n25043), .B(n36140), .C(n37202), .Y(n37201) );
  AOI22X1 U31720 ( .A(reg_A[118]), .B(n25135), .C(reg_A[117]), .D(n25252), .Y(
        n37202) );
  OAI21X1 U31721 ( .A(n25028), .B(n25771), .C(n37203), .Y(n37200) );
  AOI22X1 U31722 ( .A(reg_A[116]), .B(n25136), .C(reg_A[115]), .D(n25067), .Y(
        n37203) );
  NOR2X1 U31723 ( .A(n37204), .B(n37205), .Y(n37198) );
  OAI21X1 U31724 ( .A(n25034), .B(n25452), .C(n37206), .Y(n37205) );
  AOI22X1 U31725 ( .A(reg_A[113]), .B(n25253), .C(reg_A[112]), .D(n25628), .Y(
        n37206) );
  OAI21X1 U31726 ( .A(n25036), .B(n25474), .C(n37207), .Y(n37204) );
  AOI22X1 U31727 ( .A(reg_A[110]), .B(n25629), .C(reg_A[108]), .D(n25222), .Y(
        n37207) );
  NAND2X1 U31728 ( .A(n37208), .B(n37209), .Y(n37196) );
  NOR2X1 U31729 ( .A(n37210), .B(n37211), .Y(n37209) );
  OAI21X1 U31730 ( .A(n25039), .B(n25468), .C(n37212), .Y(n37211) );
  AOI22X1 U31731 ( .A(reg_A[105]), .B(n25234), .C(reg_A[107]), .D(n25635), .Y(
        n37212) );
  OAI21X1 U31732 ( .A(n25065), .B(n25298), .C(n37213), .Y(n37210) );
  AOI22X1 U31733 ( .A(reg_A[102]), .B(n25246), .C(reg_A[103]), .D(n25247), .Y(
        n37213) );
  NOR2X1 U31734 ( .A(n37214), .B(n37215), .Y(n37208) );
  OAI21X1 U31735 ( .A(n25238), .B(n25396), .C(n37216), .Y(n37215) );
  AOI22X1 U31736 ( .A(reg_A[100]), .B(n25487), .C(reg_A[101]), .D(n25241), .Y(
        n37216) );
  OAI21X1 U31737 ( .A(n26719), .B(n25289), .C(n37217), .Y(n37214) );
  AOI22X1 U31738 ( .A(reg_A[97]), .B(n25242), .C(n25338), .D(reg_A[96]), .Y(
        n37217) );
  NOR2X1 U31739 ( .A(n37218), .B(n37219), .Y(n37125) );
  OAI21X1 U31740 ( .A(n37220), .B(n37184), .C(n37221), .Y(n37219) );
  OAI21X1 U31741 ( .A(n37222), .B(n37223), .C(n25170), .Y(n37221) );
  OAI21X1 U31742 ( .A(n25332), .B(n37224), .C(n37225), .Y(n37223) );
  AOI22X1 U31743 ( .A(n37226), .B(n37001), .C(n37227), .D(n37228), .Y(n37225)
         );
  INVX1 U31744 ( .A(n37229), .Y(n37227) );
  NAND2X1 U31745 ( .A(n37230), .B(n37231), .Y(n37001) );
  AOI22X1 U31746 ( .A(n36315), .B(n36447), .C(n36442), .D(n36681), .Y(n37231)
         );
  OAI21X1 U31747 ( .A(n25452), .B(n36318), .C(n37232), .Y(n36447) );
  AOI22X1 U31748 ( .A(n36685), .B(reg_A[103]), .C(n36338), .D(reg_A[119]), .Y(
        n37232) );
  AOI22X1 U31749 ( .A(n36649), .B(n36901), .C(n36280), .D(n37233), .Y(n37230)
         );
  OAI21X1 U31750 ( .A(n37234), .B(n37235), .C(n37236), .Y(n37222) );
  AOI22X1 U31751 ( .A(n37237), .B(n37238), .C(n25604), .D(n37239), .Y(n37236)
         );
  OAI21X1 U31752 ( .A(n37240), .B(n36246), .C(n37241), .Y(n37239) );
  INVX1 U31753 ( .A(n37158), .Y(n37241) );
  OAI21X1 U31754 ( .A(n37242), .B(n36136), .C(n37243), .Y(n37158) );
  AOI22X1 U31755 ( .A(n25793), .B(n36780), .C(n25700), .D(n36902), .Y(n37243)
         );
  OAI22X1 U31756 ( .A(n36236), .B(n36140), .C(n25335), .D(n36247), .Y(n36780)
         );
  MUX2X1 U31757 ( .B(n25335), .A(n25483), .S(reg_B[118]), .Y(n37238) );
  NOR2X1 U31758 ( .A(reg_B[119]), .B(n37244), .Y(n37237) );
  AOI21X1 U31759 ( .A(reg_A[113]), .B(n26010), .C(n37245), .Y(n37220) );
  OAI22X1 U31760 ( .A(n31144), .B(n25332), .C(n27925), .D(n25333), .Y(n37245)
         );
  OAI21X1 U31761 ( .A(n25771), .B(n27108), .C(n37246), .Y(n37218) );
  AOI22X1 U31762 ( .A(n36271), .B(n27110), .C(n37247), .D(n36294), .Y(n37246)
         );
  INVX1 U31763 ( .A(n28053), .Y(n27110) );
  MUX2X1 U31764 ( .B(n36140), .A(n25333), .S(reg_B[4]), .Y(n36271) );
  NAND2X1 U31765 ( .A(n37248), .B(n37249), .Y(result[118]) );
  NOR2X1 U31766 ( .A(n37250), .B(n37251), .Y(n37249) );
  NAND3X1 U31767 ( .A(n37252), .B(n37253), .C(n37254), .Y(n37251) );
  NOR2X1 U31768 ( .A(n37255), .B(n37256), .Y(n37254) );
  OAI21X1 U31769 ( .A(n25332), .B(n33978), .C(n37257), .Y(n37256) );
  OAI21X1 U31770 ( .A(n37258), .B(n37259), .C(n26504), .Y(n37257) );
  INVX1 U31771 ( .A(n37260), .Y(n37259) );
  MUX2X1 U31772 ( .B(n37261), .A(n37262), .S(reg_B[119]), .Y(n37260) );
  OAI22X1 U31773 ( .A(n36747), .B(n37263), .C(n27190), .D(n36345), .Y(n37255)
         );
  NAND2X1 U31774 ( .A(n37264), .B(n37265), .Y(n36345) );
  AOI22X1 U31775 ( .A(n26601), .B(n25337), .C(n26602), .D(n25335), .Y(n37265)
         );
  AOI22X1 U31776 ( .A(n27012), .B(n25333), .C(n26597), .D(n25332), .Y(n37264)
         );
  AOI22X1 U31777 ( .A(n37247), .B(n36329), .C(reg_A[114]), .D(n31307), .Y(
        n37253) );
  AND2X1 U31778 ( .A(n37266), .B(n37267), .Y(n37247) );
  AOI22X1 U31779 ( .A(n36315), .B(n36820), .C(n36442), .D(n36821), .Y(n37267)
         );
  INVX1 U31780 ( .A(n36608), .Y(n36820) );
  NOR2X1 U31781 ( .A(n37268), .B(n37269), .Y(n36608) );
  OAI22X1 U31782 ( .A(reg_A[110]), .B(n36318), .C(reg_A[118]), .D(n36668), .Y(
        n37269) );
  OAI21X1 U31783 ( .A(reg_A[102]), .B(n36957), .C(n36958), .Y(n37268) );
  AOI22X1 U31784 ( .A(n36280), .B(n37270), .C(n36649), .D(n36959), .Y(n37266)
         );
  INVX1 U31785 ( .A(n37271), .Y(n36959) );
  AOI22X1 U31786 ( .A(reg_A[112]), .B(n27192), .C(reg_A[113]), .D(n27256), .Y(
        n37252) );
  NAND3X1 U31787 ( .A(n37272), .B(n37273), .C(n37274), .Y(n37250) );
  NOR2X1 U31788 ( .A(n37275), .B(n37276), .Y(n37274) );
  OAI22X1 U31789 ( .A(n36971), .B(n36415), .C(n25335), .D(n33975), .Y(n37276)
         );
  NAND2X1 U31790 ( .A(n25793), .B(n36702), .Y(n36415) );
  INVX1 U31791 ( .A(n36902), .Y(n36971) );
  OAI22X1 U31792 ( .A(n36236), .B(n25333), .C(n25771), .D(n36247), .Y(n36902)
         );
  OAI21X1 U31793 ( .A(n37277), .B(n25337), .C(n37278), .Y(n37275) );
  OAI21X1 U31794 ( .A(n33961), .B(n25283), .C(reg_A[118]), .Y(n37278) );
  INVX1 U31795 ( .A(n34999), .Y(n33961) );
  AOI21X1 U31796 ( .A(n37279), .B(n36286), .C(n27183), .Y(n37277) );
  NOR2X1 U31797 ( .A(n36236), .B(n36136), .Y(n37279) );
  AOI21X1 U31798 ( .A(n37280), .B(n37281), .C(n37282), .Y(n37273) );
  OAI21X1 U31799 ( .A(n37283), .B(n37284), .C(n36887), .Y(n37282) );
  NAND2X1 U31800 ( .A(n36286), .B(n37285), .Y(n36887) );
  NAND2X1 U31801 ( .A(n36286), .B(reg_B[126]), .Y(n37284) );
  NOR2X1 U31802 ( .A(reg_B[118]), .B(n37286), .Y(n37280) );
  AOI22X1 U31803 ( .A(n37287), .B(reg_B[127]), .C(n37288), .D(n25399), .Y(
        n37272) );
  NOR2X1 U31804 ( .A(n37240), .B(n25023), .Y(n37288) );
  AND2X1 U31805 ( .A(n36702), .B(n37289), .Y(n37287) );
  INVX1 U31806 ( .A(n36322), .Y(n36702) );
  NOR2X1 U31807 ( .A(n26267), .B(n36286), .Y(n36322) );
  NOR2X1 U31808 ( .A(n37290), .B(n37291), .Y(n37248) );
  NAND3X1 U31809 ( .A(n37292), .B(n37293), .C(n37294), .Y(n37291) );
  NOR2X1 U31810 ( .A(n37295), .B(n37296), .Y(n37294) );
  INVX1 U31811 ( .A(n37297), .Y(n37296) );
  AOI22X1 U31812 ( .A(n37134), .B(n37298), .C(n37262), .D(n37299), .Y(n37297)
         );
  OAI22X1 U31813 ( .A(n37300), .B(n37301), .C(n37302), .D(n37303), .Y(n37295)
         );
  INVX1 U31814 ( .A(n37228), .Y(n37302) );
  NAND2X1 U31815 ( .A(n37304), .B(n37305), .Y(n37228) );
  AOI22X1 U31816 ( .A(n36315), .B(n36582), .C(n36442), .D(n36774), .Y(n37305)
         );
  OAI21X1 U31817 ( .A(n25450), .B(n36318), .C(n37306), .Y(n36582) );
  AOI22X1 U31818 ( .A(n36685), .B(reg_A[102]), .C(n36338), .D(reg_A[118]), .Y(
        n37306) );
  AOI22X1 U31819 ( .A(n36649), .B(n37007), .C(n36280), .D(n37307), .Y(n37304)
         );
  AOI22X1 U31820 ( .A(reg_A[125]), .B(n25293), .C(reg_A[119]), .D(n25282), .Y(
        n37293) );
  AOI22X1 U31821 ( .A(n26045), .B(n37308), .C(n37309), .D(n37310), .Y(n37292)
         );
  INVX1 U31822 ( .A(n37234), .Y(n37310) );
  NOR2X1 U31823 ( .A(n37261), .B(n37258), .Y(n37234) );
  OAI21X1 U31824 ( .A(n25337), .B(n37311), .C(n37168), .Y(n37261) );
  AOI22X1 U31825 ( .A(reg_A[118]), .B(n37169), .C(reg_A[114]), .D(n37312), .Y(
        n37168) );
  NAND3X1 U31826 ( .A(n37313), .B(n37314), .C(n37315), .Y(n37308) );
  NOR2X1 U31827 ( .A(n37316), .B(n37317), .Y(n37315) );
  OAI22X1 U31828 ( .A(n27218), .B(n25332), .C(n25207), .D(n25483), .Y(n37317)
         );
  OAI21X1 U31829 ( .A(n27219), .B(n25476), .C(n37318), .Y(n37316) );
  OAI21X1 U31830 ( .A(n37319), .B(n37320), .C(n25044), .Y(n37318) );
  NAND3X1 U31831 ( .A(n37321), .B(n37322), .C(n37323), .Y(n37320) );
  NOR2X1 U31832 ( .A(n37324), .B(n37325), .Y(n37323) );
  OAI21X1 U31833 ( .A(n25036), .B(n25469), .C(n37326), .Y(n37325) );
  AOI22X1 U31834 ( .A(reg_A[110]), .B(n25124), .C(reg_A[107]), .D(n25222), .Y(
        n37326) );
  OAI21X1 U31835 ( .A(n25037), .B(n25474), .C(n37327), .Y(n37324) );
  AOI22X1 U31836 ( .A(reg_A[114]), .B(n25074), .C(reg_A[113]), .D(n25123), .Y(
        n37327) );
  AOI21X1 U31837 ( .A(reg_A[106]), .B(n25635), .C(n37328), .Y(n37322) );
  OAI22X1 U31838 ( .A(n25065), .B(n25448), .C(n25035), .D(n25298), .Y(n37328)
         );
  AOI22X1 U31839 ( .A(reg_A[105]), .B(n25325), .C(reg_A[118]), .D(n25125), .Y(
        n37321) );
  NAND2X1 U31840 ( .A(n37329), .B(n37330), .Y(n37319) );
  NOR2X1 U31841 ( .A(n37331), .B(n37332), .Y(n37330) );
  OAI21X1 U31842 ( .A(n25238), .B(n25289), .C(n37333), .Y(n37332) );
  AOI22X1 U31843 ( .A(reg_A[100]), .B(n25241), .C(reg_A[96]), .D(n25242), .Y(
        n37333) );
  OAI21X1 U31844 ( .A(n25038), .B(n25396), .C(n37334), .Y(n37331) );
  AOI22X1 U31845 ( .A(reg_A[101]), .B(n25246), .C(reg_A[102]), .D(n25247), .Y(
        n37334) );
  NOR2X1 U31846 ( .A(n37335), .B(n37336), .Y(n37329) );
  OAI21X1 U31847 ( .A(n25030), .B(n25452), .C(n37337), .Y(n37336) );
  AOI22X1 U31848 ( .A(reg_A[116]), .B(n25252), .C(reg_A[112]), .D(n25253), .Y(
        n37337) );
  OAI21X1 U31849 ( .A(n25041), .B(n25335), .C(n37338), .Y(n37335) );
  AOI22X1 U31850 ( .A(reg_A[97]), .B(n25257), .C(reg_A[117]), .D(n25135), .Y(
        n37338) );
  AOI22X1 U31851 ( .A(reg_A[115]), .B(n27241), .C(reg_A[114]), .D(n27242), .Y(
        n37314) );
  AOI22X1 U31852 ( .A(reg_A[116]), .B(n27243), .C(reg_A[118]), .D(n25434), .Y(
        n37313) );
  NAND3X1 U31853 ( .A(n37339), .B(n37340), .C(n37341), .Y(n37290) );
  NOR2X1 U31854 ( .A(n37342), .B(n37343), .Y(n37341) );
  OAI22X1 U31855 ( .A(n27938), .B(n25493), .C(n27512), .D(n25319), .Y(n37343)
         );
  OAI21X1 U31856 ( .A(n31590), .B(n25497), .C(n37344), .Y(n37342) );
  AOI22X1 U31857 ( .A(n37149), .B(n26028), .C(n37345), .D(n26260), .Y(n37344)
         );
  INVX1 U31858 ( .A(n37346), .Y(n37345) );
  AND2X1 U31859 ( .A(n37347), .B(n37348), .Y(n37149) );
  AOI22X1 U31860 ( .A(n25025), .B(n36949), .C(n25026), .D(n36800), .Y(n37348)
         );
  INVX1 U31861 ( .A(n37349), .Y(n36949) );
  AOI22X1 U31862 ( .A(n26032), .B(n36799), .C(n26530), .D(n37350), .Y(n37347)
         );
  INVX1 U31863 ( .A(n36598), .Y(n36799) );
  NOR2X1 U31864 ( .A(n37351), .B(n37352), .Y(n36598) );
  OAI22X1 U31865 ( .A(reg_A[118]), .B(n25063), .C(reg_A[110]), .D(n25058), .Y(
        n37352) );
  OAI21X1 U31866 ( .A(reg_A[102]), .B(n26982), .C(n36952), .Y(n37351) );
  INVX1 U31867 ( .A(n25301), .Y(n31590) );
  AOI22X1 U31868 ( .A(reg_A[121]), .B(n29051), .C(reg_A[122]), .D(n29029), .Y(
        n37340) );
  AOI22X1 U31869 ( .A(reg_A[123]), .B(n29030), .C(reg_A[124]), .D(n29031), .Y(
        n37339) );
  NAND3X1 U31870 ( .A(n37353), .B(n37354), .C(n37355), .Y(result[117]) );
  NOR2X1 U31871 ( .A(n37356), .B(n37357), .Y(n37355) );
  NAND3X1 U31872 ( .A(n37358), .B(n37359), .C(n37360), .Y(n37357) );
  AOI22X1 U31873 ( .A(n37361), .B(n36329), .C(reg_A[119]), .D(n26783), .Y(
        n37360) );
  INVX1 U31874 ( .A(n37263), .Y(n37361) );
  OAI21X1 U31875 ( .A(n37176), .B(n36312), .C(n37362), .Y(n37263) );
  AOI22X1 U31876 ( .A(n36315), .B(n36651), .C(reg_B[126]), .D(n37363), .Y(
        n37362) );
  INVX1 U31877 ( .A(n37173), .Y(n36651) );
  NOR2X1 U31878 ( .A(n37364), .B(n37365), .Y(n37173) );
  OAI22X1 U31879 ( .A(reg_A[109]), .B(n36318), .C(reg_A[117]), .D(n36668), .Y(
        n37365) );
  OAI21X1 U31880 ( .A(reg_A[101]), .B(n36957), .C(n36958), .Y(n37364) );
  OAI21X1 U31881 ( .A(n37366), .B(n37367), .C(n25730), .Y(n37359) );
  NAND2X1 U31882 ( .A(n37368), .B(n37369), .Y(n37367) );
  AOI22X1 U31883 ( .A(reg_A[122]), .B(n25750), .C(reg_A[126]), .D(n25614), .Y(
        n37369) );
  AOI22X1 U31884 ( .A(reg_A[125]), .B(n25615), .C(reg_A[127]), .D(n25607), .Y(
        n37368) );
  NAND2X1 U31885 ( .A(n37370), .B(n37371), .Y(n37366) );
  AOI22X1 U31886 ( .A(reg_A[120]), .B(n26804), .C(reg_A[123]), .D(n26878), .Y(
        n37371) );
  AOI22X1 U31887 ( .A(reg_A[124]), .B(n25613), .C(reg_A[121]), .D(n25749), .Y(
        n37370) );
  AOI22X1 U31888 ( .A(n37372), .B(n36294), .C(reg_A[117]), .D(n32829), .Y(
        n37358) );
  NAND2X1 U31889 ( .A(n25795), .B(n33195), .Y(n32829) );
  INVX1 U31890 ( .A(n36747), .Y(n36294) );
  NAND2X1 U31891 ( .A(reg_B[127]), .B(n25932), .Y(n36747) );
  NAND2X1 U31892 ( .A(n37373), .B(n37374), .Y(n37356) );
  AOI21X1 U31893 ( .A(n26504), .B(n37375), .C(n37376), .Y(n37374) );
  OAI21X1 U31894 ( .A(n37377), .B(n37378), .C(n37379), .Y(n37376) );
  NAND2X1 U31895 ( .A(n37289), .B(n36172), .Y(n37378) );
  OAI22X1 U31896 ( .A(reg_B[126]), .B(n37242), .C(n25335), .D(n37380), .Y(
        n37289) );
  INVX1 U31897 ( .A(n36975), .Y(n37242) );
  OAI22X1 U31898 ( .A(n36236), .B(n25332), .C(n25483), .D(n36247), .Y(n36975)
         );
  OAI21X1 U31899 ( .A(reg_B[118]), .B(n37164), .C(n37381), .Y(n37375) );
  AOI21X1 U31900 ( .A(n37382), .B(n37383), .C(n37258), .Y(n37381) );
  INVX1 U31901 ( .A(n37384), .Y(n37258) );
  NAND3X1 U31902 ( .A(reg_B[117]), .B(reg_A[112]), .C(reg_B[118]), .Y(n37384)
         );
  MUX2X1 U31903 ( .B(n25335), .A(n25771), .S(reg_B[119]), .Y(n37382) );
  INVX1 U31904 ( .A(n37385), .Y(n37164) );
  MUX2X1 U31905 ( .B(n37386), .A(n37387), .S(reg_B[119]), .Y(n37385) );
  MUX2X1 U31906 ( .B(reg_A[116]), .A(reg_A[112]), .S(reg_B[117]), .Y(n37387)
         );
  MUX2X1 U31907 ( .B(reg_A[117]), .A(reg_A[113]), .S(reg_B[117]), .Y(n37386)
         );
  AOI22X1 U31908 ( .A(n25372), .B(n37388), .C(n37389), .D(n37390), .Y(n37373)
         );
  OAI21X1 U31909 ( .A(n37391), .B(n37392), .C(n37393), .Y(n37388) );
  NAND3X1 U31910 ( .A(n36961), .B(n36437), .C(n37394), .Y(n37393) );
  NOR2X1 U31911 ( .A(n25476), .B(n37188), .Y(n37394) );
  INVX1 U31912 ( .A(n36429), .Y(n37391) );
  OAI22X1 U31913 ( .A(n25337), .B(n25568), .C(n25771), .D(n36246), .Y(n36429)
         );
  NOR2X1 U31914 ( .A(n37395), .B(n37396), .Y(n37354) );
  OAI21X1 U31915 ( .A(n37300), .B(n37303), .C(n37397), .Y(n37396) );
  OAI21X1 U31916 ( .A(n37398), .B(n37399), .C(n25310), .Y(n37397) );
  OR2X1 U31917 ( .A(n37400), .B(n37401), .Y(n37399) );
  OAI22X1 U31918 ( .A(n25043), .B(n25332), .C(n25219), .D(n25497), .Y(n37401)
         );
  OAI21X1 U31919 ( .A(n25034), .B(n25317), .C(n37402), .Y(n37400) );
  AOI22X1 U31920 ( .A(reg_A[122]), .B(n25123), .C(reg_A[126]), .D(n25629), .Y(
        n37402) );
  OR2X1 U31921 ( .A(n37403), .B(n37404), .Y(n37398) );
  OAI21X1 U31922 ( .A(n25056), .B(n25490), .C(n37405), .Y(n37404) );
  AOI22X1 U31923 ( .A(reg_A[123]), .B(n25253), .C(reg_A[124]), .D(n25628), .Y(
        n37405) );
  OAI21X1 U31924 ( .A(n25040), .B(n36140), .C(n37406), .Y(n37403) );
  AOI22X1 U31925 ( .A(reg_A[118]), .B(n25135), .C(reg_A[120]), .D(n25136), .Y(
        n37406) );
  AND2X1 U31926 ( .A(n37407), .B(n37408), .Y(n37300) );
  AOI22X1 U31927 ( .A(n36315), .B(n36681), .C(n36442), .D(n36901), .Y(n37408)
         );
  OAI21X1 U31928 ( .A(n25474), .B(n36318), .C(n37409), .Y(n36681) );
  AOI22X1 U31929 ( .A(n36685), .B(reg_A[101]), .C(n36338), .D(reg_A[117]), .Y(
        n37409) );
  AOI22X1 U31930 ( .A(n36649), .B(n37233), .C(n36280), .D(n37410), .Y(n37407)
         );
  OAI21X1 U31931 ( .A(n37411), .B(n31658), .C(n37412), .Y(n37395) );
  AOI22X1 U31932 ( .A(reg_A[118]), .B(n28923), .C(n26045), .D(n37413), .Y(
        n37412) );
  NAND3X1 U31933 ( .A(n37414), .B(n37415), .C(n37416), .Y(n37413) );
  AOI21X1 U31934 ( .A(reg_A[116]), .B(n25441), .C(n37417), .Y(n37416) );
  OAI21X1 U31935 ( .A(n25207), .B(n25476), .C(n37418), .Y(n37417) );
  OAI21X1 U31936 ( .A(n37419), .B(n37420), .C(n25044), .Y(n37418) );
  NAND3X1 U31937 ( .A(n37421), .B(n37422), .C(n37423), .Y(n37420) );
  NOR2X1 U31938 ( .A(n37424), .B(n37425), .Y(n37423) );
  OAI21X1 U31939 ( .A(n25036), .B(n25470), .C(n37426), .Y(n37425) );
  AOI22X1 U31940 ( .A(reg_A[109]), .B(n25124), .C(reg_A[106]), .D(n25222), .Y(
        n37426) );
  OAI21X1 U31941 ( .A(n25037), .B(n25469), .C(n37427), .Y(n37424) );
  AOI22X1 U31942 ( .A(reg_A[113]), .B(n25074), .C(reg_A[112]), .D(n25123), .Y(
        n37427) );
  AOI21X1 U31943 ( .A(reg_A[105]), .B(n25635), .C(n37428), .Y(n37422) );
  OAI22X1 U31944 ( .A(n25065), .B(n25361), .C(n25035), .D(n25448), .Y(n37428)
         );
  AOI22X1 U31945 ( .A(reg_A[104]), .B(n25325), .C(reg_A[117]), .D(n25125), .Y(
        n37421) );
  NAND3X1 U31946 ( .A(n37429), .B(n37430), .C(n37431), .Y(n37419) );
  NOR2X1 U31947 ( .A(n37432), .B(n37433), .Y(n37431) );
  OAI21X1 U31948 ( .A(n26719), .B(n25424), .C(n37434), .Y(n37433) );
  AOI22X1 U31949 ( .A(reg_A[99]), .B(n25241), .C(reg_A[97]), .D(n25339), .Y(
        n37434) );
  OAI21X1 U31950 ( .A(n25038), .B(n25289), .C(n37435), .Y(n37432) );
  AOI22X1 U31951 ( .A(reg_A[100]), .B(n25246), .C(reg_A[101]), .D(n25247), .Y(
        n37435) );
  AOI21X1 U31952 ( .A(reg_A[115]), .B(n25252), .C(n37436), .Y(n37430) );
  OAI22X1 U31953 ( .A(n25041), .B(n25771), .C(n25042), .D(n25337), .Y(n37436)
         );
  AOI22X1 U31954 ( .A(reg_A[111]), .B(n25253), .C(reg_A[110]), .D(n25628), .Y(
        n37429) );
  AOI22X1 U31955 ( .A(reg_A[113]), .B(n27242), .C(reg_A[117]), .D(n25434), .Y(
        n37414) );
  INVX1 U31956 ( .A(n37437), .Y(n37411) );
  NAND3X1 U31957 ( .A(n37438), .B(n37439), .C(n37440), .Y(n37437) );
  NOR2X1 U31958 ( .A(n37441), .B(n37442), .Y(n37440) );
  OAI21X1 U31959 ( .A(n25332), .B(n27442), .C(n37415), .Y(n37442) );
  AOI22X1 U31960 ( .A(n27243), .B(reg_A[115]), .C(n27241), .D(reg_A[114]), .Y(
        n37415) );
  OAI22X1 U31961 ( .A(n25483), .B(n25438), .C(n25337), .D(n28303), .Y(n37441)
         );
  INVX1 U31962 ( .A(n37443), .Y(n37439) );
  OAI22X1 U31963 ( .A(n37444), .B(n27379), .C(n37346), .D(n27377), .Y(n37443)
         );
  NAND2X1 U31964 ( .A(n25044), .B(n26863), .Y(n27377) );
  OAI21X1 U31965 ( .A(n37445), .B(n26030), .C(n37446), .Y(n37346) );
  AOI22X1 U31966 ( .A(n25025), .B(n37153), .C(n26032), .D(n36729), .Y(n37446)
         );
  OR2X1 U31967 ( .A(n37447), .B(n37448), .Y(n36729) );
  OAI22X1 U31968 ( .A(reg_A[117]), .B(n26036), .C(reg_A[109]), .D(n25058), .Y(
        n37448) );
  OAI21X1 U31969 ( .A(reg_A[101]), .B(n25055), .C(n36952), .Y(n37447) );
  INVX1 U31970 ( .A(n37449), .Y(n37153) );
  INVX1 U31971 ( .A(n37450), .Y(n37445) );
  NAND2X1 U31972 ( .A(reg_B[4]), .B(n25044), .Y(n27379) );
  AOI22X1 U31973 ( .A(n37170), .B(n29345), .C(reg_A[112]), .D(n37451), .Y(
        n37438) );
  AND2X1 U31974 ( .A(n37452), .B(n36473), .Y(n37170) );
  AOI22X1 U31975 ( .A(n25337), .B(n26295), .C(n25332), .D(n26293), .Y(n36473)
         );
  AOI22X1 U31976 ( .A(n26292), .B(n25483), .C(n26294), .D(n25476), .Y(n37452)
         );
  NOR2X1 U31977 ( .A(n37453), .B(n37454), .Y(n37353) );
  INVX1 U31978 ( .A(n37455), .Y(n37454) );
  AOI22X1 U31979 ( .A(n37134), .B(n37456), .C(n37457), .D(n37281), .Y(n37455)
         );
  OAI21X1 U31980 ( .A(n37458), .B(n37459), .C(n37460), .Y(n37453) );
  AOI22X1 U31981 ( .A(n37309), .B(n37262), .C(n25275), .D(n37461), .Y(n37460)
         );
  OAI21X1 U31982 ( .A(n25332), .B(n37462), .C(n37463), .Y(n37262) );
  AOI22X1 U31983 ( .A(n37312), .B(reg_A[113]), .C(n37383), .D(reg_A[115]), .Y(
        n37463) );
  INVX1 U31984 ( .A(n37464), .Y(n37458) );
  NAND3X1 U31985 ( .A(n37465), .B(n37466), .C(n37467), .Y(result[116]) );
  NOR2X1 U31986 ( .A(n37468), .B(n37469), .Y(n37467) );
  OR2X1 U31987 ( .A(n37470), .B(n37471), .Y(n37469) );
  OAI21X1 U31988 ( .A(n37472), .B(n37459), .C(n37473), .Y(n37471) );
  AOI22X1 U31989 ( .A(n37474), .B(n37134), .C(n25275), .D(n37475), .Y(n37473)
         );
  OAI21X1 U31990 ( .A(reg_B[123]), .B(n26996), .C(n27500), .Y(n37134) );
  NAND2X1 U31991 ( .A(n25382), .B(n25604), .Y(n27500) );
  OAI21X1 U31992 ( .A(n37476), .B(n37477), .C(n37478), .Y(n37470) );
  AOI22X1 U31993 ( .A(n25277), .B(n37461), .C(n37309), .D(n37464), .Y(n37478)
         );
  OAI21X1 U31994 ( .A(n25337), .B(n37462), .C(n37479), .Y(n37464) );
  AOI22X1 U31995 ( .A(n37312), .B(reg_A[112]), .C(n37383), .D(reg_A[114]), .Y(
        n37479) );
  NOR2X1 U31996 ( .A(n37480), .B(reg_B[118]), .Y(n37312) );
  NAND2X1 U31997 ( .A(n37481), .B(n37482), .Y(n37461) );
  AOI22X1 U31998 ( .A(n36315), .B(n36774), .C(n36442), .D(n37007), .Y(n37482)
         );
  OAI21X1 U31999 ( .A(n25469), .B(n36318), .C(n37483), .Y(n36774) );
  AOI22X1 U32000 ( .A(n36685), .B(reg_A[100]), .C(n36338), .D(reg_A[116]), .Y(
        n37483) );
  AOI22X1 U32001 ( .A(n36649), .B(n37307), .C(n36280), .D(n37484), .Y(n37481)
         );
  INVX1 U32002 ( .A(n37281), .Y(n37477) );
  NOR2X1 U32003 ( .A(n25523), .B(reg_B[117]), .Y(n37281) );
  NAND3X1 U32004 ( .A(n37485), .B(n37486), .C(n37487), .Y(n37468) );
  NOR2X1 U32005 ( .A(n37488), .B(n37489), .Y(n37487) );
  OAI22X1 U32006 ( .A(n27971), .B(n25321), .C(n25295), .D(n25494), .Y(n37489)
         );
  OAI22X1 U32007 ( .A(n25297), .B(n25490), .C(n27511), .D(n25493), .Y(n37488)
         );
  INVX1 U32008 ( .A(n29030), .Y(n25297) );
  OAI21X1 U32009 ( .A(n37490), .B(n37491), .C(n27358), .Y(n37486) );
  OAI21X1 U32010 ( .A(n25337), .B(n27442), .C(n37492), .Y(n37491) );
  OAI21X1 U32011 ( .A(n37493), .B(n37494), .C(n25044), .Y(n37492) );
  OAI22X1 U32012 ( .A(n27454), .B(n37450), .C(n27455), .D(n37495), .Y(n37494)
         );
  NOR2X1 U32013 ( .A(reg_B[4]), .B(n37444), .Y(n37493) );
  OAI21X1 U32014 ( .A(n37496), .B(n26030), .C(n37497), .Y(n37444) );
  AOI22X1 U32015 ( .A(n25025), .B(n37350), .C(n26032), .D(n36800), .Y(n37497)
         );
  OR2X1 U32016 ( .A(n37498), .B(n37499), .Y(n36800) );
  OAI22X1 U32017 ( .A(reg_A[116]), .B(n26036), .C(reg_A[108]), .D(n25058), .Y(
        n37499) );
  OAI21X1 U32018 ( .A(reg_A[100]), .B(n25055), .C(n36952), .Y(n37498) );
  OAI22X1 U32019 ( .A(n27449), .B(n36962), .C(n25476), .D(n27448), .Y(n37490)
         );
  NAND2X1 U32020 ( .A(reg_B[2]), .B(n25029), .Y(n27448) );
  NAND2X1 U32021 ( .A(n37500), .B(n37501), .Y(n36962) );
  AOI22X1 U32022 ( .A(n26601), .B(n25771), .C(n26602), .D(n25483), .Y(n37501)
         );
  AOI22X1 U32023 ( .A(n27012), .B(n25337), .C(n26597), .D(n25335), .Y(n37500)
         );
  NAND2X1 U32024 ( .A(n25029), .B(n26452), .Y(n27449) );
  AOI22X1 U32025 ( .A(reg_A[117]), .B(n25282), .C(n25372), .D(n37502), .Y(
        n37485) );
  NAND3X1 U32026 ( .A(n37503), .B(n37504), .C(n37505), .Y(n37502) );
  NOR2X1 U32027 ( .A(n37506), .B(n37507), .Y(n37505) );
  OAI22X1 U32028 ( .A(n36626), .B(n37392), .C(n37472), .D(n37235), .Y(n37507)
         );
  AOI22X1 U32029 ( .A(reg_A[116]), .B(n25793), .C(reg_A[114]), .D(n25399), .Y(
        n36626) );
  OAI21X1 U32030 ( .A(n37229), .B(n37508), .C(n37509), .Y(n37506) );
  AOI21X1 U32031 ( .A(n37510), .B(n37511), .C(n37512), .Y(n37509) );
  OAI21X1 U32032 ( .A(n37513), .B(n36172), .C(n37283), .Y(n37511) );
  MUX2X1 U32033 ( .B(n37514), .A(n37515), .S(reg_B[126]), .Y(n37508) );
  AOI22X1 U32034 ( .A(n37372), .B(n37226), .C(n37516), .D(reg_A[114]), .Y(
        n37504) );
  INVX1 U32035 ( .A(n37517), .Y(n37372) );
  OAI21X1 U32036 ( .A(n37518), .B(n25428), .C(n37519), .Y(n37517) );
  AOI22X1 U32037 ( .A(n36315), .B(n36821), .C(n36649), .D(n37270), .Y(n37519)
         );
  OR2X1 U32038 ( .A(n37520), .B(n37521), .Y(n36821) );
  OAI22X1 U32039 ( .A(reg_A[108]), .B(n36318), .C(reg_A[116]), .D(n36668), .Y(
        n37521) );
  OAI21X1 U32040 ( .A(reg_A[100]), .B(n36957), .C(n36958), .Y(n37520) );
  AOI22X1 U32041 ( .A(n37522), .B(reg_A[116]), .C(n37523), .D(reg_A[112]), .Y(
        n37503) );
  NOR2X1 U32042 ( .A(n37524), .B(n37525), .Y(n37466) );
  OAI21X1 U32043 ( .A(n25360), .B(n36140), .C(n37526), .Y(n37525) );
  AOI22X1 U32044 ( .A(reg_A[116]), .B(n31520), .C(reg_A[118]), .D(n25364), .Y(
        n37526) );
  NAND2X1 U32045 ( .A(n32946), .B(n35066), .Y(n31520) );
  INVX1 U32046 ( .A(n27622), .Y(n25360) );
  NAND3X1 U32047 ( .A(n37527), .B(n37528), .C(n37529), .Y(n37524) );
  AOI22X1 U32048 ( .A(n37389), .B(n37530), .C(reg_A[112]), .D(n31529), .Y(
        n37529) );
  OAI21X1 U32049 ( .A(n27443), .B(n26864), .C(n27431), .Y(n31529) );
  NAND2X1 U32050 ( .A(n26045), .B(n27242), .Y(n27431) );
  INVX1 U32051 ( .A(n37531), .Y(n37389) );
  NAND3X1 U32052 ( .A(n37390), .B(n36172), .C(n26267), .Y(n37528) );
  OAI22X1 U32053 ( .A(reg_B[126]), .B(n37240), .C(n25771), .D(n37380), .Y(
        n37390) );
  INVX1 U32054 ( .A(n37532), .Y(n37240) );
  OAI21X1 U32055 ( .A(n36236), .B(n25337), .C(n37283), .Y(n37532) );
  NAND2X1 U32056 ( .A(n36355), .B(reg_A[112]), .Y(n37283) );
  OAI21X1 U32057 ( .A(n37533), .B(n37534), .C(n25840), .Y(n37527) );
  NAND3X1 U32058 ( .A(n37535), .B(n37536), .C(n37537), .Y(n37534) );
  NOR2X1 U32059 ( .A(n37538), .B(n37539), .Y(n37537) );
  OAI22X1 U32060 ( .A(n25043), .B(n25337), .C(n25039), .D(n25448), .Y(n37539)
         );
  OAI21X1 U32061 ( .A(n25064), .B(n25298), .C(n37540), .Y(n37538) );
  AOI22X1 U32062 ( .A(reg_A[102]), .B(n25234), .C(reg_A[101]), .D(n25235), .Y(
        n37540) );
  AOI21X1 U32063 ( .A(reg_A[108]), .B(n25124), .C(n37541), .Y(n37536) );
  OAI22X1 U32064 ( .A(n25037), .B(n25470), .C(n25028), .D(n25452), .Y(n37541)
         );
  AOI22X1 U32065 ( .A(reg_A[105]), .B(n25222), .C(reg_A[106]), .D(n25637), .Y(
        n37535) );
  NAND3X1 U32066 ( .A(n37542), .B(n37543), .C(n37544), .Y(n37533) );
  NOR2X1 U32067 ( .A(n37545), .B(n37546), .Y(n37544) );
  OAI21X1 U32068 ( .A(n25042), .B(n25335), .C(n37547), .Y(n37546) );
  AOI22X1 U32069 ( .A(reg_A[98]), .B(n25241), .C(reg_A[96]), .D(n25339), .Y(
        n37547) );
  OAI21X1 U32070 ( .A(n25038), .B(n25287), .C(n37548), .Y(n37545) );
  AOI22X1 U32071 ( .A(reg_A[99]), .B(n25246), .C(reg_A[100]), .D(n25247), .Y(
        n37548) );
  AOI21X1 U32072 ( .A(reg_A[110]), .B(n25253), .C(n37549), .Y(n37543) );
  OAI22X1 U32073 ( .A(n25040), .B(n25771), .C(n25041), .D(n25483), .Y(n37549)
         );
  AOI22X1 U32074 ( .A(reg_A[109]), .B(n25628), .C(reg_A[112]), .D(n25067), .Y(
        n37542) );
  NOR2X1 U32075 ( .A(n37550), .B(n37551), .Y(n37465) );
  OAI21X1 U32076 ( .A(n27512), .B(n25323), .C(n37552), .Y(n37551) );
  AOI22X1 U32077 ( .A(reg_A[127]), .B(n25300), .C(reg_A[125]), .D(n25301), .Y(
        n37552) );
  NAND2X1 U32078 ( .A(n37553), .B(n37554), .Y(n37550) );
  AOI22X1 U32079 ( .A(reg_A[113]), .B(n27396), .C(reg_A[114]), .D(n27397), .Y(
        n37554) );
  OAI21X1 U32080 ( .A(n31658), .B(n25437), .C(n35473), .Y(n27397) );
  OAI21X1 U32081 ( .A(n31658), .B(n30437), .C(n27587), .Y(n27396) );
  AOI22X1 U32082 ( .A(reg_A[115]), .B(n27513), .C(reg_A[126]), .D(n25299), .Y(
        n37553) );
  INVX1 U32083 ( .A(n27394), .Y(n27513) );
  AOI21X1 U32084 ( .A(n27358), .B(n32188), .C(n27770), .Y(n27394) );
  INVX1 U32085 ( .A(n28303), .Y(n32188) );
  NAND3X1 U32086 ( .A(n37555), .B(n37556), .C(n37557), .Y(result[115]) );
  NOR2X1 U32087 ( .A(n37558), .B(n37559), .Y(n37557) );
  NAND3X1 U32088 ( .A(n37560), .B(n37561), .C(n37562), .Y(n37559) );
  AOI21X1 U32089 ( .A(n26045), .B(n37563), .C(n37564), .Y(n37562) );
  OAI21X1 U32090 ( .A(n32946), .B(n25335), .C(n37565), .Y(n37564) );
  OAI21X1 U32091 ( .A(n37563), .B(n37566), .C(n27358), .Y(n37565) );
  OAI21X1 U32092 ( .A(n37567), .B(n25476), .C(n37568), .Y(n37566) );
  OAI21X1 U32093 ( .A(n37569), .B(n37570), .C(n25044), .Y(n37568) );
  OAI22X1 U32094 ( .A(n27454), .B(n37571), .C(n26599), .D(n37450), .Y(n37570)
         );
  OAI21X1 U32095 ( .A(reg_B[2]), .B(n37152), .C(n37572), .Y(n37450) );
  AOI21X1 U32096 ( .A(n27570), .B(n37573), .C(n37574), .Y(n37572) );
  NOR2X1 U32097 ( .A(n37575), .B(n37576), .Y(n37152) );
  OAI22X1 U32098 ( .A(reg_A[115]), .B(n26036), .C(reg_A[107]), .D(n25058), .Y(
        n37576) );
  OAI21X1 U32099 ( .A(reg_A[99]), .B(n25055), .C(n36952), .Y(n37575) );
  OAI21X1 U32100 ( .A(n27575), .B(n37495), .C(n37577), .Y(n37569) );
  AOI22X1 U32101 ( .A(n37578), .B(n27577), .C(n27579), .D(reg_A[96]), .Y(
        n37577) );
  NOR2X1 U32102 ( .A(n27455), .B(n27677), .Y(n27579) );
  NOR2X1 U32103 ( .A(n27455), .B(reg_B[0]), .Y(n27577) );
  AOI21X1 U32104 ( .A(n25604), .B(n32939), .C(n35346), .Y(n37567) );
  OAI21X1 U32105 ( .A(n33395), .B(n26999), .C(n35476), .Y(n35346) );
  OAI21X1 U32106 ( .A(n25204), .B(n25335), .C(n37579), .Y(n37563) );
  AOI22X1 U32107 ( .A(reg_A[114]), .B(n25441), .C(reg_A[113]), .D(n27243), .Y(
        n37579) );
  MUX2X1 U32108 ( .B(n37580), .A(n37581), .S(reg_B[127]), .Y(n37561) );
  NOR2X1 U32109 ( .A(n37377), .B(n37513), .Y(n37580) );
  INVX1 U32110 ( .A(n37530), .Y(n37513) );
  OAI21X1 U32111 ( .A(n25483), .B(n37380), .C(n37582), .Y(n37530) );
  NAND3X1 U32112 ( .A(n36356), .B(n25428), .C(reg_A[115]), .Y(n37582) );
  AND2X1 U32113 ( .A(n25023), .B(n37583), .Y(n37377) );
  AOI22X1 U32114 ( .A(n25277), .B(n37475), .C(n37299), .D(n37584), .Y(n37560)
         );
  INVX1 U32115 ( .A(n37459), .Y(n37299) );
  NAND2X1 U32116 ( .A(n37585), .B(n37586), .Y(n37475) );
  AOI22X1 U32117 ( .A(n36315), .B(n36901), .C(n36442), .D(n37233), .Y(n37586)
         );
  OAI21X1 U32118 ( .A(n25470), .B(n36318), .C(n37587), .Y(n36901) );
  AOI22X1 U32119 ( .A(n36685), .B(reg_A[99]), .C(n36338), .D(reg_A[115]), .Y(
        n37587) );
  AOI22X1 U32120 ( .A(n36649), .B(n37410), .C(n36280), .D(n37588), .Y(n37585)
         );
  NAND3X1 U32121 ( .A(n37589), .B(n37590), .C(n37591), .Y(n37558) );
  AOI21X1 U32122 ( .A(reg_A[116]), .B(n25282), .C(n37592), .Y(n37591) );
  OAI22X1 U32123 ( .A(n27971), .B(n25494), .C(n25295), .D(n25490), .Y(n37592)
         );
  INVX1 U32124 ( .A(n25293), .Y(n27971) );
  OAI21X1 U32125 ( .A(n25042), .B(n26990), .C(n26781), .Y(n25282) );
  INVX1 U32126 ( .A(n28923), .Y(n26781) );
  AOI22X1 U32127 ( .A(reg_A[126]), .B(n25300), .C(reg_A[124]), .D(n25301), .Y(
        n37590) );
  OAI22X1 U32128 ( .A(n25037), .B(n26990), .C(n27253), .D(n27152), .Y(n25301)
         );
  OAI22X1 U32129 ( .A(n25473), .B(n26990), .C(n29558), .D(n27152), .Y(n25300)
         );
  AOI22X1 U32130 ( .A(reg_A[123]), .B(n25302), .C(reg_A[120]), .D(n29030), .Y(
        n37589) );
  AND2X1 U32131 ( .A(n37593), .B(n37594), .Y(n37556) );
  NOR2X1 U32132 ( .A(n37595), .B(n37596), .Y(n37594) );
  OAI21X1 U32133 ( .A(n37472), .B(n37597), .C(n37598), .Y(n37596) );
  OAI21X1 U32134 ( .A(n37599), .B(n37600), .C(n25840), .Y(n37598) );
  NAND3X1 U32135 ( .A(n37601), .B(n37602), .C(n37603), .Y(n37600) );
  NOR2X1 U32136 ( .A(n37604), .B(n37605), .Y(n37603) );
  OAI22X1 U32137 ( .A(n25043), .B(n25335), .C(n25039), .D(n25361), .Y(n37605)
         );
  OAI21X1 U32138 ( .A(n25064), .B(n25448), .C(n37606), .Y(n37604) );
  AOI22X1 U32139 ( .A(reg_A[101]), .B(n25234), .C(reg_A[100]), .D(n25235), .Y(
        n37606) );
  AOI21X1 U32140 ( .A(reg_A[107]), .B(n25124), .C(n37607), .Y(n37602) );
  OAI22X1 U32141 ( .A(n25037), .B(n25468), .C(n26703), .D(n25450), .Y(n37607)
         );
  AOI22X1 U32142 ( .A(reg_A[104]), .B(n25222), .C(reg_A[105]), .D(n25637), .Y(
        n37601) );
  NAND3X1 U32143 ( .A(n37608), .B(n37609), .C(n37610), .Y(n37599) );
  NOR2X1 U32144 ( .A(n37611), .B(n37612), .Y(n37610) );
  OAI22X1 U32145 ( .A(n25042), .B(n25771), .C(n25331), .D(n25287), .Y(n37612)
         );
  OAI21X1 U32146 ( .A(n25038), .B(n25424), .C(n37613), .Y(n37611) );
  AOI22X1 U32147 ( .A(reg_A[98]), .B(n25246), .C(reg_A[99]), .D(n25247), .Y(
        n37613) );
  AOI21X1 U32148 ( .A(reg_A[109]), .B(n25253), .C(n37614), .Y(n37609) );
  OAI22X1 U32149 ( .A(n25040), .B(n25483), .C(n25041), .D(n25476), .Y(n37614)
         );
  AOI22X1 U32150 ( .A(reg_A[108]), .B(n25628), .C(reg_A[111]), .D(n25066), .Y(
        n37608) );
  AOI21X1 U32151 ( .A(n26504), .B(n37615), .C(n37309), .Y(n37597) );
  INVX1 U32152 ( .A(n37616), .Y(n37309) );
  AOI22X1 U32153 ( .A(reg_A[115]), .B(n37169), .C(reg_A[113]), .D(n37383), .Y(
        n37472) );
  OAI21X1 U32154 ( .A(n25771), .B(n37617), .C(n37379), .Y(n37595) );
  NAND2X1 U32155 ( .A(n25372), .B(n37618), .Y(n37617) );
  AOI21X1 U32156 ( .A(n25932), .B(n37619), .C(n37620), .Y(n37593) );
  OAI22X1 U32157 ( .A(n37621), .B(n25476), .C(n37622), .D(n37531), .Y(n37620)
         );
  NAND2X1 U32158 ( .A(reg_B[127]), .B(n26267), .Y(n37531) );
  AOI21X1 U32159 ( .A(n26504), .B(n37623), .C(n37624), .Y(n37621) );
  OAI21X1 U32160 ( .A(n36247), .B(n37583), .C(n27587), .Y(n37624) );
  NAND2X1 U32161 ( .A(n26045), .B(n27241), .Y(n27587) );
  OAI21X1 U32162 ( .A(n37163), .B(n37615), .C(n37480), .Y(n37623) );
  NAND2X1 U32163 ( .A(n37625), .B(n37626), .Y(n37619) );
  AOI22X1 U32164 ( .A(n25355), .B(n37627), .C(n37514), .D(n25793), .Y(n37626)
         );
  INVX1 U32165 ( .A(n37363), .Y(n37514) );
  OAI21X1 U32166 ( .A(reg_B[125]), .B(n36867), .C(n37628), .Y(n37363) );
  AOI21X1 U32167 ( .A(n37629), .B(n36179), .C(n37630), .Y(n37628) );
  INVX1 U32168 ( .A(n37631), .Y(n36179) );
  NOR2X1 U32169 ( .A(n37632), .B(n37633), .Y(n36867) );
  OAI22X1 U32170 ( .A(reg_A[107]), .B(n36318), .C(reg_A[115]), .D(n36668), .Y(
        n37633) );
  OAI21X1 U32171 ( .A(reg_A[99]), .B(n36957), .C(n36958), .Y(n37632) );
  OAI21X1 U32172 ( .A(reg_B[123]), .B(n37634), .C(n37635), .Y(n37627) );
  AOI22X1 U32173 ( .A(n37518), .B(n25700), .C(n37515), .D(n25399), .Y(n37625)
         );
  INVX1 U32174 ( .A(n37636), .Y(n37515) );
  INVX1 U32175 ( .A(n37637), .Y(n37518) );
  NOR2X1 U32176 ( .A(n37638), .B(n37639), .Y(n37555) );
  OAI21X1 U32177 ( .A(n27620), .B(n25317), .C(n37640), .Y(n37639) );
  AOI22X1 U32178 ( .A(reg_A[117]), .B(n25364), .C(reg_A[118]), .D(n27622), .Y(
        n37640) );
  NAND2X1 U32179 ( .A(n27968), .B(n25718), .Y(n27622) );
  NAND2X1 U32180 ( .A(n27938), .B(n25717), .Y(n25364) );
  INVX1 U32181 ( .A(n25299), .Y(n27620) );
  OAI22X1 U32182 ( .A(n25036), .B(n26990), .C(n31398), .D(n27152), .Y(n25299)
         );
  OR2X1 U32183 ( .A(n37641), .B(n37642), .Y(n37638) );
  OAI22X1 U32184 ( .A(n27582), .B(n25497), .C(n37643), .D(n37301), .Y(n37642)
         );
  INVX1 U32185 ( .A(n25363), .Y(n27582) );
  OAI22X1 U32186 ( .A(n25064), .B(n26990), .C(n25738), .D(n27152), .Y(n25363)
         );
  OAI21X1 U32187 ( .A(n32909), .B(n36140), .C(n37644), .Y(n37641) );
  OAI21X1 U32188 ( .A(n37645), .B(n37646), .C(n25382), .Y(n37644) );
  OAI21X1 U32189 ( .A(n25337), .B(n37647), .C(n37648), .Y(n37646) );
  AOI22X1 U32190 ( .A(n37516), .B(reg_A[117]), .C(n37522), .D(reg_A[115]), .Y(
        n37648) );
  INVX1 U32191 ( .A(n37183), .Y(n37522) );
  OAI21X1 U32192 ( .A(n25333), .B(n37649), .C(n37650), .Y(n37645) );
  AOI22X1 U32193 ( .A(n37651), .B(n37166), .C(n37652), .D(n25410), .Y(n37650)
         );
  OAI21X1 U32194 ( .A(n37653), .B(n36247), .C(n37654), .Y(n25410) );
  AOI22X1 U32195 ( .A(reg_B[124]), .B(n36666), .C(n36356), .D(n37655), .Y(
        n37654) );
  INVX1 U32196 ( .A(n37656), .Y(n37166) );
  NOR2X1 U32197 ( .A(n36140), .B(n37244), .Y(n37651) );
  INVX1 U32198 ( .A(n25368), .Y(n32909) );
  NAND2X1 U32199 ( .A(n27511), .B(n32818), .Y(n25368) );
  INVX1 U32200 ( .A(n29029), .Y(n27511) );
  NAND3X1 U32201 ( .A(n37657), .B(n37658), .C(n37659), .Y(result[114]) );
  NOR2X1 U32202 ( .A(n37660), .B(n37661), .Y(n37659) );
  OR2X1 U32203 ( .A(n37662), .B(n37663), .Y(n37661) );
  OAI21X1 U32204 ( .A(n37664), .B(n25337), .C(n37665), .Y(n37663) );
  OAI21X1 U32205 ( .A(n37666), .B(n37667), .C(reg_A[112]), .Y(n37665) );
  OAI22X1 U32206 ( .A(n31658), .B(n35476), .C(n37169), .D(n25342), .Y(n37667)
         );
  NAND2X1 U32207 ( .A(n37668), .B(n35473), .Y(n37666) );
  NAND2X1 U32208 ( .A(n26045), .B(n27243), .Y(n35473) );
  OAI21X1 U32209 ( .A(n30427), .B(n30910), .C(n35474), .Y(n37668) );
  OAI21X1 U32210 ( .A(n37669), .B(n25087), .C(n37670), .Y(n37662) );
  OAI21X1 U32211 ( .A(n37671), .B(n37672), .C(reg_A[113]), .Y(n37670) );
  OAI21X1 U32212 ( .A(n37673), .B(n25517), .C(n31718), .Y(n37672) );
  NAND2X1 U32213 ( .A(n27358), .B(n25441), .Y(n31718) );
  INVX1 U32214 ( .A(n37618), .Y(n37673) );
  OAI21X1 U32215 ( .A(n25568), .B(n37392), .C(n37647), .Y(n37618) );
  AOI21X1 U32216 ( .A(n37674), .B(reg_A[115]), .C(n37675), .Y(n37669) );
  OAI21X1 U32217 ( .A(n25550), .B(n37676), .C(n37677), .Y(n37675) );
  NAND3X1 U32218 ( .A(n37678), .B(n37163), .C(n37523), .Y(n37677) );
  INVX1 U32219 ( .A(n37652), .Y(n37676) );
  AND2X1 U32220 ( .A(n37679), .B(n37680), .Y(n25550) );
  AOI22X1 U32221 ( .A(n36240), .B(n36362), .C(n36356), .D(n37681), .Y(n37680)
         );
  AOI22X1 U32222 ( .A(n36241), .B(n36790), .C(n36355), .D(n37682), .Y(n37679)
         );
  NAND3X1 U32223 ( .A(n37683), .B(n37684), .C(n37685), .Y(n37660) );
  AOI21X1 U32224 ( .A(n37686), .B(n26267), .C(n37687), .Y(n37685) );
  NAND2X1 U32225 ( .A(n37379), .B(n37688), .Y(n37687) );
  NAND2X1 U32226 ( .A(n37512), .B(n25372), .Y(n37379) );
  INVX1 U32227 ( .A(n37689), .Y(n37512) );
  NOR2X1 U32228 ( .A(reg_B[127]), .B(n37622), .Y(n37686) );
  INVX1 U32229 ( .A(n37690), .Y(n37622) );
  OAI21X1 U32230 ( .A(n25476), .B(n37380), .C(n37691), .Y(n37690) );
  NAND3X1 U32231 ( .A(n36356), .B(n25428), .C(reg_A[114]), .Y(n37691) );
  NAND2X1 U32232 ( .A(reg_B[126]), .B(n36356), .Y(n37380) );
  OAI21X1 U32233 ( .A(n37692), .B(n37693), .C(n25840), .Y(n37684) );
  NAND3X1 U32234 ( .A(n37694), .B(n37695), .C(n37696), .Y(n37693) );
  NOR2X1 U32235 ( .A(n37697), .B(n37698), .Y(n37696) );
  OAI22X1 U32236 ( .A(n25035), .B(n25436), .C(n25036), .D(n25298), .Y(n37698)
         );
  OAI21X1 U32237 ( .A(n25027), .B(n25448), .C(n37699), .Y(n37697) );
  AOI22X1 U32238 ( .A(reg_A[105]), .B(n25629), .C(reg_A[106]), .D(n25124), .Y(
        n37699) );
  AOI22X1 U32239 ( .A(reg_A[99]), .B(n25235), .C(reg_A[102]), .D(n25635), .Y(
        n37695) );
  AOI22X1 U32240 ( .A(reg_A[101]), .B(n25325), .C(reg_A[114]), .D(n25125), .Y(
        n37694) );
  NAND3X1 U32241 ( .A(n37700), .B(n37701), .C(n37702), .Y(n37692) );
  NOR2X1 U32242 ( .A(n37703), .B(n37704), .Y(n37702) );
  OAI22X1 U32243 ( .A(n25041), .B(n25452), .C(n25042), .D(n25483), .Y(n37704)
         );
  OAI21X1 U32244 ( .A(n25051), .B(n25424), .C(n37705), .Y(n37703) );
  AOI22X1 U32245 ( .A(reg_A[97]), .B(n25246), .C(reg_A[98]), .D(n25247), .Y(
        n37705) );
  AOI21X1 U32246 ( .A(reg_A[107]), .B(n25628), .C(n37706), .Y(n37701) );
  OAI22X1 U32247 ( .A(n25033), .B(n25469), .C(n25040), .D(n25476), .Y(n37706)
         );
  AOI22X1 U32248 ( .A(reg_A[110]), .B(n25073), .C(reg_A[109]), .D(n25123), .Y(
        n37700) );
  OAI21X1 U32249 ( .A(n27687), .B(n37707), .C(reg_A[114]), .Y(n37683) );
  OAI21X1 U32250 ( .A(n25204), .B(n31658), .C(n35066), .Y(n27687) );
  NOR2X1 U32251 ( .A(n37708), .B(n37709), .Y(n37658) );
  OAI22X1 U32252 ( .A(n37710), .B(n37616), .C(n37643), .D(n37303), .Y(n37709)
         );
  AND2X1 U32253 ( .A(n37711), .B(n37712), .Y(n37643) );
  AOI22X1 U32254 ( .A(n36315), .B(n37007), .C(n36442), .D(n37307), .Y(n37712)
         );
  OAI21X1 U32255 ( .A(n36318), .B(n25468), .C(n37713), .Y(n37007) );
  AOI22X1 U32256 ( .A(n36685), .B(reg_A[98]), .C(n36338), .D(reg_A[114]), .Y(
        n37713) );
  AOI22X1 U32257 ( .A(n36649), .B(n37484), .C(n36280), .D(n37714), .Y(n37711)
         );
  INVX1 U32258 ( .A(n37584), .Y(n37710) );
  OAI22X1 U32259 ( .A(n25771), .B(n37462), .C(n25476), .D(n37311), .Y(n37584)
         );
  OAI21X1 U32260 ( .A(n36140), .B(n25652), .C(n37715), .Y(n37708) );
  AOI22X1 U32261 ( .A(reg_A[117]), .B(n37716), .C(n25508), .D(reg_A[118]), .Y(
        n37715) );
  NOR2X1 U32262 ( .A(n37717), .B(n37718), .Y(n37657) );
  OAI21X1 U32263 ( .A(n37719), .B(n37301), .C(n37720), .Y(n37718) );
  OAI21X1 U32264 ( .A(n37721), .B(n37722), .C(n25932), .Y(n37720) );
  OAI22X1 U32265 ( .A(n25568), .B(n37636), .C(n25397), .D(n37637), .Y(n37722)
         );
  OAI21X1 U32266 ( .A(reg_B[125]), .B(n37271), .C(n37723), .Y(n37637) );
  AOI21X1 U32267 ( .A(n37629), .B(n36337), .C(n37630), .Y(n37723) );
  NOR2X1 U32268 ( .A(n37724), .B(n37725), .Y(n37271) );
  OAI22X1 U32269 ( .A(reg_A[106]), .B(n36318), .C(reg_A[114]), .D(n36668), .Y(
        n37725) );
  OAI21X1 U32270 ( .A(reg_A[98]), .B(n36957), .C(n36958), .Y(n37724) );
  OAI21X1 U32271 ( .A(n36136), .B(n37726), .C(n37727), .Y(n37721) );
  OAI21X1 U32272 ( .A(n37728), .B(n37006), .C(n25355), .Y(n37727) );
  NOR2X1 U32273 ( .A(reg_B[123]), .B(n37729), .Y(n37728) );
  MUX2X1 U32274 ( .B(n37730), .A(n37731), .S(reg_B[125]), .Y(n37726) );
  OAI21X1 U32275 ( .A(reg_B[123]), .B(n36612), .C(n37635), .Y(n37731) );
  INVX1 U32276 ( .A(n37270), .Y(n37730) );
  OAI21X1 U32277 ( .A(reg_A[96]), .B(n25551), .C(n37732), .Y(n37270) );
  AOI22X1 U32278 ( .A(n36338), .B(n25476), .C(n36686), .D(n25298), .Y(n37732)
         );
  OAI21X1 U32279 ( .A(n37733), .B(n37734), .C(n37735), .Y(n37717) );
  OAI21X1 U32280 ( .A(n37736), .B(n37737), .C(n25203), .Y(n37735) );
  NAND3X1 U32281 ( .A(n37738), .B(n37739), .C(n37740), .Y(n37737) );
  AOI21X1 U32282 ( .A(reg_A[116]), .B(n27637), .C(n37741), .Y(n37740) );
  OAI22X1 U32283 ( .A(n25599), .B(n25332), .C(n25600), .D(n36140), .Y(n37741)
         );
  AOI22X1 U32284 ( .A(reg_A[114]), .B(n27639), .C(reg_A[115]), .D(n25617), .Y(
        n37739) );
  AOI22X1 U32285 ( .A(reg_A[118]), .B(n25650), .C(reg_A[120]), .D(n25651), .Y(
        n37738) );
  NAND3X1 U32286 ( .A(n37742), .B(n37743), .C(n37744), .Y(n37736) );
  AOI21X1 U32287 ( .A(reg_A[125]), .B(n27643), .C(n37745), .Y(n37744) );
  OAI22X1 U32288 ( .A(n27645), .B(n25323), .C(n27646), .D(n25321), .Y(n37745)
         );
  AOI21X1 U32289 ( .A(n25044), .B(n25629), .C(n25500), .Y(n27646) );
  AOI21X1 U32290 ( .A(n25097), .B(n25637), .C(n25439), .Y(n27645) );
  INVX1 U32291 ( .A(n28362), .Y(n25439) );
  OAI21X1 U32292 ( .A(n25403), .B(n25473), .C(n28363), .Y(n27643) );
  AOI22X1 U32293 ( .A(reg_A[126]), .B(n27647), .C(reg_A[127]), .D(n27648), .Y(
        n37743) );
  OAI21X1 U32294 ( .A(n25403), .B(n25231), .C(n25451), .Y(n27647) );
  AOI22X1 U32295 ( .A(reg_A[121]), .B(n27649), .C(reg_A[122]), .D(n27650), .Y(
        n37742) );
  OAI21X1 U32296 ( .A(n25403), .B(n25467), .C(n30444), .Y(n27650) );
  OAI21X1 U32297 ( .A(n25403), .B(n25129), .C(n30443), .Y(n27649) );
  NAND2X1 U32298 ( .A(n37746), .B(n27676), .Y(n37734) );
  AOI22X1 U32299 ( .A(n26597), .B(n37495), .C(n26009), .D(n37350), .Y(n37746)
         );
  OAI21X1 U32300 ( .A(reg_A[96]), .B(n27677), .C(n37747), .Y(n37350) );
  AOI22X1 U32301 ( .A(n26038), .B(n25298), .C(n26664), .D(n25476), .Y(n37747)
         );
  OAI21X1 U32302 ( .A(n37496), .B(n26599), .C(n37748), .Y(n37733) );
  AOI22X1 U32303 ( .A(n27680), .B(n25424), .C(n37749), .D(n27677), .Y(n37748)
         );
  OAI21X1 U32304 ( .A(n37750), .B(n25754), .C(n37751), .Y(n37749) );
  AOI22X1 U32305 ( .A(n26002), .B(n36731), .C(n26008), .D(n37573), .Y(n37751)
         );
  AOI21X1 U32306 ( .A(n27455), .B(n26208), .C(n27677), .Y(n27680) );
  INVX1 U32307 ( .A(n37571), .Y(n37496) );
  OAI21X1 U32308 ( .A(reg_B[2]), .B(n37349), .C(n37752), .Y(n37571) );
  AOI21X1 U32309 ( .A(n27570), .B(n36407), .C(n37574), .Y(n37752) );
  NOR2X1 U32310 ( .A(n37753), .B(n37754), .Y(n37349) );
  OAI22X1 U32311 ( .A(reg_A[114]), .B(n26036), .C(reg_A[106]), .D(n25058), .Y(
        n37754) );
  OAI21X1 U32312 ( .A(reg_A[98]), .B(n25055), .C(n36952), .Y(n37753) );
  OR2X1 U32313 ( .A(n37755), .B(n37756), .Y(result[113]) );
  NAND3X1 U32314 ( .A(n37757), .B(n37758), .C(n37759), .Y(n37756) );
  NOR2X1 U32315 ( .A(n37760), .B(n37761), .Y(n37759) );
  OAI21X1 U32316 ( .A(n37762), .B(n37301), .C(n37763), .Y(n37761) );
  OAI21X1 U32317 ( .A(n37764), .B(n37765), .C(n25372), .Y(n37763) );
  OAI21X1 U32318 ( .A(n37766), .B(n37229), .C(n37767), .Y(n37765) );
  OAI21X1 U32319 ( .A(n37768), .B(n37769), .C(n37226), .Y(n37767) );
  MUX2X1 U32320 ( .B(n37636), .A(n37635), .S(reg_B[126]), .Y(n37769) );
  OAI21X1 U32321 ( .A(reg_B[125]), .B(n37176), .C(n37770), .Y(n37636) );
  AOI21X1 U32322 ( .A(n37629), .B(n36458), .C(n37630), .Y(n37770) );
  INVX1 U32323 ( .A(n37771), .Y(n37630) );
  NAND3X1 U32324 ( .A(reg_B[125]), .B(n25424), .C(reg_B[123]), .Y(n37771) );
  INVX1 U32325 ( .A(n37772), .Y(n36458) );
  NOR2X1 U32326 ( .A(n36177), .B(reg_B[123]), .Y(n37629) );
  NOR2X1 U32327 ( .A(n37773), .B(n37774), .Y(n37176) );
  OAI22X1 U32328 ( .A(reg_A[105]), .B(n36318), .C(reg_A[113]), .D(n36668), .Y(
        n37774) );
  OAI21X1 U32329 ( .A(reg_A[97]), .B(n36957), .C(n36958), .Y(n37773) );
  NAND2X1 U32330 ( .A(n36684), .B(n25424), .Y(n36958) );
  NOR2X1 U32331 ( .A(n25551), .B(n36291), .Y(n36684) );
  NOR2X1 U32332 ( .A(reg_B[123]), .B(n37775), .Y(n37768) );
  AOI22X1 U32333 ( .A(n36648), .B(n36280), .C(n36442), .D(n37631), .Y(n37775)
         );
  AOI21X1 U32334 ( .A(n37776), .B(n25551), .C(n37006), .Y(n37766) );
  OAI21X1 U32335 ( .A(n25476), .B(n37777), .C(n37689), .Y(n37764) );
  NAND2X1 U32336 ( .A(n37510), .B(n37285), .Y(n37689) );
  NOR2X1 U32337 ( .A(n36291), .B(n25476), .Y(n37285) );
  NAND2X1 U32338 ( .A(n25029), .B(n37462), .Y(n37777) );
  INVX1 U32339 ( .A(n37778), .Y(n37762) );
  OAI21X1 U32340 ( .A(n37719), .B(n37303), .C(n37779), .Y(n37760) );
  OAI21X1 U32341 ( .A(n37780), .B(n37781), .C(n25203), .Y(n37779) );
  NAND3X1 U32342 ( .A(n37782), .B(n37783), .C(n37784), .Y(n37781) );
  AOI22X1 U32343 ( .A(reg_A[116]), .B(n27740), .C(reg_A[115]), .D(n27637), .Y(
        n37784) );
  OAI21X1 U32344 ( .A(n37785), .B(n37786), .C(n25044), .Y(n37783) );
  NAND2X1 U32345 ( .A(n37787), .B(n37788), .Y(n37786) );
  AOI22X1 U32346 ( .A(reg_A[123]), .B(n25637), .C(reg_A[127]), .D(n25234), .Y(
        n37788) );
  AOI22X1 U32347 ( .A(reg_A[125]), .B(n25635), .C(reg_A[126]), .D(n25325), .Y(
        n37787) );
  NAND2X1 U32348 ( .A(n37789), .B(n37790), .Y(n37785) );
  AOI22X1 U32349 ( .A(reg_A[120]), .B(n25628), .C(reg_A[122]), .D(n25629), .Y(
        n37790) );
  AOI22X1 U32350 ( .A(reg_A[121]), .B(n25124), .C(reg_A[124]), .D(n25222), .Y(
        n37789) );
  OAI21X1 U32351 ( .A(n37791), .B(n37792), .C(n25604), .Y(n37782) );
  NAND2X1 U32352 ( .A(n37793), .B(n37794), .Y(n37792) );
  AOI22X1 U32353 ( .A(reg_A[123]), .B(n25607), .C(reg_A[127]), .D(n25608), .Y(
        n37794) );
  AOI22X1 U32354 ( .A(reg_A[125]), .B(n25609), .C(reg_A[126]), .D(n25610), .Y(
        n37793) );
  NAND2X1 U32355 ( .A(n37795), .B(n37796), .Y(n37791) );
  AOI22X1 U32356 ( .A(reg_A[120]), .B(n25613), .C(reg_A[122]), .D(n25614), .Y(
        n37796) );
  AOI22X1 U32357 ( .A(reg_A[121]), .B(n25615), .C(reg_A[124]), .D(n25616), .Y(
        n37795) );
  OR2X1 U32358 ( .A(n37797), .B(n37798), .Y(n37780) );
  OAI22X1 U32359 ( .A(n25600), .B(n25333), .C(n27755), .D(n36140), .Y(n37798)
         );
  INVX1 U32360 ( .A(n25651), .Y(n27755) );
  OAI21X1 U32361 ( .A(n25403), .B(n25131), .C(n28311), .Y(n25651) );
  INVX1 U32362 ( .A(n30721), .Y(n25600) );
  OAI21X1 U32363 ( .A(n25403), .B(n26703), .C(n25449), .Y(n30721) );
  OAI21X1 U32364 ( .A(n27756), .B(n25332), .C(n37799), .Y(n37797) );
  AOI22X1 U32365 ( .A(reg_A[113]), .B(n27639), .C(reg_A[114]), .D(n25617), .Y(
        n37799) );
  NAND2X1 U32366 ( .A(n29467), .B(n30791), .Y(n25617) );
  INVX1 U32367 ( .A(n25619), .Y(n27639) );
  NOR2X1 U32368 ( .A(n29466), .B(n30792), .Y(n25619) );
  INVX1 U32369 ( .A(n25650), .Y(n27756) );
  AND2X1 U32370 ( .A(n37800), .B(n37801), .Y(n37719) );
  AOI22X1 U32371 ( .A(n36315), .B(n37233), .C(n36442), .D(n37410), .Y(n37801)
         );
  OAI21X1 U32372 ( .A(n36318), .B(n25296), .C(n37802), .Y(n37233) );
  AOI22X1 U32373 ( .A(n36685), .B(reg_A[97]), .C(n36338), .D(reg_A[113]), .Y(
        n37802) );
  AOI22X1 U32374 ( .A(n36649), .B(n37588), .C(n36280), .D(n37803), .Y(n37800)
         );
  AOI21X1 U32375 ( .A(reg_A[116]), .B(n37716), .C(n37804), .Y(n37758) );
  OAI21X1 U32376 ( .A(n37664), .B(n25335), .C(n37805), .Y(n37804) );
  OAI21X1 U32377 ( .A(n37806), .B(n37807), .C(reg_A[112]), .Y(n37805) );
  NAND2X1 U32378 ( .A(n37808), .B(n35229), .Y(n37807) );
  AOI22X1 U32379 ( .A(n25736), .B(n30910), .C(n26943), .D(n30427), .Y(n35229)
         );
  INVX1 U32380 ( .A(n37671), .Y(n37808) );
  OAI21X1 U32381 ( .A(n37462), .B(n37459), .C(n37809), .Y(n37671) );
  AOI21X1 U32382 ( .A(n37810), .B(n25700), .C(n27770), .Y(n37809) );
  NOR2X1 U32383 ( .A(n27523), .B(n27218), .Y(n27770) );
  NOR2X1 U32384 ( .A(n25023), .B(n36236), .Y(n37810) );
  NAND2X1 U32385 ( .A(reg_B[119]), .B(n26186), .Y(n37459) );
  OAI22X1 U32386 ( .A(n25031), .B(n37615), .C(n36172), .D(n37583), .Y(n37806)
         );
  NAND2X1 U32387 ( .A(n37510), .B(n25372), .Y(n37583) );
  AOI21X1 U32388 ( .A(n25382), .B(n37516), .C(n25506), .Y(n37664) );
  INVX1 U32389 ( .A(n29766), .Y(n25506) );
  NAND2X1 U32390 ( .A(n27388), .B(n25203), .Y(n29766) );
  INVX1 U32391 ( .A(n37224), .Y(n37516) );
  OAI21X1 U32392 ( .A(n25087), .B(n37649), .C(n29765), .Y(n37716) );
  NAND2X1 U32393 ( .A(n27386), .B(n25203), .Y(n29765) );
  INVX1 U32394 ( .A(n36451), .Y(n27386) );
  INVX1 U32395 ( .A(n37811), .Y(n37649) );
  AOI22X1 U32396 ( .A(n25508), .B(reg_A[117]), .C(n25509), .D(reg_A[118]), .Y(
        n37757) );
  INVX1 U32397 ( .A(n25652), .Y(n25509) );
  NAND2X1 U32398 ( .A(n30177), .B(n25203), .Y(n25652) );
  INVX1 U32399 ( .A(n30355), .Y(n30177) );
  INVX1 U32400 ( .A(n29782), .Y(n25508) );
  NAND2X1 U32401 ( .A(n30357), .B(n25203), .Y(n29782) );
  NAND3X1 U32402 ( .A(n37812), .B(n37813), .C(n37814), .Y(n37755) );
  NOR2X1 U32403 ( .A(n37815), .B(n37816), .Y(n37814) );
  OAI21X1 U32404 ( .A(n27820), .B(n36731), .C(n37817), .Y(n37816) );
  OAI21X1 U32405 ( .A(n37818), .B(n37819), .C(reg_A[113]), .Y(n37817) );
  OAI21X1 U32406 ( .A(n25204), .B(n25279), .C(n37820), .Y(n37819) );
  INVX1 U32407 ( .A(n37707), .Y(n37820) );
  OAI21X1 U32408 ( .A(n34089), .B(n37183), .C(n37821), .Y(n37707) );
  NAND3X1 U32409 ( .A(n25793), .B(n25372), .C(n37822), .Y(n37821) );
  INVX1 U32410 ( .A(n37392), .Y(n37822) );
  NAND2X1 U32411 ( .A(n37510), .B(n36356), .Y(n37392) );
  NOR2X1 U32412 ( .A(n37188), .B(n25415), .Y(n37510) );
  INVX1 U32413 ( .A(n31887), .Y(n34089) );
  NAND2X1 U32414 ( .A(n25517), .B(n25087), .Y(n31887) );
  INVX1 U32415 ( .A(n37823), .Y(n36731) );
  NAND2X1 U32416 ( .A(n27921), .B(n26010), .Y(n27820) );
  OAI21X1 U32417 ( .A(n37824), .B(n30951), .C(n37825), .Y(n37815) );
  AOI21X1 U32418 ( .A(n37826), .B(reg_A[96]), .C(n37581), .Y(n37825) );
  INVX1 U32419 ( .A(n37688), .Y(n37581) );
  NAND3X1 U32420 ( .A(n36961), .B(n25372), .C(n36906), .Y(n37688) );
  INVX1 U32421 ( .A(n37827), .Y(n36906) );
  NAND3X1 U32422 ( .A(reg_A[112]), .B(n36359), .C(n36235), .Y(n37827) );
  INVX1 U32423 ( .A(n36667), .Y(n36961) );
  NAND2X1 U32424 ( .A(n25604), .B(n36291), .Y(n36667) );
  AOI21X1 U32425 ( .A(n26012), .B(n25939), .C(n27677), .Y(n37826) );
  NAND2X1 U32426 ( .A(n26028), .B(reg_B[3]), .Y(n25939) );
  NOR2X1 U32427 ( .A(n37828), .B(n37829), .Y(n37824) );
  NAND3X1 U32428 ( .A(n37830), .B(n37831), .C(n37832), .Y(n37829) );
  NOR2X1 U32429 ( .A(n37833), .B(n37834), .Y(n37832) );
  OAI22X1 U32430 ( .A(n25035), .B(n25396), .C(n25036), .D(n25448), .Y(n37834)
         );
  OAI21X1 U32431 ( .A(n25027), .B(n25361), .C(n37835), .Y(n37833) );
  AOI22X1 U32432 ( .A(reg_A[104]), .B(n25629), .C(reg_A[105]), .D(n25124), .Y(
        n37835) );
  AOI22X1 U32433 ( .A(reg_A[98]), .B(n25235), .C(reg_A[101]), .D(n25635), .Y(
        n37831) );
  AOI22X1 U32434 ( .A(reg_A[100]), .B(n25325), .C(reg_A[113]), .D(n25125), .Y(
        n37830) );
  NAND3X1 U32435 ( .A(n37836), .B(n37837), .C(n37838), .Y(n37828) );
  NOR2X1 U32436 ( .A(n37839), .B(n37840), .Y(n37838) );
  OAI22X1 U32437 ( .A(n25040), .B(n25452), .C(n25041), .D(n25450), .Y(n37840)
         );
  OAI21X1 U32438 ( .A(n25042), .B(n25476), .C(n37841), .Y(n37839) );
  AOI22X1 U32439 ( .A(reg_A[96]), .B(n25246), .C(reg_A[97]), .D(n25247), .Y(
        n37841) );
  AOI22X1 U32440 ( .A(reg_A[107]), .B(n25253), .C(reg_A[106]), .D(n25628), .Y(
        n37837) );
  AOI22X1 U32441 ( .A(reg_A[109]), .B(n25074), .C(reg_A[108]), .D(n25123), .Y(
        n37836) );
  AOI21X1 U32442 ( .A(n36262), .B(n37842), .C(n37843), .Y(n37813) );
  OAI22X1 U32443 ( .A(n27825), .B(n37495), .C(n27821), .D(n37844), .Y(n37843)
         );
  NAND2X1 U32444 ( .A(n26260), .B(n27677), .Y(n27821) );
  INVX1 U32445 ( .A(n26012), .Y(n26260) );
  NAND2X1 U32446 ( .A(n27676), .B(reg_B[4]), .Y(n26012) );
  OAI21X1 U32447 ( .A(reg_B[2]), .B(n37449), .C(n37845), .Y(n37495) );
  AOI21X1 U32448 ( .A(n27570), .B(n36466), .C(n37574), .Y(n37845) );
  AND2X1 U32449 ( .A(n27828), .B(n25424), .Y(n37574) );
  NOR2X1 U32450 ( .A(n27677), .B(n26452), .Y(n27828) );
  NOR2X1 U32451 ( .A(n26452), .B(reg_B[0]), .Y(n27570) );
  NOR2X1 U32452 ( .A(n37846), .B(n37847), .Y(n37449) );
  OAI22X1 U32453 ( .A(reg_A[113]), .B(n26036), .C(reg_A[105]), .D(n25058), .Y(
        n37847) );
  NAND2X1 U32454 ( .A(reg_B[1]), .B(n27677), .Y(n26981) );
  OAI21X1 U32455 ( .A(reg_A[97]), .B(n25055), .C(n36952), .Y(n37846) );
  NAND2X1 U32456 ( .A(n26662), .B(n25424), .Y(n36952) );
  NOR2X1 U32457 ( .A(n26596), .B(n27677), .Y(n26662) );
  NAND2X1 U32458 ( .A(reg_B[0]), .B(n26596), .Y(n26982) );
  NAND2X1 U32459 ( .A(n27012), .B(n27676), .Y(n27825) );
  INVX1 U32460 ( .A(n27826), .Y(n37842) );
  NAND2X1 U32461 ( .A(n27921), .B(n26009), .Y(n27826) );
  AOI22X1 U32462 ( .A(n29779), .B(reg_A[119]), .C(n25382), .D(n37848), .Y(
        n37812) );
  OAI21X1 U32463 ( .A(n25771), .B(n37647), .C(n37849), .Y(n37848) );
  AOI22X1 U32464 ( .A(n37652), .B(n25688), .C(n37523), .D(n37457), .Y(n37849)
         );
  OAI21X1 U32465 ( .A(n25332), .B(n37656), .C(n37850), .Y(n37457) );
  MUX2X1 U32466 ( .B(n37851), .A(n37852), .S(reg_B[119]), .Y(n37850) );
  NOR2X1 U32467 ( .A(reg_B[118]), .B(n25333), .Y(n37852) );
  NOR2X1 U32468 ( .A(n36140), .B(n37163), .Y(n37851) );
  INVX1 U32469 ( .A(n37244), .Y(n37523) );
  NAND2X1 U32470 ( .A(n37853), .B(n37854), .Y(n25688) );
  AOI22X1 U32471 ( .A(n36240), .B(n36911), .C(n36356), .D(n37855), .Y(n37854)
         );
  AOI22X1 U32472 ( .A(n36241), .B(n36877), .C(n36355), .D(n37856), .Y(n37853)
         );
  INVX1 U32473 ( .A(n25702), .Y(n29779) );
  NAND2X1 U32474 ( .A(n30722), .B(n25203), .Y(n25702) );
  INVX1 U32475 ( .A(n30179), .Y(n30722) );
  OR2X1 U32476 ( .A(n37857), .B(n37858), .Y(result[112]) );
  NAND3X1 U32477 ( .A(n37859), .B(n37860), .C(n37861), .Y(n37858) );
  NOR2X1 U32478 ( .A(n37862), .B(n37863), .Y(n37861) );
  OAI22X1 U32479 ( .A(n25771), .B(n25717), .C(n25335), .D(n25718), .Y(n37863)
         );
  OAI21X1 U32480 ( .A(n25483), .B(n25719), .C(n37864), .Y(n37862) );
  AOI22X1 U32481 ( .A(n25277), .B(n37778), .C(n25275), .D(n37865), .Y(n37864)
         );
  OAI21X1 U32482 ( .A(n37866), .B(n36312), .C(n37867), .Y(n37778) );
  AOI22X1 U32483 ( .A(n36315), .B(n37307), .C(n37868), .D(reg_B[126]), .Y(
        n37867) );
  OAI21X1 U32484 ( .A(n36318), .B(n25298), .C(n37869), .Y(n37307) );
  AOI22X1 U32485 ( .A(n36685), .B(reg_A[96]), .C(n36338), .D(reg_A[112]), .Y(
        n37869) );
  AOI21X1 U32486 ( .A(reg_A[112]), .B(n37870), .C(n37871), .Y(n37860) );
  OAI21X1 U32487 ( .A(n37872), .B(n25726), .C(n37873), .Y(n37871) );
  OAI21X1 U32488 ( .A(n37874), .B(n37875), .C(n25382), .Y(n37873) );
  OAI22X1 U32489 ( .A(n37476), .B(n37244), .C(n25483), .D(n37647), .Y(n37875)
         );
  INVX1 U32490 ( .A(n37674), .Y(n37647) );
  NOR2X1 U32491 ( .A(n37235), .B(n37462), .Y(n37674) );
  NAND2X1 U32492 ( .A(reg_B[117]), .B(n25029), .Y(n37244) );
  INVX1 U32493 ( .A(n37876), .Y(n37476) );
  OAI21X1 U32494 ( .A(n25337), .B(n37656), .C(n37877), .Y(n37876) );
  MUX2X1 U32495 ( .B(n37878), .A(n37678), .S(reg_B[118]), .Y(n37877) );
  INVX1 U32496 ( .A(n37286), .Y(n37678) );
  MUX2X1 U32497 ( .B(reg_A[118]), .A(reg_A[119]), .S(reg_B[119]), .Y(n37286)
         );
  NOR2X1 U32498 ( .A(n25332), .B(n37615), .Y(n37878) );
  NAND2X1 U32499 ( .A(n37163), .B(n37615), .Y(n37656) );
  OAI21X1 U32500 ( .A(n25771), .B(n37224), .C(n37879), .Y(n37874) );
  AOI22X1 U32501 ( .A(n37652), .B(n25813), .C(n37811), .D(reg_A[115]), .Y(
        n37879) );
  NOR2X1 U32502 ( .A(n37235), .B(n37311), .Y(n37811) );
  NAND2X1 U32503 ( .A(reg_B[119]), .B(n25029), .Y(n37235) );
  NAND2X1 U32504 ( .A(n37880), .B(n37881), .Y(n25813) );
  AOI22X1 U32505 ( .A(n36240), .B(n36619), .C(n36356), .D(n37882), .Y(n37881)
         );
  AOI22X1 U32506 ( .A(n36241), .B(n37883), .C(n36355), .D(n37884), .Y(n37880)
         );
  OAI21X1 U32507 ( .A(reg_B[123]), .B(n25403), .C(n25415), .Y(n37652) );
  NAND3X1 U32508 ( .A(n25589), .B(n37615), .C(n37383), .Y(n37224) );
  INVX1 U32509 ( .A(n37311), .Y(n37383) );
  NAND2X1 U32510 ( .A(reg_B[118]), .B(n37480), .Y(n37311) );
  AOI21X1 U32511 ( .A(reg_A[117]), .B(n25751), .C(n37885), .Y(n37872) );
  OAI22X1 U32512 ( .A(n25753), .B(n36140), .C(n25754), .D(n25333), .Y(n37885)
         );
  NAND3X1 U32513 ( .A(n37886), .B(n25795), .C(n37887), .Y(n37870) );
  NOR2X1 U32514 ( .A(n37818), .B(n37888), .Y(n37887) );
  OAI21X1 U32515 ( .A(n25087), .B(n37183), .C(n37889), .Y(n37888) );
  INVX1 U32516 ( .A(n35639), .Y(n37889) );
  NAND3X1 U32517 ( .A(n29998), .B(n25031), .C(n35066), .Y(n35639) );
  NAND2X1 U32518 ( .A(n26045), .B(n25434), .Y(n35066) );
  NAND3X1 U32519 ( .A(n25589), .B(n37615), .C(n37169), .Y(n37183) );
  INVX1 U32520 ( .A(n37462), .Y(n37169) );
  OAI21X1 U32521 ( .A(n37462), .B(n37616), .C(n37890), .Y(n37818) );
  NAND3X1 U32522 ( .A(n36356), .B(n26267), .C(n25793), .Y(n37890) );
  NAND2X1 U32523 ( .A(n26186), .B(n37615), .Y(n37616) );
  INVX1 U32524 ( .A(reg_B[119]), .Y(n37615) );
  NOR2X1 U32525 ( .A(n30910), .B(n36286), .Y(n37886) );
  NOR2X1 U32526 ( .A(n37188), .B(n25032), .Y(n36286) );
  INVX1 U32527 ( .A(n36235), .Y(n37188) );
  NOR2X1 U32528 ( .A(n37891), .B(n37892), .Y(n36235) );
  NAND3X1 U32529 ( .A(n37893), .B(n37894), .C(n37895), .Y(n37892) );
  NOR2X1 U32530 ( .A(n37462), .B(n37896), .Y(n37895) );
  NAND2X1 U32531 ( .A(n25561), .B(n25522), .Y(n37896) );
  NAND2X1 U32532 ( .A(n37480), .B(n37163), .Y(n37462) );
  INVX1 U32533 ( .A(reg_B[118]), .Y(n37163) );
  INVX1 U32534 ( .A(reg_B[117]), .Y(n37480) );
  NOR2X1 U32535 ( .A(reg_B[114]), .B(reg_B[113]), .Y(n37894) );
  NOR2X1 U32536 ( .A(reg_B[112]), .B(n25591), .Y(n37893) );
  NAND3X1 U32537 ( .A(n37897), .B(n37898), .C(n37899), .Y(n37891) );
  NOR2X1 U32538 ( .A(reg_B[115]), .B(n37900), .Y(n37899) );
  OR2X1 U32539 ( .A(reg_B[119]), .B(reg_B[116]), .Y(n37900) );
  NOR2X1 U32540 ( .A(reg_B[123]), .B(reg_B[122]), .Y(n37898) );
  NOR2X1 U32541 ( .A(reg_B[121]), .B(reg_B[120]), .Y(n37897) );
  AOI22X1 U32542 ( .A(n32020), .B(reg_A[96]), .C(n25722), .D(reg_A[116]), .Y(
        n37859) );
  INVX1 U32543 ( .A(n32818), .Y(n25722) );
  NAND2X1 U32544 ( .A(n26928), .B(n26003), .Y(n32818) );
  INVX1 U32545 ( .A(n31636), .Y(n32020) );
  NAND3X1 U32546 ( .A(n37901), .B(n37902), .C(n37903), .Y(n37857) );
  NOR2X1 U32547 ( .A(n37904), .B(n37905), .Y(n37903) );
  OAI21X1 U32548 ( .A(reg_B[123]), .B(n37906), .C(n37907), .Y(n37905) );
  OAI21X1 U32549 ( .A(n37908), .B(n37909), .C(n25310), .Y(n37907) );
  NAND3X1 U32550 ( .A(n37910), .B(n37911), .C(n37912), .Y(n37909) );
  NOR2X1 U32551 ( .A(n37913), .B(n37914), .Y(n37912) );
  OAI22X1 U32552 ( .A(n25043), .B(n25476), .C(n25039), .D(n25317), .Y(n37914)
         );
  OAI22X1 U32553 ( .A(n25064), .B(n25323), .C(n25482), .D(n25497), .Y(n37913)
         );
  AOI22X1 U32554 ( .A(reg_A[120]), .B(n25124), .C(reg_A[123]), .D(n25222), .Y(
        n37911) );
  AOI22X1 U32555 ( .A(reg_A[122]), .B(n25637), .C(reg_A[126]), .D(n25234), .Y(
        n37910) );
  NAND3X1 U32556 ( .A(n37915), .B(n37916), .C(n37917), .Y(n37908) );
  NOR2X1 U32557 ( .A(n37918), .B(n37919), .Y(n37917) );
  OAI22X1 U32558 ( .A(n25033), .B(n25333), .C(n25040), .D(n25771), .Y(n37919)
         );
  OAI22X1 U32559 ( .A(n25041), .B(n25335), .C(n25784), .D(n25483), .Y(n37918)
         );
  AOI22X1 U32560 ( .A(reg_A[119]), .B(n25628), .C(reg_A[116]), .D(n25067), .Y(
        n37916) );
  AOI22X1 U32561 ( .A(reg_A[117]), .B(n25123), .C(reg_A[121]), .D(n25629), .Y(
        n37915) );
  AOI22X1 U32562 ( .A(n37920), .B(n37921), .C(n37776), .D(n36329), .Y(n37906)
         );
  AOI21X1 U32563 ( .A(n25428), .B(n37634), .C(n37922), .Y(n37776) );
  INVX1 U32564 ( .A(n37923), .Y(n37922) );
  AOI22X1 U32565 ( .A(n37924), .B(n36280), .C(n36442), .D(n36337), .Y(n37923)
         );
  MUX2X1 U32566 ( .B(reg_A[102]), .A(reg_A[110]), .S(n36291), .Y(n36337) );
  MUX2X1 U32567 ( .B(reg_A[106]), .A(reg_A[98]), .S(reg_B[124]), .Y(n37924) );
  OAI21X1 U32568 ( .A(reg_A[112]), .B(n36236), .C(n37925), .Y(n37634) );
  AOI22X1 U32569 ( .A(reg_B[125]), .B(n36612), .C(n36241), .D(n25298), .Y(
        n37925) );
  MUX2X1 U32570 ( .B(reg_A[100]), .A(reg_A[108]), .S(n36291), .Y(n36612) );
  INVX1 U32571 ( .A(n37729), .Y(n37921) );
  MUX2X1 U32572 ( .B(n37631), .A(n36648), .S(reg_B[125]), .Y(n37729) );
  MUX2X1 U32573 ( .B(n25470), .A(n25396), .S(reg_B[124]), .Y(n36648) );
  MUX2X1 U32574 ( .B(n25452), .A(n25448), .S(reg_B[124]), .Y(n37631) );
  NAND3X1 U32575 ( .A(n37926), .B(n37927), .C(n37928), .Y(n37904) );
  OAI21X1 U32576 ( .A(n37929), .B(n37930), .C(n25730), .Y(n37928) );
  NAND3X1 U32577 ( .A(n37931), .B(n37932), .C(n37933), .Y(n37930) );
  NOR2X1 U32578 ( .A(n37934), .B(n37935), .Y(n37933) );
  OAI22X1 U32579 ( .A(n25736), .B(n25476), .C(n25737), .D(n25317), .Y(n37935)
         );
  OAI22X1 U32580 ( .A(n25738), .B(n25323), .C(n25739), .D(n25497), .Y(n37934)
         );
  AOI22X1 U32581 ( .A(reg_A[120]), .B(n25615), .C(reg_A[123]), .D(n25616), .Y(
        n37932) );
  AOI22X1 U32582 ( .A(reg_A[122]), .B(n25607), .C(reg_A[126]), .D(n25608), .Y(
        n37931) );
  NAND3X1 U32583 ( .A(n37936), .B(n37937), .C(n37938), .Y(n37929) );
  NOR2X1 U32584 ( .A(n37939), .B(n37940), .Y(n37938) );
  OAI22X1 U32585 ( .A(n25061), .B(n25333), .C(n25746), .D(n25771), .Y(n37940)
         );
  INVX1 U32586 ( .A(reg_A[118]), .Y(n25333) );
  OAI22X1 U32587 ( .A(n25747), .B(n25335), .C(n25748), .D(n25483), .Y(n37939)
         );
  AOI22X1 U32588 ( .A(reg_A[119]), .B(n25613), .C(reg_A[116]), .D(n25749), .Y(
        n37937) );
  AOI22X1 U32589 ( .A(reg_A[117]), .B(n25750), .C(reg_A[121]), .D(n25614), .Y(
        n37936) );
  OAI21X1 U32590 ( .A(n37941), .B(n37942), .C(n25840), .Y(n37926) );
  NAND3X1 U32591 ( .A(n37943), .B(n37944), .C(n37945), .Y(n37942) );
  NOR2X1 U32592 ( .A(n37946), .B(n37947), .Y(n37945) );
  OAI22X1 U32593 ( .A(n25043), .B(n25476), .C(n25229), .D(n25396), .Y(n37947)
         );
  OAI22X1 U32594 ( .A(n25064), .B(n25436), .C(n25482), .D(n25287), .Y(n37946)
         );
  AOI22X1 U32595 ( .A(reg_A[104]), .B(n25124), .C(reg_A[101]), .D(n25222), .Y(
        n37944) );
  AOI22X1 U32596 ( .A(reg_A[102]), .B(n25637), .C(reg_A[98]), .D(n25234), .Y(
        n37943) );
  NAND3X1 U32597 ( .A(n37948), .B(n37949), .C(n37950), .Y(n37941) );
  NOR2X1 U32598 ( .A(n37951), .B(n37952), .Y(n37950) );
  OAI22X1 U32599 ( .A(n25033), .B(n25468), .C(n25040), .D(n25450), .Y(n37952)
         );
  OAI21X1 U32600 ( .A(n25041), .B(n25474), .C(n37953), .Y(n37951) );
  AOI22X1 U32601 ( .A(reg_A[96]), .B(n25247), .C(reg_A[111]), .D(n25135), .Y(
        n37953) );
  AOI22X1 U32602 ( .A(reg_A[105]), .B(n25628), .C(reg_A[108]), .D(n25067), .Y(
        n37949) );
  AOI22X1 U32603 ( .A(reg_A[107]), .B(n25123), .C(reg_A[103]), .D(n25629), .Y(
        n37948) );
  AOI21X1 U32604 ( .A(n27860), .B(reg_A[105]), .C(n37954), .Y(n37902) );
  OAI21X1 U32605 ( .A(n27839), .B(n37844), .C(n37955), .Y(n37954) );
  OAI21X1 U32606 ( .A(n37956), .B(n37957), .C(n37958), .Y(n37955) );
  OAI21X1 U32607 ( .A(n25287), .B(n25546), .C(n37959), .Y(n37957) );
  NAND3X1 U32608 ( .A(n25551), .B(n36177), .C(n37772), .Y(n37959) );
  MUX2X1 U32609 ( .B(n25474), .A(n25670), .S(reg_B[124]), .Y(n37772) );
  NOR2X1 U32610 ( .A(n25296), .B(n25544), .Y(n37956) );
  OAI21X1 U32611 ( .A(reg_B[3]), .B(n37578), .C(n37960), .Y(n37844) );
  AOI22X1 U32612 ( .A(n26530), .B(n37961), .C(n25026), .D(n36407), .Y(n37960)
         );
  MUX2X1 U32613 ( .B(reg_A[102]), .A(reg_A[110]), .S(n26596), .Y(n36407) );
  NOR2X1 U32614 ( .A(n26030), .B(reg_B[2]), .Y(n26210) );
  INVX1 U32615 ( .A(n37962), .Y(n37961) );
  INVX1 U32616 ( .A(n37963), .Y(n37578) );
  OAI21X1 U32617 ( .A(n37750), .B(n26452), .C(n37964), .Y(n37963) );
  AOI22X1 U32618 ( .A(n27859), .B(n25298), .C(n27443), .D(n25476), .Y(n37964)
         );
  NOR2X1 U32619 ( .A(n26596), .B(reg_B[2]), .Y(n27859) );
  NAND2X1 U32620 ( .A(n26028), .B(n27677), .Y(n27839) );
  INVX1 U32621 ( .A(n26525), .Y(n26028) );
  NAND2X1 U32622 ( .A(n27676), .B(n26863), .Y(n26525) );
  INVX1 U32623 ( .A(n35674), .Y(n27860) );
  NAND3X1 U32624 ( .A(n27676), .B(n26002), .C(n26664), .Y(n35674) );
  AOI22X1 U32625 ( .A(n27861), .B(reg_A[97]), .C(n27921), .D(n37965), .Y(
        n37901) );
  OAI21X1 U32626 ( .A(n27925), .B(n37573), .C(n37966), .Y(n37965) );
  AOI22X1 U32627 ( .A(n37967), .B(n26008), .C(n37823), .D(n25751), .Y(n37966)
         );
  INVX1 U32628 ( .A(n36262), .Y(n37573) );
  MUX2X1 U32629 ( .B(n25452), .A(n25448), .S(reg_B[1]), .Y(n36262) );
  NOR2X1 U32630 ( .A(n25835), .B(reg_B[0]), .Y(n27921) );
  NOR2X1 U32631 ( .A(n25835), .B(n25065), .Y(n27861) );
  NAND3X1 U32632 ( .A(n37968), .B(n37969), .C(n37970), .Y(result[111]) );
  NOR2X1 U32633 ( .A(n37971), .B(n37972), .Y(n37970) );
  NAND3X1 U32634 ( .A(n37973), .B(n37974), .C(n37975), .Y(n37972) );
  INVX1 U32635 ( .A(n37976), .Y(n37975) );
  OAI21X1 U32636 ( .A(n25424), .B(n28066), .C(n37977), .Y(n37976) );
  AOI22X1 U32637 ( .A(n25406), .B(n37978), .C(n26262), .D(n37979), .Y(n37977)
         );
  INVX1 U32638 ( .A(n37980), .Y(n28066) );
  OAI21X1 U32639 ( .A(n37981), .B(n25835), .C(n26625), .Y(n37980) );
  NAND2X1 U32640 ( .A(n25840), .B(n25235), .Y(n26625) );
  NOR2X1 U32641 ( .A(reg_B[0]), .B(n37982), .Y(n37981) );
  AOI22X1 U32642 ( .A(n37983), .B(n32116), .C(n37984), .D(n37655), .Y(n37974)
         );
  INVX1 U32643 ( .A(n25945), .Y(n32116) );
  AOI22X1 U32644 ( .A(n25696), .B(n37985), .C(n37986), .D(n37987), .Y(n37973)
         );
  NAND3X1 U32645 ( .A(n37988), .B(n37989), .C(n37990), .Y(n37971) );
  AOI21X1 U32646 ( .A(n32052), .B(reg_A[110]), .C(n37991), .Y(n37990) );
  OAI21X1 U32647 ( .A(n37992), .B(n37993), .C(n37994), .Y(n37991) );
  OAI21X1 U32648 ( .A(n37995), .B(n37996), .C(n25999), .Y(n37994) );
  OAI21X1 U32649 ( .A(n26943), .B(n25452), .C(n37997), .Y(n37996) );
  AOI22X1 U32650 ( .A(reg_A[105]), .B(n26010), .C(reg_A[104]), .D(n26002), .Y(
        n37997) );
  OAI21X1 U32651 ( .A(n31144), .B(n25474), .C(n37998), .Y(n37995) );
  AOI22X1 U32652 ( .A(reg_A[110]), .B(n26007), .C(reg_A[108]), .D(n26008), .Y(
        n37998) );
  INVX1 U32653 ( .A(n28194), .Y(n32052) );
  AOI22X1 U32654 ( .A(reg_A[107]), .B(n37999), .C(n26480), .D(n38000), .Y(
        n37989) );
  OAI21X1 U32655 ( .A(n37653), .B(n25549), .C(n38001), .Y(n38000) );
  AOI22X1 U32656 ( .A(n36148), .B(n36321), .C(n25407), .D(n38002), .Y(n38001)
         );
  OAI21X1 U32657 ( .A(n38003), .B(n38004), .C(n38005), .Y(n37999) );
  AOI21X1 U32658 ( .A(n38006), .B(n38007), .C(n27132), .Y(n38005) );
  INVX1 U32659 ( .A(n27995), .Y(n27132) );
  INVX1 U32660 ( .A(n38008), .Y(n38007) );
  AOI22X1 U32661 ( .A(n28050), .B(reg_A[106]), .C(n38009), .D(n37865), .Y(
        n37988) );
  NAND2X1 U32662 ( .A(n38010), .B(n38011), .Y(n37865) );
  AOI22X1 U32663 ( .A(n36315), .B(n37410), .C(n36442), .D(n37588), .Y(n38011)
         );
  OAI22X1 U32664 ( .A(n25448), .B(n36318), .C(n25452), .D(n36668), .Y(n37410)
         );
  AOI22X1 U32665 ( .A(n36649), .B(n37803), .C(n36280), .D(n38012), .Y(n38010)
         );
  INVX1 U32666 ( .A(n27108), .Y(n28050) );
  NOR2X1 U32667 ( .A(n38013), .B(n38014), .Y(n37969) );
  NAND3X1 U32668 ( .A(n38015), .B(n38016), .C(n38017), .Y(n38014) );
  OAI21X1 U32669 ( .A(n38018), .B(n38019), .C(n25918), .Y(n38017) );
  NAND3X1 U32670 ( .A(n38020), .B(n38021), .C(n38022), .Y(n38019) );
  NOR2X1 U32671 ( .A(n38023), .B(n38024), .Y(n38022) );
  OAI22X1 U32672 ( .A(n25736), .B(n25452), .C(n25737), .D(n25289), .Y(n38024)
         );
  OAI22X1 U32673 ( .A(n25738), .B(n25396), .C(n25739), .D(n25424), .Y(n38023)
         );
  AOI22X1 U32674 ( .A(reg_A[103]), .B(n25615), .C(reg_A[100]), .D(n25616), .Y(
        n38021) );
  AOI22X1 U32675 ( .A(reg_A[101]), .B(n25607), .C(reg_A[97]), .D(n25608), .Y(
        n38020) );
  NAND3X1 U32676 ( .A(n38025), .B(n38026), .C(n38027), .Y(n38018) );
  NOR2X1 U32677 ( .A(n38028), .B(n38029), .Y(n38027) );
  OAI22X1 U32678 ( .A(n25061), .B(n25296), .C(n25746), .D(n25474), .Y(n38029)
         );
  OAI22X1 U32679 ( .A(n25747), .B(n25469), .C(n25748), .D(n25450), .Y(n38028)
         );
  AOI22X1 U32680 ( .A(reg_A[104]), .B(n25613), .C(reg_A[107]), .D(n25749), .Y(
        n38026) );
  AOI22X1 U32681 ( .A(reg_A[106]), .B(n25750), .C(reg_A[102]), .D(n25614), .Y(
        n38025) );
  NAND2X1 U32682 ( .A(n38030), .B(n38031), .Y(n38016) );
  OAI22X1 U32683 ( .A(n25448), .B(n38032), .C(n25396), .D(n25827), .Y(n38030)
         );
  OAI21X1 U32684 ( .A(n38033), .B(n38034), .C(n25119), .Y(n38015) );
  NAND3X1 U32685 ( .A(n38035), .B(n38036), .C(n38037), .Y(n38034) );
  AOI21X1 U32686 ( .A(reg_A[111]), .B(n25125), .C(n38038), .Y(n38037) );
  OAI22X1 U32687 ( .A(n25039), .B(n25289), .C(n25231), .D(n25396), .Y(n38038)
         );
  AOI22X1 U32688 ( .A(reg_A[103]), .B(n25124), .C(reg_A[100]), .D(n25222), .Y(
        n38036) );
  AOI22X1 U32689 ( .A(reg_A[101]), .B(n25637), .C(reg_A[97]), .D(n25234), .Y(
        n38035) );
  NAND3X1 U32690 ( .A(n38039), .B(n38040), .C(n38041), .Y(n38033) );
  NOR2X1 U32691 ( .A(n38042), .B(n38043), .Y(n38041) );
  OAI22X1 U32692 ( .A(n25033), .B(n25296), .C(n25133), .D(n25474), .Y(n38043)
         );
  OAI22X1 U32693 ( .A(n25041), .B(n25469), .C(n25784), .D(n25450), .Y(n38042)
         );
  AOI22X1 U32694 ( .A(reg_A[104]), .B(n25628), .C(reg_A[107]), .D(n25067), .Y(
        n38040) );
  AOI22X1 U32695 ( .A(reg_A[106]), .B(n25123), .C(reg_A[102]), .D(n25629), .Y(
        n38039) );
  OR2X1 U32696 ( .A(n38044), .B(n38045), .Y(n38013) );
  OAI21X1 U32697 ( .A(n25668), .B(n38046), .C(n38047), .Y(n38045) );
  OAI21X1 U32698 ( .A(n38048), .B(n38049), .C(n37958), .Y(n38047) );
  INVX1 U32699 ( .A(n38050), .Y(n38048) );
  OR2X1 U32700 ( .A(n26151), .B(n38051), .Y(n38046) );
  OAI21X1 U32701 ( .A(n25672), .B(n38052), .C(n37927), .Y(n38044) );
  NAND2X1 U32702 ( .A(n26504), .B(n38053), .Y(n38052) );
  NOR2X1 U32703 ( .A(n38054), .B(n38055), .Y(n37968) );
  OAI21X1 U32704 ( .A(n29958), .B(n38056), .C(n38057), .Y(n38055) );
  AOI22X1 U32705 ( .A(n37920), .B(n37868), .C(n36778), .D(n38058), .Y(n38057)
         );
  NAND2X1 U32706 ( .A(n37014), .B(n26032), .Y(n29958) );
  NAND3X1 U32707 ( .A(n38059), .B(n38060), .C(n38061), .Y(n38054) );
  AOI22X1 U32708 ( .A(reg_B[110]), .B(n38062), .C(n38063), .D(n28138), .Y(
        n38061) );
  INVX1 U32709 ( .A(n25941), .Y(n28138) );
  NAND2X1 U32710 ( .A(n25025), .B(n30910), .Y(n25941) );
  OAI21X1 U32711 ( .A(n25031), .B(n38064), .C(n38065), .Y(n38062) );
  INVX1 U32712 ( .A(n38066), .Y(n38064) );
  OAI21X1 U32713 ( .A(n38067), .B(n38068), .C(n25310), .Y(n38060) );
  NAND3X1 U32714 ( .A(n38069), .B(n38070), .C(n38071), .Y(n38068) );
  NOR2X1 U32715 ( .A(n38072), .B(n38073), .Y(n38071) );
  OAI22X1 U32716 ( .A(n25043), .B(n25452), .C(n25039), .D(n25323), .Y(n38073)
         );
  OAI22X1 U32717 ( .A(n25064), .B(n25321), .C(n25482), .D(n25319), .Y(n38072)
         );
  AOI22X1 U32718 ( .A(reg_A[119]), .B(n25124), .C(reg_A[122]), .D(n25222), .Y(
        n38070) );
  AOI22X1 U32719 ( .A(reg_A[121]), .B(n25637), .C(reg_A[125]), .D(n25234), .Y(
        n38069) );
  NAND3X1 U32720 ( .A(n38074), .B(n38075), .C(n38076), .Y(n38067) );
  NOR2X1 U32721 ( .A(n38077), .B(n38078), .Y(n38076) );
  OAI22X1 U32722 ( .A(n25033), .B(n25332), .C(n25040), .D(n25483), .Y(n38078)
         );
  OAI21X1 U32723 ( .A(n25041), .B(n25771), .C(n38079), .Y(n38077) );
  AOI22X1 U32724 ( .A(reg_A[127]), .B(n25247), .C(reg_A[112]), .D(n25135), .Y(
        n38079) );
  AOI22X1 U32725 ( .A(reg_A[118]), .B(n25628), .C(reg_A[115]), .D(n25067), .Y(
        n38075) );
  AOI22X1 U32726 ( .A(reg_A[116]), .B(n25123), .C(reg_A[120]), .D(n25629), .Y(
        n38074) );
  OAI21X1 U32727 ( .A(n28082), .B(n38080), .C(reg_A[111]), .Y(n38059) );
  OAI21X1 U32728 ( .A(n25820), .B(n38004), .C(n38081), .Y(n38080) );
  NAND2X1 U32729 ( .A(n25561), .B(n38082), .Y(n38081) );
  OAI21X1 U32730 ( .A(reg_B[109]), .B(n38008), .C(n38083), .Y(n38082) );
  AOI21X1 U32731 ( .A(n38084), .B(n25170), .C(n26504), .Y(n38008) );
  NAND3X1 U32732 ( .A(n38085), .B(n38086), .C(n38087), .Y(result[110]) );
  NOR2X1 U32733 ( .A(n38088), .B(n38089), .Y(n38087) );
  NAND3X1 U32734 ( .A(n38090), .B(n38091), .C(n38092), .Y(n38089) );
  NOR2X1 U32735 ( .A(n38093), .B(n38094), .Y(n38092) );
  OAI21X1 U32736 ( .A(n38095), .B(n38083), .C(n38096), .Y(n38094) );
  MUX2X1 U32737 ( .B(n37992), .A(n38097), .S(reg_B[111]), .Y(n38093) );
  NAND2X1 U32738 ( .A(n38098), .B(n29315), .Y(n38097) );
  INVX1 U32739 ( .A(n38099), .Y(n37992) );
  OAI22X1 U32740 ( .A(n38100), .B(n26151), .C(n26147), .D(n38101), .Y(n38099)
         );
  MUX2X1 U32741 ( .B(n38102), .A(n38103), .S(reg_B[110]), .Y(n38101) );
  NAND2X1 U32742 ( .A(n38104), .B(n38105), .Y(n38102) );
  INVX1 U32743 ( .A(n38106), .Y(n38105) );
  AOI22X1 U32744 ( .A(n38107), .B(reg_A[106]), .C(reg_A[110]), .D(n25522), .Y(
        n38104) );
  AOI22X1 U32745 ( .A(n37978), .B(n38108), .C(n25277), .D(n38058), .Y(n38091)
         );
  OAI21X1 U32746 ( .A(n38109), .B(n36439), .C(n38110), .Y(n38058) );
  AOI22X1 U32747 ( .A(n36442), .B(n37714), .C(n37868), .D(n25428), .Y(n38110)
         );
  INVX1 U32748 ( .A(n36360), .Y(n36442) );
  NAND2X1 U32749 ( .A(reg_B[126]), .B(n36177), .Y(n36360) );
  INVX1 U32750 ( .A(n36987), .Y(n37978) );
  AOI22X1 U32751 ( .A(n26045), .B(n38111), .C(n25275), .D(n38112), .Y(n38090)
         );
  INVX1 U32752 ( .A(n37301), .Y(n25275) );
  NAND3X1 U32753 ( .A(n38113), .B(n38114), .C(n38115), .Y(n38111) );
  NOR2X1 U32754 ( .A(n38116), .B(n38117), .Y(n38115) );
  OAI21X1 U32755 ( .A(n25474), .B(n28303), .C(n38118), .Y(n38117) );
  OAI21X1 U32756 ( .A(n38119), .B(n38120), .C(n25604), .Y(n38118) );
  NAND2X1 U32757 ( .A(n38121), .B(n38122), .Y(n38120) );
  AOI22X1 U32758 ( .A(reg_A[100]), .B(n25607), .C(reg_A[96]), .D(n25608), .Y(
        n38122) );
  AOI22X1 U32759 ( .A(reg_A[98]), .B(n25609), .C(reg_A[97]), .D(n25610), .Y(
        n38121) );
  NAND2X1 U32760 ( .A(n38123), .B(n38124), .Y(n38119) );
  AOI22X1 U32761 ( .A(reg_A[103]), .B(n25613), .C(reg_A[101]), .D(n25614), .Y(
        n38124) );
  AOI22X1 U32762 ( .A(reg_A[102]), .B(n25615), .C(reg_A[99]), .D(n25616), .Y(
        n38123) );
  OAI22X1 U32763 ( .A(n25298), .B(n28311), .C(n25296), .D(n25449), .Y(n38116)
         );
  AOI22X1 U32764 ( .A(n25442), .B(reg_A[107]), .C(n27387), .D(reg_A[106]), .Y(
        n38114) );
  INVX1 U32765 ( .A(n25438), .Y(n27387) );
  INVX1 U32766 ( .A(n30437), .Y(n25442) );
  AOI22X1 U32767 ( .A(n28312), .B(reg_A[108]), .C(reg_A[110]), .D(n25434), .Y(
        n38113) );
  INVX1 U32768 ( .A(n25437), .Y(n28312) );
  NAND3X1 U32769 ( .A(n38125), .B(n38126), .C(n38127), .Y(n38088) );
  NOR2X1 U32770 ( .A(n38128), .B(n38129), .Y(n38127) );
  OAI22X1 U32771 ( .A(n32135), .B(n25450), .C(n26041), .D(n25296), .Y(n38129)
         );
  INVX1 U32772 ( .A(n28282), .Y(n26041) );
  OAI21X1 U32773 ( .A(n27523), .B(n30355), .C(n32117), .Y(n28282) );
  OAI22X1 U32774 ( .A(n32203), .B(n25298), .C(n38130), .D(n38131), .Y(n38128)
         );
  INVX1 U32775 ( .A(n26043), .Y(n32203) );
  OAI21X1 U32776 ( .A(n27523), .B(n30179), .C(n28434), .Y(n26043) );
  OAI21X1 U32777 ( .A(n38132), .B(n38133), .C(n25119), .Y(n38126) );
  NAND3X1 U32778 ( .A(n38134), .B(n38135), .C(n38136), .Y(n38133) );
  AOI21X1 U32779 ( .A(reg_A[110]), .B(n25125), .C(n38137), .Y(n38136) );
  OAI22X1 U32780 ( .A(n25039), .B(n25287), .C(n25231), .D(n25289), .Y(n38137)
         );
  AOI22X1 U32781 ( .A(reg_A[101]), .B(n25629), .C(reg_A[102]), .D(n25124), .Y(
        n38135) );
  AOI22X1 U32782 ( .A(reg_A[99]), .B(n25222), .C(reg_A[100]), .D(n25637), .Y(
        n38134) );
  NAND3X1 U32783 ( .A(n38138), .B(n38139), .C(n38140), .Y(n38132) );
  AOI21X1 U32784 ( .A(reg_A[105]), .B(n25123), .C(n38141), .Y(n38140) );
  OAI22X1 U32785 ( .A(n26431), .B(n25468), .C(n25129), .D(n25448), .Y(n38141)
         );
  AOI22X1 U32786 ( .A(reg_A[109]), .B(n25135), .C(reg_A[107]), .D(n25136), .Y(
        n38139) );
  AOI22X1 U32787 ( .A(reg_A[108]), .B(n25252), .C(reg_A[104]), .D(n25253), .Y(
        n38138) );
  AOI22X1 U32788 ( .A(reg_A[107]), .B(n28206), .C(reg_A[109]), .D(n28332), .Y(
        n38125) );
  NOR2X1 U32789 ( .A(n38142), .B(n38143), .Y(n38086) );
  OAI21X1 U32790 ( .A(n38144), .B(n38145), .C(n38146), .Y(n38143) );
  AOI22X1 U32791 ( .A(n38147), .B(n28253), .C(n38148), .D(n36280), .Y(n38146)
         );
  INVX1 U32792 ( .A(n26145), .Y(n28253) );
  NAND2X1 U32793 ( .A(reg_B[2]), .B(n30910), .Y(n26145) );
  OR2X1 U32794 ( .A(n38149), .B(n38150), .Y(n38142) );
  OAI21X1 U32795 ( .A(n38151), .B(n38152), .C(n38153), .Y(n38150) );
  OAI21X1 U32796 ( .A(n38154), .B(n36555), .C(reg_A[108]), .Y(n38153) );
  INVX1 U32797 ( .A(n37985), .Y(n38151) );
  OAI21X1 U32798 ( .A(reg_B[108]), .B(n38100), .C(n38155), .Y(n37985) );
  MUX2X1 U32799 ( .B(n38106), .A(n38156), .S(reg_B[110]), .Y(n38155) );
  NOR2X1 U32800 ( .A(n25436), .B(n38032), .Y(n38156) );
  OAI22X1 U32801 ( .A(n25361), .B(n38032), .C(n25289), .D(n25827), .Y(n38106)
         );
  MUX2X1 U32802 ( .B(n38053), .A(n38157), .S(reg_B[110]), .Y(n38100) );
  INVX1 U32803 ( .A(n38158), .Y(n38157) );
  MUX2X1 U32804 ( .B(n25468), .A(n25450), .S(n38159), .Y(n38053) );
  OAI21X1 U32805 ( .A(n38160), .B(n25468), .C(n38161), .Y(n38149) );
  OAI21X1 U32806 ( .A(n38162), .B(n38163), .C(n25310), .Y(n38161) );
  NAND3X1 U32807 ( .A(n38164), .B(n38165), .C(n38166), .Y(n38163) );
  NOR2X1 U32808 ( .A(n38167), .B(n38168), .Y(n38166) );
  OAI22X1 U32809 ( .A(n25035), .B(n25323), .C(n25036), .D(n25493), .Y(n38168)
         );
  OAI21X1 U32810 ( .A(n25027), .B(n25490), .C(n38169), .Y(n38167) );
  AOI22X1 U32811 ( .A(reg_A[119]), .B(n25629), .C(reg_A[118]), .D(n25124), .Y(
        n38169) );
  AOI22X1 U32812 ( .A(reg_A[125]), .B(n25235), .C(reg_A[122]), .D(n25635), .Y(
        n38165) );
  AOI22X1 U32813 ( .A(reg_A[123]), .B(n25325), .C(reg_A[110]), .D(n25125), .Y(
        n38164) );
  NAND3X1 U32814 ( .A(n38170), .B(n38171), .C(n38172), .Y(n38162) );
  NOR2X1 U32815 ( .A(n38173), .B(n38174), .Y(n38172) );
  OAI22X1 U32816 ( .A(n25040), .B(n25476), .C(n25254), .D(n25483), .Y(n38174)
         );
  OAI21X1 U32817 ( .A(n25042), .B(n25452), .C(n38175), .Y(n38173) );
  AOI22X1 U32818 ( .A(reg_A[127]), .B(n25246), .C(reg_A[126]), .D(n25247), .Y(
        n38175) );
  AOI22X1 U32819 ( .A(reg_A[116]), .B(n25253), .C(reg_A[117]), .D(n25628), .Y(
        n38171) );
  AOI22X1 U32820 ( .A(reg_A[114]), .B(n25074), .C(reg_A[115]), .D(n25123), .Y(
        n38170) );
  AOI21X1 U32821 ( .A(n38006), .B(n26504), .C(n26026), .Y(n38160) );
  NAND2X1 U32822 ( .A(n28122), .B(n30932), .Y(n26026) );
  NOR2X1 U32823 ( .A(n38176), .B(n38177), .Y(n38085) );
  OAI21X1 U32824 ( .A(n38178), .B(n38179), .C(n38180), .Y(n38177) );
  AOI22X1 U32825 ( .A(reg_A[111]), .B(n28280), .C(reg_A[96]), .D(n28281), .Y(
        n38180) );
  OAI22X1 U32826 ( .A(n25035), .B(n30951), .C(n25835), .D(n38181), .Y(n28281)
         );
  OAI21X1 U32827 ( .A(reg_B[0]), .B(n26530), .C(n25063), .Y(n38181) );
  INVX1 U32828 ( .A(n37987), .Y(n38178) );
  NAND2X1 U32829 ( .A(n38182), .B(n38183), .Y(n38176) );
  AOI22X1 U32830 ( .A(n26480), .B(n38184), .C(n25932), .D(n38185), .Y(n38183)
         );
  OAI21X1 U32831 ( .A(n38186), .B(n36136), .C(n38187), .Y(n38185) );
  AOI22X1 U32832 ( .A(n37868), .B(n25793), .C(reg_B[127]), .D(n38112), .Y(
        n38187) );
  MUX2X1 U32833 ( .B(n38188), .A(n38189), .S(reg_B[125]), .Y(n37868) );
  INVX1 U32834 ( .A(n37484), .Y(n38188) );
  OAI22X1 U32835 ( .A(n36318), .B(n25361), .C(n25450), .D(n36668), .Y(n37484)
         );
  INVX1 U32836 ( .A(n38049), .Y(n38186) );
  OAI21X1 U32837 ( .A(n38190), .B(n25549), .C(n38191), .Y(n38184) );
  AOI22X1 U32838 ( .A(n36321), .B(n36362), .C(n25407), .D(n36790), .Y(n38191)
         );
  AOI22X1 U32839 ( .A(n38192), .B(n26139), .C(n37984), .D(n37681), .Y(n38182)
         );
  INVX1 U32840 ( .A(n26421), .Y(n26139) );
  INVX1 U32841 ( .A(n38193), .Y(n38192) );
  NAND2X1 U32842 ( .A(n38194), .B(n38195), .Y(result[10]) );
  NOR2X1 U32843 ( .A(n38196), .B(n38197), .Y(n38195) );
  NAND3X1 U32844 ( .A(n38198), .B(n38199), .C(n38200), .Y(n38197) );
  NOR2X1 U32845 ( .A(n38201), .B(n38202), .Y(n38200) );
  OAI21X1 U32846 ( .A(n38203), .B(n25794), .C(n38204), .Y(n38202) );
  OAI21X1 U32847 ( .A(n38205), .B(n38206), .C(n26480), .Y(n38204) );
  OAI22X1 U32848 ( .A(n29239), .B(n25099), .C(n34906), .D(n25106), .Y(n38206)
         );
  INVX1 U32849 ( .A(n35466), .Y(n34906) );
  NAND2X1 U32850 ( .A(n38207), .B(n38208), .Y(n35466) );
  AOI22X1 U32851 ( .A(reg_A[22]), .B(n25156), .C(n25142), .D(reg_A[23]), .Y(
        n38208) );
  AOI22X1 U32852 ( .A(reg_A[24]), .B(n25258), .C(reg_A[25]), .D(n26761), .Y(
        n38207) );
  INVX1 U32853 ( .A(n35467), .Y(n29239) );
  NAND2X1 U32854 ( .A(n38209), .B(n38210), .Y(n35467) );
  AOI22X1 U32855 ( .A(reg_A[18]), .B(n25156), .C(n25142), .D(reg_A[19]), .Y(
        n38210) );
  AOI22X1 U32856 ( .A(reg_A[20]), .B(n25258), .C(reg_A[21]), .D(n26761), .Y(
        n38209) );
  OAI21X1 U32857 ( .A(n29240), .B(n28033), .C(n38211), .Y(n38205) );
  AOI22X1 U32858 ( .A(n25108), .B(n34908), .C(n25103), .D(n34909), .Y(n38211)
         );
  NAND2X1 U32859 ( .A(n38212), .B(n38213), .Y(n34909) );
  AOI22X1 U32860 ( .A(reg_A[26]), .B(n25156), .C(n25142), .D(reg_A[27]), .Y(
        n38213) );
  AOI22X1 U32861 ( .A(reg_A[28]), .B(n25258), .C(reg_A[29]), .D(n26761), .Y(
        n38212) );
  INVX1 U32862 ( .A(n35907), .Y(n25103) );
  NAND2X1 U32863 ( .A(n34189), .B(reg_B[27]), .Y(n35907) );
  OAI22X1 U32864 ( .A(n27954), .B(n26758), .C(n25262), .D(n29286), .Y(n34908)
         );
  INVX1 U32865 ( .A(reg_A[30]), .Y(n29286) );
  NOR2X1 U32866 ( .A(n34009), .B(n31782), .Y(n25108) );
  INVX1 U32867 ( .A(n34147), .Y(n29240) );
  NAND2X1 U32868 ( .A(n38214), .B(n38215), .Y(n34147) );
  AOI22X1 U32869 ( .A(reg_A[14]), .B(n25156), .C(n25142), .D(reg_A[15]), .Y(
        n38215) );
  AOI22X1 U32870 ( .A(reg_A[16]), .B(n25258), .C(reg_A[17]), .D(n26761), .Y(
        n38214) );
  AOI21X1 U32871 ( .A(n38216), .B(n26723), .C(n38217), .Y(n38203) );
  OAI21X1 U32872 ( .A(n30552), .B(n35887), .C(n36050), .Y(n38217) );
  NAND2X1 U32873 ( .A(n25193), .B(reg_B[13]), .Y(n36050) );
  NAND2X1 U32874 ( .A(n38218), .B(n38219), .Y(n35887) );
  AOI22X1 U32875 ( .A(n26733), .B(n30569), .C(n25172), .D(n29265), .Y(n38219)
         );
  AOI22X1 U32876 ( .A(n26734), .B(n25130), .C(n25116), .D(n26677), .Y(n38218)
         );
  INVX1 U32877 ( .A(n26691), .Y(n30552) );
  INVX1 U32878 ( .A(n35903), .Y(n38216) );
  NAND2X1 U32879 ( .A(n38220), .B(n38221), .Y(n35903) );
  MUX2X1 U32880 ( .B(n38222), .A(n38223), .S(reg_B[12]), .Y(n38221) );
  NOR2X1 U32881 ( .A(reg_A[0]), .B(n29256), .Y(n38223) );
  OAI22X1 U32882 ( .A(reg_A[7]), .B(n25194), .C(reg_A[8]), .D(n25189), .Y(
        n38222) );
  AOI22X1 U32883 ( .A(n25172), .B(n37086), .C(n25116), .D(n37080), .Y(n38220)
         );
  MUX2X1 U32884 ( .B(reg_A[10]), .A(reg_A[2]), .S(reg_B[12]), .Y(n37080) );
  MUX2X1 U32885 ( .B(reg_A[9]), .A(reg_A[1]), .S(reg_B[12]), .Y(n37086) );
  OAI21X1 U32886 ( .A(n32934), .B(n25157), .C(n38224), .Y(n38201) );
  AOI22X1 U32887 ( .A(n25168), .B(n37030), .C(n25159), .D(n25169), .Y(n38224)
         );
  OAI21X1 U32888 ( .A(n29304), .B(n25132), .C(n25190), .Y(n25169) );
  NAND2X1 U32889 ( .A(reg_A[3]), .B(n26691), .Y(n25190) );
  NOR2X1 U32890 ( .A(n25194), .B(n26147), .Y(n25159) );
  OAI21X1 U32891 ( .A(n26701), .B(n29304), .C(n38225), .Y(n37030) );
  AOI22X1 U32892 ( .A(n25193), .B(n26723), .C(reg_A[4]), .D(n26691), .Y(n38225) );
  INVX1 U32893 ( .A(n30548), .Y(n25193) );
  NAND2X1 U32894 ( .A(reg_B[12]), .B(reg_A[0]), .Y(n30548) );
  NOR2X1 U32895 ( .A(n25189), .B(n26147), .Y(n25168) );
  NAND2X1 U32896 ( .A(n35754), .B(n25932), .Y(n25157) );
  INVX1 U32897 ( .A(n36023), .Y(n35754) );
  NAND2X1 U32898 ( .A(reg_A[0]), .B(n33807), .Y(n36023) );
  AOI22X1 U32899 ( .A(n25172), .B(n25115), .C(n25116), .D(n35957), .Y(n38199)
         );
  INVX1 U32900 ( .A(n38226), .Y(n35957) );
  AOI22X1 U32901 ( .A(n36045), .B(n26267), .C(reg_A[10]), .D(n38227), .Y(
        n38226) );
  OAI21X1 U32902 ( .A(n29304), .B(n25147), .C(n38228), .Y(n36045) );
  AOI22X1 U32903 ( .A(n35865), .B(reg_A[2]), .C(reg_A[6]), .D(n26691), .Y(
        n38228) );
  OAI21X1 U32904 ( .A(n37028), .B(n26147), .C(n38229), .Y(n25115) );
  OAI21X1 U32905 ( .A(n38230), .B(n38227), .C(reg_A[9]), .Y(n38229) );
  INVX1 U32906 ( .A(n35992), .Y(n38227) );
  NAND2X1 U32907 ( .A(n26504), .B(n26723), .Y(n35992) );
  NOR2X1 U32908 ( .A(reg_B[13]), .B(n26151), .Y(n38230) );
  INVX1 U32909 ( .A(n36044), .Y(n37028) );
  OAI21X1 U32910 ( .A(n29304), .B(n25146), .C(n38231), .Y(n36044) );
  AOI22X1 U32911 ( .A(n35865), .B(reg_A[1]), .C(reg_A[5]), .D(n26691), .Y(
        n38231) );
  INVX1 U32912 ( .A(n31796), .Y(n29304) );
  AOI22X1 U32913 ( .A(n28572), .B(reg_A[1]), .C(n29324), .D(n28575), .Y(n38198) );
  INVX1 U32914 ( .A(n35839), .Y(n29324) );
  NAND2X1 U32915 ( .A(n38232), .B(n38233), .Y(n35839) );
  AOI22X1 U32916 ( .A(n26601), .B(n30569), .C(n26602), .D(n25130), .Y(n38233)
         );
  AOI22X1 U32917 ( .A(n27012), .B(n26677), .C(n26597), .D(n29265), .Y(n38232)
         );
  INVX1 U32918 ( .A(n36789), .Y(n28572) );
  NAND3X1 U32919 ( .A(n38234), .B(n38235), .C(n38236), .Y(n38196) );
  NOR2X1 U32920 ( .A(n38237), .B(n38238), .Y(n38236) );
  OAI21X1 U32921 ( .A(n38239), .B(n26990), .C(n38240), .Y(n38238) );
  OAI21X1 U32922 ( .A(n31792), .B(n28772), .C(reg_A[8]), .Y(n38240) );
  OR2X1 U32923 ( .A(n36768), .B(n25138), .Y(n28772) );
  AND2X1 U32924 ( .A(n29316), .B(n25110), .Y(n31792) );
  NOR2X1 U32925 ( .A(n29305), .B(n25024), .Y(n29316) );
  NOR2X1 U32926 ( .A(n38241), .B(n38242), .Y(n38239) );
  NAND3X1 U32927 ( .A(n38243), .B(n38244), .C(n38245), .Y(n38242) );
  NOR2X1 U32928 ( .A(n38246), .B(n38247), .Y(n38245) );
  OAI21X1 U32929 ( .A(n30587), .B(n25219), .C(n38248), .Y(n38247) );
  AOI22X1 U32930 ( .A(n25124), .B(reg_A[18]), .C(reg_A[21]), .D(n25222), .Y(
        n38248) );
  OAI21X1 U32931 ( .A(n25037), .B(n25220), .C(n38249), .Y(n38246) );
  AOI22X1 U32932 ( .A(reg_A[14]), .B(n25074), .C(n25123), .D(reg_A[15]), .Y(
        n38249) );
  AOI21X1 U32933 ( .A(reg_A[22]), .B(n25635), .C(n38250), .Y(n38244) );
  OAI22X1 U32934 ( .A(n27960), .B(n25482), .C(n25475), .D(n27962), .Y(n38250)
         );
  AOI22X1 U32935 ( .A(n25325), .B(reg_A[23]), .C(n25125), .D(reg_A[10]), .Y(
        n38243) );
  NAND3X1 U32936 ( .A(n38251), .B(n38252), .C(n38253), .Y(n38241) );
  NOR2X1 U32937 ( .A(n38254), .B(n38255), .Y(n38253) );
  OAI21X1 U32938 ( .A(n27954), .B(n26719), .C(n38256), .Y(n38255) );
  AOI22X1 U32939 ( .A(n25241), .B(reg_A[28]), .C(reg_A[30]), .D(n25339), .Y(
        n38256) );
  INVX1 U32940 ( .A(reg_A[31]), .Y(n27954) );
  OAI21X1 U32941 ( .A(n25038), .B(n25239), .C(n38257), .Y(n38254) );
  AOI22X1 U32942 ( .A(reg_A[27]), .B(n25246), .C(n25247), .D(reg_A[26]), .Y(
        n38257) );
  INVX1 U32943 ( .A(reg_A[29]), .Y(n25239) );
  AOI21X1 U32944 ( .A(n25252), .B(reg_A[12]), .C(n38258), .Y(n38252) );
  OAI22X1 U32945 ( .A(n25041), .B(n25206), .C(n25042), .D(n27967), .Y(n38258)
         );
  INVX1 U32946 ( .A(reg_A[11]), .Y(n27967) );
  AOI22X1 U32947 ( .A(reg_A[16]), .B(n25253), .C(reg_A[17]), .D(n25628), .Y(
        n38251) );
  OAI21X1 U32948 ( .A(n36000), .B(n38259), .C(n38260), .Y(n38237) );
  AOI21X1 U32949 ( .A(n38261), .B(n25382), .C(n38262), .Y(n38260) );
  INVX1 U32950 ( .A(n35646), .Y(n38262) );
  NAND2X1 U32951 ( .A(n25932), .B(n35321), .Y(n35646) );
  INVX1 U32952 ( .A(n35439), .Y(n35321) );
  NAND2X1 U32953 ( .A(reg_B[27]), .B(reg_A[0]), .Y(n35439) );
  NOR2X1 U32954 ( .A(n38263), .B(n25093), .Y(n38261) );
  NAND2X1 U32955 ( .A(reg_B[13]), .B(n37075), .Y(n25093) );
  INVX1 U32956 ( .A(n29246), .Y(n38263) );
  OAI22X1 U32957 ( .A(n25208), .B(n26692), .C(n26731), .D(n29279), .Y(n29246)
         );
  NAND2X1 U32958 ( .A(n25170), .B(n37082), .Y(n38259) );
  OAI22X1 U32959 ( .A(n26701), .B(n35857), .C(n25147), .D(n35888), .Y(n37082)
         );
  NAND2X1 U32960 ( .A(reg_B[14]), .B(n26723), .Y(n35857) );
  NAND2X1 U32961 ( .A(n25029), .B(n29302), .Y(n36000) );
  AOI22X1 U32962 ( .A(n35900), .B(n28735), .C(n35895), .D(n29247), .Y(n38235)
         );
  NAND2X1 U32963 ( .A(n38264), .B(n38265), .Y(n29247) );
  AOI22X1 U32964 ( .A(reg_A[12]), .B(n26733), .C(reg_A[11]), .D(n25172), .Y(
        n38265) );
  AOI22X1 U32965 ( .A(reg_A[13]), .B(n26734), .C(n25116), .D(reg_A[10]), .Y(
        n38264) );
  NOR2X1 U32966 ( .A(n25087), .B(n25112), .Y(n35895) );
  NAND2X1 U32967 ( .A(n26723), .B(n37075), .Y(n25112) );
  OAI21X1 U32968 ( .A(reg_B[12]), .B(n25415), .C(n26999), .Y(n37075) );
  NOR2X1 U32969 ( .A(n38266), .B(n38267), .Y(n35900) );
  OAI22X1 U32970 ( .A(n37124), .B(n27454), .C(n35642), .D(n26599), .Y(n38267)
         );
  MUX2X1 U32971 ( .B(n25147), .A(n25128), .S(reg_B[1]), .Y(n35642) );
  MUX2X1 U32972 ( .B(n25146), .A(n25177), .S(reg_B[1]), .Y(n37124) );
  OAI21X1 U32973 ( .A(reg_A[0]), .B(n28739), .C(n38268), .Y(n38266) );
  AOI22X1 U32974 ( .A(n28741), .B(n25132), .C(n28742), .D(n26701), .Y(n38268)
         );
  AOI22X1 U32975 ( .A(n28726), .B(reg_A[15]), .C(n28802), .D(reg_A[14]), .Y(
        n38234) );
  NOR2X1 U32976 ( .A(n38269), .B(n38270), .Y(n38194) );
  NAND3X1 U32977 ( .A(n38271), .B(n38272), .C(n38273), .Y(n38270) );
  NOR2X1 U32978 ( .A(n38274), .B(n38275), .Y(n38273) );
  OAI22X1 U32979 ( .A(n38276), .B(n37095), .C(n25130), .D(n28562), .Y(n38275)
         );
  NAND2X1 U32980 ( .A(reg_A[8]), .B(n26504), .Y(n37095) );
  INVX1 U32981 ( .A(n35888), .Y(n38276) );
  NAND2X1 U32982 ( .A(n26723), .B(n29256), .Y(n35888) );
  OAI21X1 U32983 ( .A(n29241), .B(n30559), .C(n38277), .Y(n38274) );
  OAI21X1 U32984 ( .A(n38278), .B(n38279), .C(n25119), .Y(n38277) );
  OR2X1 U32985 ( .A(n38280), .B(n38281), .Y(n38279) );
  OAI22X1 U32986 ( .A(n25147), .B(n25228), .C(n25128), .D(n25467), .Y(n38281)
         );
  OAI21X1 U32987 ( .A(n25177), .B(n25223), .C(n38282), .Y(n38280) );
  AOI22X1 U32988 ( .A(n25075), .B(reg_A[6]), .C(n25123), .D(reg_A[5]), .Y(
        n38282) );
  OR2X1 U32989 ( .A(n38283), .B(n38284), .Y(n38278) );
  OAI22X1 U32990 ( .A(n25130), .B(n25129), .C(n30569), .D(n25131), .Y(n38284)
         );
  OAI21X1 U32991 ( .A(n26701), .B(n25133), .C(n38285), .Y(n38283) );
  AOI22X1 U32992 ( .A(n25135), .B(reg_A[9]), .C(n25136), .D(reg_A[7]), .Y(
        n38285) );
  NAND2X1 U32993 ( .A(n26480), .B(n25110), .Y(n30559) );
  INVX1 U32994 ( .A(n34146), .Y(n29241) );
  NAND2X1 U32995 ( .A(n38286), .B(n38287), .Y(n34146) );
  AOI22X1 U32996 ( .A(reg_A[10]), .B(n25156), .C(n25142), .D(reg_A[11]), .Y(
        n38287) );
  AOI22X1 U32997 ( .A(reg_A[12]), .B(n25258), .C(reg_A[13]), .D(n26761), .Y(
        n38286) );
  AOI22X1 U32998 ( .A(reg_A[0]), .B(n28700), .C(reg_A[10]), .D(n28661), .Y(
        n38272) );
  NAND2X1 U32999 ( .A(n38288), .B(n28512), .Y(n28700) );
  AOI22X1 U33000 ( .A(reg_A[9]), .B(n26626), .C(n38289), .D(n26756), .Y(n38271) );
  OAI21X1 U33001 ( .A(n26757), .B(n25264), .C(n38290), .Y(n38289) );
  AOI22X1 U33002 ( .A(n25156), .B(n37110), .C(n25142), .D(n36098), .Y(n38290)
         );
  OAI22X1 U33003 ( .A(n35675), .B(reg_B[29]), .C(n28033), .D(n29265), .Y(
        n36098) );
  INVX1 U33004 ( .A(n35743), .Y(n35675) );
  OAI22X1 U33005 ( .A(n33807), .B(n25146), .C(n34465), .D(n25177), .Y(n35743)
         );
  INVX1 U33006 ( .A(reg_A[9]), .Y(n25146) );
  INVX1 U33007 ( .A(n35920), .Y(n37110) );
  AOI22X1 U33008 ( .A(n35616), .B(n33955), .C(reg_A[6]), .D(n25101), .Y(n35920) );
  OAI22X1 U33009 ( .A(n33807), .B(n25147), .C(n25128), .D(n34465), .Y(n35616)
         );
  INVX1 U33010 ( .A(reg_A[10]), .Y(n25147) );
  INVX1 U33011 ( .A(n25259), .Y(n26757) );
  OAI22X1 U33012 ( .A(n25132), .B(n26775), .C(n25130), .D(n28033), .Y(n25259)
         );
  NAND3X1 U33013 ( .A(n38291), .B(n38292), .C(n38293), .Y(n38269) );
  NOR2X1 U33014 ( .A(n38294), .B(n38295), .Y(n38293) );
  OAI22X1 U33015 ( .A(n29265), .B(n28571), .C(n25128), .D(n25178), .Y(n38295)
         );
  OAI21X1 U33016 ( .A(n26677), .B(n28679), .C(n38296), .Y(n38294) );
  AOI22X1 U33017 ( .A(n25180), .B(reg_A[7]), .C(n28576), .D(reg_A[4]), .Y(
        n38296) );
  INVX1 U33018 ( .A(n28715), .Y(n25180) );
  AOI22X1 U33019 ( .A(n25152), .B(reg_A[13]), .C(n25153), .D(reg_A[12]), .Y(
        n38292) );
  AOI22X1 U33020 ( .A(n28280), .B(reg_A[11]), .C(n25258), .D(n25143), .Y(
        n38291) );
  OAI21X1 U33021 ( .A(n27438), .B(n38297), .C(n38298), .Y(n25143) );
  OAI21X1 U33022 ( .A(n38299), .B(n38300), .C(n25699), .Y(n38298) );
  INVX1 U33023 ( .A(n38297), .Y(n38300) );
  AND2X1 U33024 ( .A(n33955), .B(n35846), .Y(n38299) );
  OAI22X1 U33025 ( .A(n26701), .B(n33807), .C(n26742), .D(n34465), .Y(n35846)
         );
  NAND2X1 U33026 ( .A(n25101), .B(reg_A[4]), .Y(n38297) );
  NAND3X1 U33027 ( .A(n38301), .B(n38302), .C(n38303), .Y(result[109]) );
  NOR2X1 U33028 ( .A(n38304), .B(n38305), .Y(n38303) );
  NAND3X1 U33029 ( .A(n38306), .B(n38096), .C(n38307), .Y(n38305) );
  NOR2X1 U33030 ( .A(n38308), .B(n38309), .Y(n38307) );
  OAI21X1 U33031 ( .A(n25474), .B(n38310), .C(n38311), .Y(n38309) );
  OAI21X1 U33032 ( .A(n38312), .B(n38313), .C(n26045), .Y(n38311) );
  NAND3X1 U33033 ( .A(n38314), .B(n38315), .C(n38316), .Y(n38313) );
  AOI21X1 U33034 ( .A(reg_A[109]), .B(n25434), .C(n38317), .Y(n38316) );
  OAI22X1 U33035 ( .A(n28353), .B(n25470), .C(n25205), .D(n25296), .Y(n38317)
         );
  INVX1 U33036 ( .A(n27242), .Y(n25205) );
  AOI22X1 U33037 ( .A(n25097), .B(n38318), .C(reg_A[104]), .D(n28355), .Y(
        n38315) );
  AOI22X1 U33038 ( .A(reg_A[108]), .B(n25441), .C(reg_A[106]), .D(n27241), .Y(
        n38314) );
  NAND3X1 U33039 ( .A(n38319), .B(n38320), .C(n38321), .Y(n38312) );
  NOR2X1 U33040 ( .A(n38322), .B(n38323), .Y(n38321) );
  OAI22X1 U33041 ( .A(n28361), .B(n25424), .C(n25448), .D(n28311), .Y(n38323)
         );
  INVX1 U33042 ( .A(n27648), .Y(n28361) );
  OAI21X1 U33043 ( .A(n25403), .B(n25229), .C(n25453), .Y(n27648) );
  NAND2X1 U33044 ( .A(n25610), .B(n25604), .Y(n25453) );
  OAI22X1 U33045 ( .A(n25396), .B(n28362), .C(n25289), .D(n28363), .Y(n38322)
         );
  NAND2X1 U33046 ( .A(n25616), .B(n25604), .Y(n28363) );
  NAND2X1 U33047 ( .A(n25607), .B(n25604), .Y(n28362) );
  AOI22X1 U33048 ( .A(n28364), .B(reg_A[97]), .C(n25500), .D(reg_A[100]), .Y(
        n38320) );
  INVX1 U33049 ( .A(n26229), .Y(n25500) );
  NAND2X1 U33050 ( .A(n25614), .B(n25604), .Y(n26229) );
  INVX1 U33051 ( .A(n25451), .Y(n28364) );
  NAND2X1 U33052 ( .A(n25609), .B(n25604), .Y(n25451) );
  AOI22X1 U33053 ( .A(n25501), .B(reg_A[101]), .C(n25502), .D(reg_A[102]), .Y(
        n38319) );
  INVX1 U33054 ( .A(n30443), .Y(n25502) );
  NAND2X1 U33055 ( .A(n25613), .B(n25604), .Y(n30443) );
  INVX1 U33056 ( .A(n30444), .Y(n25501) );
  NAND2X1 U33057 ( .A(n25615), .B(n25604), .Y(n30444) );
  OAI22X1 U33058 ( .A(n38324), .B(n36987), .C(n25994), .D(n38325), .Y(n38308)
         );
  AOI21X1 U33059 ( .A(reg_B[110]), .B(n38326), .C(n38327), .Y(n38096) );
  AOI22X1 U33060 ( .A(n27676), .B(n38318), .C(n38328), .D(n25689), .Y(n38306)
         );
  NAND3X1 U33061 ( .A(n38329), .B(n38330), .C(n38331), .Y(n38318) );
  NOR2X1 U33062 ( .A(n38332), .B(n38333), .Y(n38331) );
  OAI21X1 U33063 ( .A(n25043), .B(n25474), .C(n38334), .Y(n38333) );
  AOI22X1 U33064 ( .A(reg_A[99]), .B(n25637), .C(reg_A[97]), .D(n25635), .Y(
        n38334) );
  OAI21X1 U33065 ( .A(n25027), .B(n25289), .C(n38335), .Y(n38332) );
  AOI22X1 U33066 ( .A(reg_A[100]), .B(n25629), .C(reg_A[101]), .D(n25124), .Y(
        n38335) );
  NOR2X1 U33067 ( .A(n38336), .B(n38337), .Y(n38330) );
  OAI22X1 U33068 ( .A(n25033), .B(n25448), .C(n25040), .D(n25470), .Y(n38337)
         );
  OAI22X1 U33069 ( .A(n25041), .B(n25468), .C(n25042), .D(n25469), .Y(n38336)
         );
  AOI21X1 U33070 ( .A(reg_A[104]), .B(n25123), .C(n38338), .Y(n38329) );
  OAI22X1 U33071 ( .A(n26431), .B(n25296), .C(n25030), .D(n25361), .Y(n38338)
         );
  NAND3X1 U33072 ( .A(n38339), .B(n38340), .C(n38341), .Y(n38304) );
  AOI21X1 U33073 ( .A(n38031), .B(n37987), .C(n38342), .Y(n38341) );
  OAI22X1 U33074 ( .A(n38343), .B(n38130), .C(n25148), .D(n25450), .Y(n38342)
         );
  NAND2X1 U33075 ( .A(n38344), .B(n38345), .Y(n37987) );
  AOI22X1 U33076 ( .A(n38346), .B(reg_A[97]), .C(n38347), .D(reg_A[101]), .Y(
        n38345) );
  AOI22X1 U33077 ( .A(n38107), .B(reg_A[105]), .C(reg_A[109]), .D(n25522), .Y(
        n38344) );
  AOI22X1 U33078 ( .A(n25560), .B(n38348), .C(n37979), .D(n25150), .Y(n38340)
         );
  AOI21X1 U33079 ( .A(n38349), .B(reg_B[2]), .C(n38350), .Y(n37979) );
  INVX1 U33080 ( .A(n38351), .Y(n38350) );
  AOI22X1 U33081 ( .A(n26293), .B(n36466), .C(n26295), .D(n36604), .Y(n38351)
         );
  INVX1 U33082 ( .A(n37750), .Y(n36604) );
  MUX2X1 U33083 ( .B(n25469), .A(n25436), .S(reg_B[1]), .Y(n37750) );
  INVX1 U33084 ( .A(n37967), .Y(n36466) );
  MUX2X1 U33085 ( .B(n25474), .A(n25670), .S(reg_B[1]), .Y(n37967) );
  AOI22X1 U33086 ( .A(n37984), .B(n37855), .C(reg_A[111]), .D(n25153), .Y(
        n38339) );
  NOR2X1 U33087 ( .A(n38352), .B(n38353), .Y(n38302) );
  NAND3X1 U33088 ( .A(n38354), .B(n38355), .C(n38356), .Y(n38353) );
  AOI22X1 U33089 ( .A(n37983), .B(n32319), .C(n36778), .D(n38357), .Y(n38356)
         );
  NOR2X1 U33090 ( .A(n37229), .B(n25697), .Y(n36778) );
  INVX1 U33091 ( .A(n26278), .Y(n32319) );
  NAND2X1 U33092 ( .A(n30427), .B(n26030), .Y(n26278) );
  AND2X1 U33093 ( .A(n38358), .B(n38359), .Y(n37983) );
  AOI22X1 U33094 ( .A(n26292), .B(n25296), .C(n26293), .D(n25474), .Y(n38359)
         );
  AOI22X1 U33095 ( .A(n26294), .B(n25298), .C(n26295), .D(n25469), .Y(n38358)
         );
  OAI21X1 U33096 ( .A(n38360), .B(n38361), .C(n25310), .Y(n38355) );
  NAND3X1 U33097 ( .A(n38362), .B(n38363), .C(n38364), .Y(n38361) );
  NOR2X1 U33098 ( .A(n38365), .B(n38366), .Y(n38364) );
  OAI22X1 U33099 ( .A(n25035), .B(n25321), .C(n25036), .D(n36140), .Y(n38366)
         );
  OAI21X1 U33100 ( .A(n25027), .B(n25493), .C(n38367), .Y(n38365) );
  AOI22X1 U33101 ( .A(reg_A[118]), .B(n25629), .C(reg_A[117]), .D(n25124), .Y(
        n38367) );
  AOI22X1 U33102 ( .A(reg_A[124]), .B(n25235), .C(reg_A[121]), .D(n25635), .Y(
        n38363) );
  AOI22X1 U33103 ( .A(reg_A[122]), .B(n25325), .C(reg_A[109]), .D(n25125), .Y(
        n38362) );
  NAND3X1 U33104 ( .A(n38368), .B(n38369), .C(n38370), .Y(n38360) );
  NOR2X1 U33105 ( .A(n38371), .B(n38372), .Y(n38370) );
  OAI22X1 U33106 ( .A(n25041), .B(n25476), .C(n25042), .D(n25450), .Y(n38372)
         );
  OAI21X1 U33107 ( .A(n25051), .B(n25497), .C(n38373), .Y(n38371) );
  AOI22X1 U33108 ( .A(reg_A[126]), .B(n25246), .C(reg_A[125]), .D(n25247), .Y(
        n38373) );
  AOI21X1 U33109 ( .A(reg_A[116]), .B(n25628), .C(n38374), .Y(n38369) );
  OAI22X1 U33110 ( .A(n25033), .B(n25335), .C(n25040), .D(n25452), .Y(n38374)
         );
  AOI22X1 U33111 ( .A(reg_A[113]), .B(n25074), .C(reg_A[114]), .D(n25123), .Y(
        n38368) );
  OAI21X1 U33112 ( .A(n38154), .B(n38375), .C(reg_A[107]), .Y(n38354) );
  INVX1 U33113 ( .A(n28415), .Y(n38375) );
  NAND2X1 U33114 ( .A(n30427), .B(n26009), .Y(n28415) );
  NOR2X1 U33115 ( .A(n38144), .B(n25668), .Y(n38154) );
  NAND3X1 U33116 ( .A(n38376), .B(n38065), .C(n38377), .Y(n38352) );
  AOI22X1 U33117 ( .A(n38378), .B(n25559), .C(n38379), .D(n26186), .Y(n38377)
         );
  INVX1 U33118 ( .A(n38380), .Y(n38379) );
  MUX2X1 U33119 ( .B(n38098), .A(n38381), .S(reg_B[111]), .Y(n38380) );
  OAI22X1 U33120 ( .A(reg_B[110]), .B(n38051), .C(n25470), .D(n38382), .Y(
        n38098) );
  AND2X1 U33121 ( .A(n38103), .B(n26267), .Y(n38378) );
  NAND3X1 U33122 ( .A(reg_B[109]), .B(n25696), .C(n38383), .Y(n38065) );
  NAND3X1 U33123 ( .A(n26504), .B(n25521), .C(n38066), .Y(n38376) );
  MUX2X1 U33124 ( .B(n38051), .A(n38158), .S(reg_B[111]), .Y(n38066) );
  MUX2X1 U33125 ( .B(reg_A[109]), .A(reg_A[105]), .S(reg_B[109]), .Y(n38051)
         );
  NOR2X1 U33126 ( .A(n38384), .B(n38385), .Y(n38301) );
  OAI21X1 U33127 ( .A(n38386), .B(n38387), .C(n38388), .Y(n38385) );
  AOI22X1 U33128 ( .A(n38112), .B(n38009), .C(n32356), .D(reg_A[106]), .Y(
        n38388) );
  INVX1 U33129 ( .A(n28379), .Y(n32356) );
  NAND2X1 U33130 ( .A(n30427), .B(n26008), .Y(n28379) );
  OR2X1 U33131 ( .A(n36329), .B(n36436), .Y(n38009) );
  OAI21X1 U33132 ( .A(n38389), .B(n25428), .C(n38390), .Y(n38112) );
  AOI22X1 U33133 ( .A(n36315), .B(n37588), .C(n36649), .D(n38012), .Y(n38390)
         );
  INVX1 U33134 ( .A(n36312), .Y(n36649) );
  OAI22X1 U33135 ( .A(n36318), .B(n25670), .C(n25474), .D(n36668), .Y(n37588)
         );
  INVX1 U33136 ( .A(n36359), .Y(n36315) );
  INVX1 U33137 ( .A(n38391), .Y(n38386) );
  NAND2X1 U33138 ( .A(n38392), .B(n38393), .Y(n38384) );
  AOI22X1 U33139 ( .A(n28453), .B(reg_A[96]), .C(n26480), .D(n38394), .Y(
        n38393) );
  OAI21X1 U33140 ( .A(n38395), .B(n25549), .C(n38396), .Y(n38394) );
  AOI22X1 U33141 ( .A(n36321), .B(n36911), .C(n25407), .D(n36877), .Y(n38396)
         );
  NOR2X1 U33142 ( .A(n25835), .B(n38397), .Y(n28453) );
  OAI21X1 U33143 ( .A(reg_B[0]), .B(n38398), .C(n25063), .Y(n38397) );
  AOI22X1 U33144 ( .A(n25932), .B(n38399), .C(n32292), .D(reg_A[104]), .Y(
        n38392) );
  INVX1 U33145 ( .A(n28434), .Y(n32292) );
  OAI21X1 U33146 ( .A(n25793), .B(n38050), .C(n38400), .Y(n38399) );
  AOI22X1 U33147 ( .A(n25700), .B(n38049), .C(n25355), .D(n38401), .Y(n38400)
         );
  NAND2X1 U33148 ( .A(n38402), .B(n38403), .Y(result[108]) );
  NOR2X1 U33149 ( .A(n38404), .B(n38405), .Y(n38403) );
  NAND3X1 U33150 ( .A(n38406), .B(n38407), .C(n38408), .Y(n38405) );
  NOR2X1 U33151 ( .A(n38409), .B(n38410), .Y(n38408) );
  OAI22X1 U33152 ( .A(n26421), .B(n38411), .C(n25396), .D(n36789), .Y(n38410)
         );
  NAND2X1 U33153 ( .A(n37014), .B(n26452), .Y(n26421) );
  OAI22X1 U33154 ( .A(n32432), .B(n25468), .C(n32433), .D(n25296), .Y(n38409)
         );
  INVX1 U33155 ( .A(n28495), .Y(n32433) );
  NAND2X1 U33156 ( .A(n35859), .B(n28715), .Y(n28495) );
  INVX1 U33157 ( .A(n28206), .Y(n35859) );
  OAI22X1 U33158 ( .A(n27523), .B(n36451), .C(n38412), .D(n30090), .Y(n28206)
         );
  INVX1 U33159 ( .A(n28496), .Y(n32432) );
  NAND2X1 U33160 ( .A(n28276), .B(n32817), .Y(n28496) );
  INVX1 U33161 ( .A(n36555), .Y(n28276) );
  OAI21X1 U33162 ( .A(n38412), .B(n31144), .C(n30486), .Y(n36555) );
  NAND2X1 U33163 ( .A(n27388), .B(n26045), .Y(n30486) );
  INVX1 U33164 ( .A(n38413), .Y(n27388) );
  INVX1 U33165 ( .A(n38414), .Y(n38412) );
  AOI22X1 U33166 ( .A(n28649), .B(reg_A[98]), .C(n26480), .D(n38415), .Y(
        n38407) );
  OAI21X1 U33167 ( .A(n38416), .B(n25549), .C(n38417), .Y(n38415) );
  AOI22X1 U33168 ( .A(n36321), .B(n36619), .C(n25407), .D(n37883), .Y(n38417)
         );
  INVX1 U33169 ( .A(n36141), .Y(n36321) );
  INVX1 U33170 ( .A(n28512), .Y(n28649) );
  AOI22X1 U33171 ( .A(n25562), .B(n38348), .C(reg_A[96]), .D(n28494), .Y(
        n38406) );
  NAND3X1 U33172 ( .A(n38418), .B(n26917), .C(n38419), .Y(n28494) );
  INVX1 U33173 ( .A(n36558), .Y(n38419) );
  OAI21X1 U33174 ( .A(n30990), .B(n25738), .C(n30827), .Y(n36558) );
  NAND2X1 U33175 ( .A(n25840), .B(n25635), .Y(n26917) );
  OAI21X1 U33176 ( .A(n26455), .B(reg_B[0]), .C(n27676), .Y(n38418) );
  OAI22X1 U33177 ( .A(n38420), .B(n26147), .C(n25468), .D(n38144), .Y(n38348)
         );
  NAND3X1 U33178 ( .A(n38421), .B(n38422), .C(n38423), .Y(n38404) );
  NOR2X1 U33179 ( .A(n38424), .B(n38425), .Y(n38423) );
  OAI21X1 U33180 ( .A(n38426), .B(n25469), .C(n38427), .Y(n38425) );
  OAI21X1 U33181 ( .A(n38428), .B(n38429), .C(n25310), .Y(n38427) );
  NAND3X1 U33182 ( .A(n38430), .B(n38431), .C(n38432), .Y(n38429) );
  NOR2X1 U33183 ( .A(n38433), .B(n38434), .Y(n38432) );
  OAI22X1 U33184 ( .A(n25043), .B(n25469), .C(n25039), .D(n25490), .Y(n38434)
         );
  OAI21X1 U33185 ( .A(n25064), .B(n25493), .C(n38435), .Y(n38433) );
  AOI22X1 U33186 ( .A(reg_A[122]), .B(n25234), .C(reg_A[123]), .D(n25235), .Y(
        n38435) );
  AOI21X1 U33187 ( .A(reg_A[116]), .B(n25124), .C(n38436), .Y(n38431) );
  OAI22X1 U33188 ( .A(n25037), .B(n25332), .C(n26703), .D(n25483), .Y(n38436)
         );
  AOI22X1 U33189 ( .A(reg_A[119]), .B(n25222), .C(reg_A[118]), .D(n25637), .Y(
        n38430) );
  NAND3X1 U33190 ( .A(n38437), .B(n38438), .C(n38439), .Y(n38428) );
  NOR2X1 U33191 ( .A(n38440), .B(n38441), .Y(n38439) );
  OAI22X1 U33192 ( .A(n25042), .B(n25474), .C(n25331), .D(n25319), .Y(n38441)
         );
  OAI21X1 U33193 ( .A(n25038), .B(n25497), .C(n38442), .Y(n38440) );
  AOI22X1 U33194 ( .A(reg_A[125]), .B(n25246), .C(reg_A[124]), .D(n25247), .Y(
        n38442) );
  AOI21X1 U33195 ( .A(reg_A[114]), .B(n25253), .C(n38443), .Y(n38438) );
  OAI22X1 U33196 ( .A(n25040), .B(n25450), .C(n25254), .D(n25452), .Y(n38443)
         );
  AOI22X1 U33197 ( .A(reg_A[115]), .B(n25628), .C(reg_A[112]), .D(n25066), .Y(
        n38437) );
  INVX1 U33198 ( .A(n38444), .Y(n38426) );
  OAI21X1 U33199 ( .A(n38144), .B(n25669), .C(n32495), .Y(n38444) );
  INVX1 U33200 ( .A(n28563), .Y(n32495) );
  NAND3X1 U33201 ( .A(n32827), .B(n30908), .C(n32135), .Y(n28563) );
  INVX1 U33202 ( .A(n28082), .Y(n32135) );
  NAND2X1 U33203 ( .A(n38310), .B(n36307), .Y(n28082) );
  NAND2X1 U33204 ( .A(n26004), .B(n38414), .Y(n36307) );
  NAND2X1 U33205 ( .A(n30792), .B(n26045), .Y(n30908) );
  NAND2X1 U33206 ( .A(n26504), .B(n38159), .Y(n38144) );
  OAI21X1 U33207 ( .A(n38445), .B(n27438), .C(n38446), .Y(n38424) );
  AOI22X1 U33208 ( .A(n25119), .B(n38447), .C(n38448), .D(n26756), .Y(n38446)
         );
  OAI22X1 U33209 ( .A(n38449), .B(n36246), .C(n38389), .D(n25568), .Y(n38448)
         );
  NAND2X1 U33210 ( .A(n38450), .B(n38451), .Y(n38447) );
  NOR2X1 U33211 ( .A(n38452), .B(n38453), .Y(n38451) );
  OAI21X1 U33212 ( .A(n25043), .B(n25469), .C(n38454), .Y(n38453) );
  AOI22X1 U33213 ( .A(reg_A[107]), .B(n25135), .C(reg_A[106]), .D(n25252), .Y(
        n38454) );
  OAI21X1 U33214 ( .A(n25028), .B(n25448), .C(n38455), .Y(n38452) );
  AOI22X1 U33215 ( .A(reg_A[105]), .B(n25136), .C(reg_A[104]), .D(n25066), .Y(
        n38455) );
  NOR2X1 U33216 ( .A(n38456), .B(n38457), .Y(n38450) );
  OAI21X1 U33217 ( .A(n25034), .B(n25436), .C(n38458), .Y(n38457) );
  AOI22X1 U33218 ( .A(reg_A[102]), .B(n25253), .C(reg_A[101]), .D(n25628), .Y(
        n38458) );
  OAI21X1 U33219 ( .A(n25036), .B(n25289), .C(n38459), .Y(n38456) );
  AOI22X1 U33220 ( .A(reg_A[99]), .B(n25629), .C(reg_A[97]), .D(n25222), .Y(
        n38459) );
  AOI22X1 U33221 ( .A(n25793), .B(n38049), .C(n25399), .D(n38401), .Y(n38445)
         );
  OAI22X1 U33222 ( .A(n37866), .B(reg_B[125]), .C(n25298), .D(n25544), .Y(
        n38049) );
  AOI22X1 U33223 ( .A(n38460), .B(n38391), .C(n38461), .D(n38103), .Y(n38422)
         );
  NAND2X1 U33224 ( .A(n38462), .B(n38463), .Y(n38103) );
  AOI22X1 U33225 ( .A(n38346), .B(reg_A[96]), .C(n38347), .D(reg_A[100]), .Y(
        n38463) );
  INVX1 U33226 ( .A(n25827), .Y(n38346) );
  NAND2X1 U33227 ( .A(reg_B[108]), .B(reg_B[109]), .Y(n25827) );
  AOI22X1 U33228 ( .A(n38107), .B(reg_A[104]), .C(reg_A[108]), .D(n25522), .Y(
        n38462) );
  OAI21X1 U33229 ( .A(n38032), .B(n38464), .C(n38465), .Y(n38391) );
  AOI22X1 U33230 ( .A(n38466), .B(n38107), .C(n38381), .D(n38467), .Y(n38465)
         );
  NOR2X1 U33231 ( .A(n25521), .B(n25361), .Y(n38466) );
  INVX1 U33232 ( .A(n38468), .Y(n38464) );
  INVX1 U33233 ( .A(n38152), .Y(n38460) );
  AOI22X1 U33234 ( .A(n36436), .B(n38357), .C(n28549), .D(reg_A[97]), .Y(
        n38421) );
  INVX1 U33235 ( .A(n38469), .Y(n38357) );
  AOI21X1 U33236 ( .A(n38401), .B(reg_B[126]), .C(n38470), .Y(n38469) );
  OAI22X1 U33237 ( .A(n36359), .B(n37866), .C(n36312), .D(n38109), .Y(n38470)
         );
  NAND2X1 U33238 ( .A(reg_B[125]), .B(n25428), .Y(n36312) );
  INVX1 U33239 ( .A(n37714), .Y(n37866) );
  OAI22X1 U33240 ( .A(n36318), .B(n25436), .C(n25469), .D(n36668), .Y(n37714)
         );
  NAND2X1 U33241 ( .A(n36177), .B(n25428), .Y(n36359) );
  NOR2X1 U33242 ( .A(n25375), .B(n25697), .Y(n36436) );
  INVX1 U33243 ( .A(n37226), .Y(n25375) );
  NOR2X1 U33244 ( .A(n25403), .B(reg_B[127]), .Y(n37226) );
  NOR2X1 U33245 ( .A(n38471), .B(n38472), .Y(n38402) );
  NAND3X1 U33246 ( .A(n38473), .B(n38474), .C(n38475), .Y(n38472) );
  NOR2X1 U33247 ( .A(n38476), .B(n38477), .Y(n38475) );
  OAI22X1 U33248 ( .A(n25808), .B(n36987), .C(n32494), .D(n25298), .Y(n38477)
         );
  INVX1 U33249 ( .A(n26348), .Y(n32494) );
  OAI21X1 U33250 ( .A(n26452), .B(n29998), .C(n38478), .Y(n26348) );
  NOR2X1 U33251 ( .A(n25181), .B(n26269), .Y(n38478) );
  INVX1 U33252 ( .A(n30932), .Y(n26269) );
  NAND2X1 U33253 ( .A(n30357), .B(n26045), .Y(n30932) );
  INVX1 U33254 ( .A(n31058), .Y(n30357) );
  INVX1 U33255 ( .A(n28679), .Y(n25181) );
  NAND2X1 U33256 ( .A(n26480), .B(n25427), .Y(n36987) );
  OAI22X1 U33257 ( .A(n38131), .B(n38479), .C(n32496), .D(n25470), .Y(n38476)
         );
  NOR2X1 U33258 ( .A(n28332), .B(n32880), .Y(n32496) );
  OAI21X1 U33259 ( .A(n27523), .B(n30791), .C(n28194), .Y(n28332) );
  NAND2X1 U33260 ( .A(n26007), .B(n38414), .Y(n28194) );
  OAI21X1 U33261 ( .A(reg_B[1]), .B(n26864), .C(n29998), .Y(n38414) );
  AOI22X1 U33262 ( .A(n32498), .B(reg_A[101]), .C(n38328), .D(n25825), .Y(
        n38474) );
  NOR2X1 U33263 ( .A(n38480), .B(n38481), .Y(n38473) );
  MUX2X1 U33264 ( .B(n38482), .A(n38483), .S(reg_B[111]), .Y(n38481) );
  NAND2X1 U33265 ( .A(n38484), .B(n29315), .Y(n38483) );
  NAND2X1 U33266 ( .A(n26186), .B(n38381), .Y(n38482) );
  OAI22X1 U33267 ( .A(reg_B[110]), .B(n38158), .C(n25468), .D(n38382), .Y(
        n38381) );
  MUX2X1 U33268 ( .B(reg_A[108]), .A(reg_A[104]), .S(reg_B[109]), .Y(n38158)
         );
  NAND3X1 U33269 ( .A(n38485), .B(n38486), .C(n38487), .Y(n38471) );
  NOR2X1 U33270 ( .A(n38488), .B(n38489), .Y(n38487) );
  OAI22X1 U33271 ( .A(n38490), .B(n36960), .C(n28571), .D(n25448), .Y(n38489)
         );
  OAI21X1 U33272 ( .A(n25178), .B(n25436), .C(n38491), .Y(n38488) );
  AOI22X1 U33273 ( .A(n38492), .B(n28575), .C(n28576), .D(reg_A[102]), .Y(
        n38491) );
  INVX1 U33274 ( .A(n28714), .Y(n28576) );
  AOI22X1 U33275 ( .A(reg_A[111]), .B(n25152), .C(reg_A[110]), .D(n25153), .Y(
        n38486) );
  AOI22X1 U33276 ( .A(reg_A[109]), .B(n28280), .C(n38493), .D(n38494), .Y(
        n38485) );
  NAND2X1 U33277 ( .A(n38495), .B(n38496), .Y(result[107]) );
  NOR2X1 U33278 ( .A(n38497), .B(n38498), .Y(n38496) );
  NAND3X1 U33279 ( .A(n38499), .B(n38500), .C(n38501), .Y(n38498) );
  NOR2X1 U33280 ( .A(n38502), .B(n38503), .Y(n38501) );
  OAI22X1 U33281 ( .A(n25178), .B(n25396), .C(n28679), .D(n25448), .Y(n38503)
         );
  NAND2X1 U33282 ( .A(n25749), .B(n25918), .Y(n28679) );
  NAND2X1 U33283 ( .A(n25615), .B(n25918), .Y(n25178) );
  OAI22X1 U33284 ( .A(n25670), .B(n28714), .C(n25289), .D(n36789), .Y(n38502)
         );
  NAND2X1 U33285 ( .A(n25614), .B(n25918), .Y(n36789) );
  NAND2X1 U33286 ( .A(n26878), .B(n25918), .Y(n28714) );
  AOI22X1 U33287 ( .A(n28802), .B(reg_A[111]), .C(n26480), .D(n38504), .Y(
        n38500) );
  OAI21X1 U33288 ( .A(n37653), .B(n25546), .C(n38505), .Y(n38504) );
  AOI22X1 U33289 ( .A(n36685), .B(n36666), .C(n25409), .D(n37655), .Y(n38505)
         );
  MUX2X1 U33290 ( .B(n38506), .A(n36170), .S(reg_B[125]), .Y(n36666) );
  INVX1 U33291 ( .A(n36957), .Y(n36685) );
  NAND2X1 U33292 ( .A(reg_B[123]), .B(n36291), .Y(n36957) );
  INVX1 U33293 ( .A(n28592), .Y(n28802) );
  AOI22X1 U33294 ( .A(reg_A[96]), .B(n28590), .C(reg_A[105]), .D(n32528), .Y(
        n38499) );
  INVX1 U33295 ( .A(n28586), .Y(n32528) );
  NOR2X1 U33296 ( .A(n36669), .B(n25138), .Y(n28586) );
  INVX1 U33297 ( .A(n32817), .Y(n25138) );
  NAND2X1 U33298 ( .A(n26927), .B(n25918), .Y(n32817) );
  NOR2X1 U33299 ( .A(n38413), .B(n25279), .Y(n36669) );
  OAI21X1 U33300 ( .A(n38507), .B(n25835), .C(n36614), .Y(n28590) );
  NOR2X1 U33301 ( .A(n28549), .B(n26627), .Y(n36614) );
  INVX1 U33302 ( .A(n31000), .Y(n26627) );
  NAND2X1 U33303 ( .A(n25840), .B(n25222), .Y(n31000) );
  NOR2X1 U33304 ( .A(n29558), .B(n30990), .Y(n28549) );
  AOI21X1 U33305 ( .A(reg_B[1]), .B(n32939), .C(reg_B[0]), .Y(n38507) );
  INVX1 U33306 ( .A(n33395), .Y(n32939) );
  NAND2X1 U33307 ( .A(n38508), .B(n38509), .Y(n38497) );
  NOR2X1 U33308 ( .A(n38510), .B(n38511), .Y(n38509) );
  NAND2X1 U33309 ( .A(n38512), .B(n38513), .Y(n38511) );
  OAI21X1 U33310 ( .A(n38514), .B(n38515), .C(n25560), .Y(n38513) );
  OAI21X1 U33311 ( .A(n38516), .B(n38517), .C(n25310), .Y(n38512) );
  NAND3X1 U33312 ( .A(n38518), .B(n38519), .C(n38520), .Y(n38517) );
  NOR2X1 U33313 ( .A(n38521), .B(n38522), .Y(n38520) );
  OAI22X1 U33314 ( .A(n25043), .B(n25470), .C(n25039), .D(n25493), .Y(n38522)
         );
  OAI21X1 U33315 ( .A(n25064), .B(n36140), .C(n38523), .Y(n38521) );
  AOI22X1 U33316 ( .A(reg_A[121]), .B(n25234), .C(reg_A[122]), .D(n25235), .Y(
        n38523) );
  AOI21X1 U33317 ( .A(reg_A[115]), .B(n25124), .C(n38524), .Y(n38519) );
  OAI22X1 U33318 ( .A(n25037), .B(n25337), .C(n26703), .D(n25476), .Y(n38524)
         );
  AOI22X1 U33319 ( .A(reg_A[118]), .B(n25222), .C(reg_A[117]), .D(n25637), .Y(
        n38518) );
  NAND3X1 U33320 ( .A(n38525), .B(n38526), .C(n38527), .Y(n38516) );
  NOR2X1 U33321 ( .A(n38528), .B(n38529), .Y(n38527) );
  OAI21X1 U33322 ( .A(n25042), .B(n25469), .C(n38530), .Y(n38529) );
  AOI22X1 U33323 ( .A(reg_A[125]), .B(n25241), .C(reg_A[127]), .D(n25339), .Y(
        n38530) );
  OAI21X1 U33324 ( .A(n25038), .B(n25319), .C(n38531), .Y(n38528) );
  AOI22X1 U33325 ( .A(reg_A[124]), .B(n25246), .C(reg_A[123]), .D(n25247), .Y(
        n38531) );
  AOI21X1 U33326 ( .A(reg_A[113]), .B(n25253), .C(n38532), .Y(n38526) );
  OAI22X1 U33327 ( .A(n25040), .B(n25474), .C(n25254), .D(n25450), .Y(n38532)
         );
  AOI22X1 U33328 ( .A(reg_A[114]), .B(n25628), .C(reg_A[111]), .D(n25066), .Y(
        n38525) );
  NAND3X1 U33329 ( .A(n38533), .B(n38534), .C(n38535), .Y(n38510) );
  OAI21X1 U33330 ( .A(n38148), .B(n38536), .C(n25355), .Y(n38535) );
  NAND3X1 U33331 ( .A(n29315), .B(n37993), .C(n38484), .Y(n38534) );
  OAI21X1 U33332 ( .A(n25296), .B(n38382), .C(n38537), .Y(n38484) );
  NAND3X1 U33333 ( .A(n38159), .B(n25521), .C(reg_A[107]), .Y(n38537) );
  NAND2X1 U33334 ( .A(reg_B[110]), .B(n38159), .Y(n38382) );
  OAI21X1 U33335 ( .A(n38538), .B(n38383), .C(n38539), .Y(n38533) );
  INVX1 U33336 ( .A(n25344), .Y(n38539) );
  NOR2X1 U33337 ( .A(n38540), .B(n38541), .Y(n38508) );
  OAI22X1 U33338 ( .A(n25287), .B(n28512), .C(n38542), .D(n38543), .Y(n38541)
         );
  INVX1 U33339 ( .A(n25408), .Y(n38542) );
  NAND2X1 U33340 ( .A(n25607), .B(n25918), .Y(n28512) );
  OAI21X1 U33341 ( .A(n25414), .B(n38544), .C(n38545), .Y(n38540) );
  OAI21X1 U33342 ( .A(n38546), .B(n26626), .C(reg_A[106]), .Y(n38545) );
  INVX1 U33343 ( .A(n26483), .Y(n26626) );
  NOR2X1 U33344 ( .A(n38547), .B(n32880), .Y(n26483) );
  NOR2X1 U33345 ( .A(n25748), .B(n30990), .Y(n32880) );
  AOI22X1 U33346 ( .A(n38159), .B(n38548), .C(n38006), .D(reg_A[111]), .Y(
        n25414) );
  NOR2X1 U33347 ( .A(n38159), .B(n25669), .Y(n38006) );
  NOR2X1 U33348 ( .A(n38549), .B(n38550), .Y(n38495) );
  NAND3X1 U33349 ( .A(n38551), .B(n38552), .C(n38553), .Y(n38550) );
  NOR2X1 U33350 ( .A(n38554), .B(n38555), .Y(n38553) );
  OAI22X1 U33351 ( .A(n28698), .B(n25470), .C(n25994), .D(n38556), .Y(n38555)
         );
  INVX1 U33352 ( .A(n28661), .Y(n28698) );
  NAND2X1 U33353 ( .A(n25145), .B(n38310), .Y(n28661) );
  INVX1 U33354 ( .A(n28835), .Y(n25145) );
  NAND2X1 U33355 ( .A(n36750), .B(n32827), .Y(n28835) );
  NAND2X1 U33356 ( .A(n26924), .B(n25918), .Y(n32827) );
  OAI22X1 U33357 ( .A(n38179), .B(n38420), .C(n28664), .D(n25298), .Y(n38554)
         );
  INVX1 U33358 ( .A(n32603), .Y(n28664) );
  NAND2X1 U33359 ( .A(n26473), .B(n28715), .Y(n32603) );
  NAND2X1 U33360 ( .A(n26804), .B(n25918), .Y(n28715) );
  OAI21X1 U33361 ( .A(n26008), .B(n38557), .C(n38558), .Y(n26473) );
  INVX1 U33362 ( .A(n38559), .Y(n38558) );
  NOR2X1 U33363 ( .A(n33395), .B(n31658), .Y(n38557) );
  NOR2X1 U33364 ( .A(reg_B[2]), .B(n35348), .Y(n33395) );
  NOR2X1 U33365 ( .A(n26863), .B(n26032), .Y(n35348) );
  AOI22X1 U33366 ( .A(n38560), .B(n26756), .C(n38561), .D(n25119), .Y(n38552)
         );
  NAND3X1 U33367 ( .A(n38562), .B(n38563), .C(n38564), .Y(n38561) );
  NOR2X1 U33368 ( .A(n38565), .B(n38566), .Y(n38564) );
  OAI21X1 U33369 ( .A(n26431), .B(n25448), .C(n38567), .Y(n38566) );
  AOI22X1 U33370 ( .A(reg_A[101]), .B(n25253), .C(reg_A[100]), .D(n25628), .Y(
        n38567) );
  OAI21X1 U33371 ( .A(n25040), .B(n25296), .C(n38568), .Y(n38565) );
  AOI22X1 U33372 ( .A(reg_A[106]), .B(n25135), .C(reg_A[104]), .D(n25136), .Y(
        n38568) );
  AOI21X1 U33373 ( .A(reg_A[99]), .B(n25124), .C(n38569), .Y(n38563) );
  OAI22X1 U33374 ( .A(n25037), .B(n25289), .C(n26703), .D(n25361), .Y(n38569)
         );
  AOI22X1 U33375 ( .A(reg_A[97]), .B(n25637), .C(reg_A[107]), .D(n25125), .Y(
        n38562) );
  OAI21X1 U33376 ( .A(n38449), .B(n36136), .C(n38570), .Y(n38560) );
  AOI22X1 U33377 ( .A(n25793), .B(n38571), .C(n25700), .D(n38401), .Y(n38570)
         );
  INVX1 U33378 ( .A(n38389), .Y(n38571) );
  AOI22X1 U33379 ( .A(n37803), .B(n36177), .C(reg_A[103]), .D(n25405), .Y(
        n38389) );
  OAI22X1 U33380 ( .A(n25396), .B(n36318), .C(n25470), .D(n36668), .Y(n37803)
         );
  AOI21X1 U33381 ( .A(n32498), .B(reg_A[100]), .C(n38480), .Y(n38551) );
  INVX1 U33382 ( .A(n28562), .Y(n32498) );
  NAND3X1 U33383 ( .A(n38572), .B(n38573), .C(n38574), .Y(n38549) );
  NOR2X1 U33384 ( .A(n38575), .B(n38576), .Y(n38574) );
  OAI22X1 U33385 ( .A(n38577), .B(n38130), .C(n38343), .D(n38479), .Y(n38576)
         );
  INVX1 U33386 ( .A(n38494), .Y(n38130) );
  OAI21X1 U33387 ( .A(n25820), .B(n25470), .C(n38578), .Y(n38494) );
  AOI22X1 U33388 ( .A(n38347), .B(reg_A[99]), .C(n38107), .D(reg_A[103]), .Y(
        n38578) );
  OAI22X1 U33389 ( .A(n25148), .B(n25469), .C(n28569), .D(n25474), .Y(n38575)
         );
  AOI22X1 U33390 ( .A(reg_A[102]), .B(n25149), .C(n38579), .D(n25150), .Y(
        n38573) );
  INVX1 U33391 ( .A(n26854), .Y(n25150) );
  INVX1 U33392 ( .A(n38325), .Y(n38579) );
  OAI21X1 U33393 ( .A(reg_B[2]), .B(n38063), .C(n38580), .Y(n38325) );
  AOI22X1 U33394 ( .A(n26455), .B(n25424), .C(n26456), .D(n38056), .Y(n38580)
         );
  INVX1 U33395 ( .A(n38581), .Y(n38063) );
  OAI21X1 U33396 ( .A(reg_B[4]), .B(n37823), .C(n38582), .Y(n38581) );
  AOI22X1 U33397 ( .A(n26462), .B(n25468), .C(n26463), .D(n25289), .Y(n38582)
         );
  INVX1 U33398 ( .A(n26861), .Y(n26463) );
  MUX2X1 U33399 ( .B(n25470), .A(n25396), .S(reg_B[1]), .Y(n37823) );
  INVX1 U33400 ( .A(n28571), .Y(n25149) );
  NAND2X1 U33401 ( .A(n25750), .B(n25918), .Y(n28571) );
  AOI22X1 U33402 ( .A(n37984), .B(n25406), .C(reg_A[110]), .D(n25152), .Y(
        n38572) );
  NAND2X1 U33403 ( .A(n38583), .B(n38584), .Y(result[106]) );
  NOR2X1 U33404 ( .A(n38585), .B(n38586), .Y(n38584) );
  NAND2X1 U33405 ( .A(n38587), .B(n38588), .Y(n38586) );
  NOR2X1 U33406 ( .A(n38589), .B(n38590), .Y(n38588) );
  OAI21X1 U33407 ( .A(n38288), .B(n25424), .C(n38591), .Y(n38590) );
  OAI21X1 U33408 ( .A(n38592), .B(n38593), .C(n26480), .Y(n38591) );
  OAI22X1 U33409 ( .A(n38190), .B(n25546), .C(n38594), .D(n25549), .Y(n38593)
         );
  INVX1 U33410 ( .A(n37681), .Y(n38594) );
  OAI22X1 U33411 ( .A(n38595), .B(n36141), .C(n38596), .D(n38597), .Y(n38592)
         );
  INVX1 U33412 ( .A(n38598), .Y(n38288) );
  NAND3X1 U33413 ( .A(n30827), .B(n31636), .C(n38599), .Y(n38598) );
  AOI22X1 U33414 ( .A(n38600), .B(n27676), .C(n25840), .D(n25637), .Y(n38599)
         );
  NOR2X1 U33415 ( .A(n26032), .B(n26596), .Y(n38600) );
  NAND2X1 U33416 ( .A(n37014), .B(reg_B[2]), .Y(n30827) );
  OAI22X1 U33417 ( .A(n38095), .B(n38601), .C(n25450), .D(n28592), .Y(n38589)
         );
  NAND2X1 U33418 ( .A(n25203), .B(n27242), .Y(n28592) );
  INVX1 U33419 ( .A(n38602), .Y(n38601) );
  AOI21X1 U33420 ( .A(n37984), .B(n38108), .C(n38603), .Y(n38587) );
  OAI22X1 U33421 ( .A(n26420), .B(n38193), .C(n38604), .D(n25668), .Y(n38603)
         );
  NAND3X1 U33422 ( .A(n38605), .B(n38606), .C(n38607), .Y(n38585) );
  NOR2X1 U33423 ( .A(n38608), .B(n38609), .Y(n38607) );
  OAI21X1 U33424 ( .A(n38610), .B(n25468), .C(n38611), .Y(n38609) );
  OAI21X1 U33425 ( .A(n38546), .B(n38547), .C(reg_A[105]), .Y(n38611) );
  NOR2X1 U33426 ( .A(n30791), .B(n25279), .Y(n38547) );
  INVX1 U33427 ( .A(n38612), .Y(n38546) );
  NAND3X1 U33428 ( .A(n29315), .B(n38159), .C(n25559), .Y(n38612) );
  NOR2X1 U33429 ( .A(n28343), .B(n38613), .Y(n38610) );
  INVX1 U33430 ( .A(n38310), .Y(n28343) );
  NAND2X1 U33431 ( .A(n25203), .B(n25434), .Y(n38310) );
  INVX1 U33432 ( .A(n25204), .Y(n25434) );
  OAI21X1 U33433 ( .A(n38614), .B(n38615), .C(n38616), .Y(n38608) );
  OAI21X1 U33434 ( .A(n38617), .B(n38618), .C(n25310), .Y(n38616) );
  NAND3X1 U33435 ( .A(n38619), .B(n38620), .C(n38621), .Y(n38618) );
  NOR2X1 U33436 ( .A(n38622), .B(n38623), .Y(n38621) );
  OAI21X1 U33437 ( .A(n25036), .B(n25337), .C(n38624), .Y(n38623) );
  AOI22X1 U33438 ( .A(reg_A[114]), .B(n25124), .C(reg_A[117]), .D(n25222), .Y(
        n38624) );
  OAI21X1 U33439 ( .A(n25037), .B(n25335), .C(n38625), .Y(n38622) );
  AOI22X1 U33440 ( .A(reg_A[110]), .B(n25074), .C(reg_A[111]), .D(n25123), .Y(
        n38625) );
  AOI21X1 U33441 ( .A(reg_A[118]), .B(n25635), .C(n38626), .Y(n38620) );
  OAI22X1 U33442 ( .A(n25065), .B(n25490), .C(n25035), .D(n25493), .Y(n38626)
         );
  AOI22X1 U33443 ( .A(reg_A[119]), .B(n25325), .C(reg_A[106]), .D(n25125), .Y(
        n38619) );
  NAND3X1 U33444 ( .A(n38627), .B(n38628), .C(n38629), .Y(n38617) );
  NOR2X1 U33445 ( .A(n38630), .B(n38631), .Y(n38629) );
  OAI21X1 U33446 ( .A(n26719), .B(n25497), .C(n38632), .Y(n38631) );
  AOI22X1 U33447 ( .A(reg_A[124]), .B(n25241), .C(reg_A[126]), .D(n25339), .Y(
        n38632) );
  OAI21X1 U33448 ( .A(n25038), .B(n25317), .C(n38633), .Y(n38630) );
  AOI22X1 U33449 ( .A(reg_A[123]), .B(n25246), .C(reg_A[122]), .D(n25247), .Y(
        n38633) );
  AOI21X1 U33450 ( .A(reg_A[108]), .B(n25252), .C(n38634), .Y(n38628) );
  OAI22X1 U33451 ( .A(n25041), .B(n25474), .C(n25042), .D(n25470), .Y(n38634)
         );
  AOI22X1 U33452 ( .A(reg_A[112]), .B(n25253), .C(reg_A[113]), .D(n25628), .Y(
        n38627) );
  OR2X1 U33453 ( .A(n38635), .B(n25032), .Y(n38615) );
  AOI22X1 U33454 ( .A(n38147), .B(n28735), .C(n38148), .D(reg_B[126]), .Y(
        n38606) );
  INVX1 U33455 ( .A(n38636), .Y(n38148) );
  INVX1 U33456 ( .A(n26584), .Y(n28735) );
  NAND2X1 U33457 ( .A(n30910), .B(n26452), .Y(n26584) );
  NOR2X1 U33458 ( .A(n38637), .B(n38638), .Y(n38147) );
  OAI22X1 U33459 ( .A(n38639), .B(n27454), .C(n37962), .D(n26599), .Y(n38638)
         );
  MUX2X1 U33460 ( .B(n25468), .A(n25289), .S(reg_B[1]), .Y(n37962) );
  OAI21X1 U33461 ( .A(reg_A[96]), .B(n28739), .C(n38640), .Y(n38637) );
  AOI22X1 U33462 ( .A(n28741), .B(n25448), .C(n28742), .D(n25298), .Y(n38640)
         );
  NOR2X1 U33463 ( .A(n27575), .B(reg_B[1]), .Y(n28742) );
  NOR2X1 U33464 ( .A(n27455), .B(reg_B[1]), .Y(n28741) );
  NAND2X1 U33465 ( .A(reg_B[1]), .B(reg_B[3]), .Y(n28739) );
  AOI22X1 U33466 ( .A(n38641), .B(n25552), .C(n28726), .D(reg_A[111]), .Y(
        n38605) );
  NOR2X1 U33467 ( .A(n30931), .B(n25207), .Y(n28726) );
  INVX1 U33468 ( .A(n38543), .Y(n38641) );
  NOR2X1 U33469 ( .A(n38642), .B(n38643), .Y(n38583) );
  NAND3X1 U33470 ( .A(n38644), .B(n38645), .C(n38646), .Y(n38643) );
  NOR2X1 U33471 ( .A(n38647), .B(n38648), .Y(n38646) );
  OAI21X1 U33472 ( .A(n25521), .B(n38649), .C(n38650), .Y(n38648) );
  OAI21X1 U33473 ( .A(n38651), .B(n38652), .C(n25918), .Y(n38650) );
  OR2X1 U33474 ( .A(n38653), .B(n38654), .Y(n38652) );
  OAI22X1 U33475 ( .A(n25736), .B(n25468), .C(n31398), .D(n25424), .Y(n38654)
         );
  OAI21X1 U33476 ( .A(n27252), .B(n25289), .C(n38655), .Y(n38653) );
  AOI22X1 U33477 ( .A(reg_A[101]), .B(n25750), .C(reg_A[97]), .D(n25614), .Y(
        n38655) );
  OR2X1 U33478 ( .A(n38656), .B(n38657), .Y(n38651) );
  OAI21X1 U33479 ( .A(n26801), .B(n25361), .C(n38658), .Y(n38657) );
  AOI22X1 U33480 ( .A(reg_A[100]), .B(n26878), .C(reg_A[99]), .D(n25613), .Y(
        n38658) );
  OAI21X1 U33481 ( .A(n25062), .B(n25298), .C(n38659), .Y(n38656) );
  AOI22X1 U33482 ( .A(reg_A[105]), .B(n26803), .C(reg_A[103]), .D(n26804), .Y(
        n38659) );
  AOI22X1 U33483 ( .A(n38660), .B(n26756), .C(n38661), .D(n25119), .Y(n38645)
         );
  NAND3X1 U33484 ( .A(n38662), .B(n38663), .C(n38664), .Y(n38661) );
  NOR2X1 U33485 ( .A(n38665), .B(n38666), .Y(n38664) );
  OAI22X1 U33486 ( .A(n25043), .B(n25468), .C(n25467), .D(n25289), .Y(n38666)
         );
  OAI21X1 U33487 ( .A(n25037), .B(n25287), .C(n38667), .Y(n38665) );
  AOI22X1 U33488 ( .A(reg_A[102]), .B(n25074), .C(reg_A[101]), .D(n25123), .Y(
        n38667) );
  AOI21X1 U33489 ( .A(reg_A[104]), .B(n25252), .C(n38668), .Y(n38663) );
  OAI22X1 U33490 ( .A(n25041), .B(n25448), .C(n25042), .D(n25296), .Y(n38668)
         );
  AOI22X1 U33491 ( .A(reg_A[100]), .B(n25253), .C(reg_A[99]), .D(n25628), .Y(
        n38662) );
  OAI21X1 U33492 ( .A(n38669), .B(n36246), .C(n38670), .Y(n38660) );
  AOI22X1 U33493 ( .A(n25793), .B(n38401), .C(n25700), .D(n38671), .Y(n38670)
         );
  OAI22X1 U33494 ( .A(n38189), .B(reg_B[125]), .C(n25544), .D(n25361), .Y(
        n38401) );
  AOI22X1 U33495 ( .A(reg_A[98]), .B(n36686), .C(reg_A[106]), .D(n36338), .Y(
        n38189) );
  AOI22X1 U33496 ( .A(n38328), .B(n25535), .C(n36768), .D(reg_A[104]), .Y(
        n38644) );
  NOR2X1 U33497 ( .A(n38559), .B(n38672), .Y(n36768) );
  OAI21X1 U33498 ( .A(n27358), .B(n26009), .C(n35474), .Y(n38672) );
  NAND3X1 U33499 ( .A(n38673), .B(n38674), .C(n38675), .Y(n38642) );
  AOI21X1 U33500 ( .A(n38676), .B(n38677), .C(n38678), .Y(n38675) );
  OAI22X1 U33501 ( .A(n38179), .B(n38479), .C(n38577), .D(n38420), .Y(n38678)
         );
  INVX1 U33502 ( .A(n38679), .Y(n38420) );
  OAI21X1 U33503 ( .A(n25820), .B(n25468), .C(n38680), .Y(n38679) );
  AOI22X1 U33504 ( .A(n38347), .B(reg_A[98]), .C(n38107), .D(reg_A[102]), .Y(
        n38680) );
  AOI22X1 U33505 ( .A(reg_A[109]), .B(n25152), .C(reg_A[108]), .D(n25153), .Y(
        n38674) );
  INVX1 U33506 ( .A(n28569), .Y(n25153) );
  NAND2X1 U33507 ( .A(n25203), .B(n27243), .Y(n28569) );
  AOI22X1 U33508 ( .A(reg_A[107]), .B(n28280), .C(n25399), .D(n38536), .Y(
        n38673) );
  INVX1 U33509 ( .A(n25148), .Y(n28280) );
  NAND2X1 U33510 ( .A(n25203), .B(n25441), .Y(n25148) );
  NAND2X1 U33511 ( .A(n38681), .B(n38682), .Y(result[105]) );
  NOR2X1 U33512 ( .A(n38683), .B(n38684), .Y(n38682) );
  NAND2X1 U33513 ( .A(n38685), .B(n38686), .Y(n38684) );
  AOI21X1 U33514 ( .A(reg_A[105]), .B(n38613), .C(n38687), .Y(n38686) );
  OAI21X1 U33515 ( .A(n38688), .B(n26864), .C(n38689), .Y(n38687) );
  OAI21X1 U33516 ( .A(n38690), .B(n38691), .C(n25203), .Y(n38689) );
  OAI21X1 U33517 ( .A(n25204), .B(n25296), .C(n38692), .Y(n38691) );
  AOI22X1 U33518 ( .A(reg_A[109]), .B(n27242), .C(reg_A[107]), .D(n27243), .Y(
        n38692) );
  OR2X1 U33519 ( .A(n38693), .B(n38694), .Y(n38690) );
  OAI22X1 U33520 ( .A(n27218), .B(n25468), .C(n25207), .D(n25450), .Y(n38694)
         );
  OAI21X1 U33521 ( .A(n27219), .B(n25452), .C(n38695), .Y(n38693) );
  OAI21X1 U33522 ( .A(n38696), .B(n38697), .C(n25044), .Y(n38695) );
  NAND3X1 U33523 ( .A(n38698), .B(n38699), .C(n38700), .Y(n38697) );
  NOR2X1 U33524 ( .A(n38701), .B(n38702), .Y(n38700) );
  OAI21X1 U33525 ( .A(n25036), .B(n25335), .C(n38703), .Y(n38702) );
  AOI22X1 U33526 ( .A(reg_A[113]), .B(n25124), .C(reg_A[116]), .D(n25222), .Y(
        n38703) );
  OAI21X1 U33527 ( .A(n25037), .B(n25771), .C(n38704), .Y(n38701) );
  AOI22X1 U33528 ( .A(reg_A[109]), .B(n25074), .C(reg_A[110]), .D(n25123), .Y(
        n38704) );
  AOI21X1 U33529 ( .A(reg_A[117]), .B(n25635), .C(n38705), .Y(n38699) );
  OAI22X1 U33530 ( .A(n25065), .B(n25493), .C(n25475), .D(n36140), .Y(n38705)
         );
  AOI22X1 U33531 ( .A(reg_A[118]), .B(n25325), .C(reg_A[105]), .D(n25125), .Y(
        n38698) );
  NAND2X1 U33532 ( .A(n38706), .B(n38707), .Y(n38696) );
  NOR2X1 U33533 ( .A(n38708), .B(n38709), .Y(n38707) );
  OAI21X1 U33534 ( .A(n25238), .B(n25317), .C(n38710), .Y(n38709) );
  AOI22X1 U33535 ( .A(reg_A[123]), .B(n25241), .C(reg_A[127]), .D(n25242), .Y(
        n38710) );
  OAI21X1 U33536 ( .A(n25038), .B(n25323), .C(n38711), .Y(n38708) );
  AOI22X1 U33537 ( .A(reg_A[122]), .B(n25246), .C(reg_A[121]), .D(n25247), .Y(
        n38711) );
  NOR2X1 U33538 ( .A(n38712), .B(n38713), .Y(n38706) );
  OAI21X1 U33539 ( .A(n25030), .B(n25476), .C(n38714), .Y(n38713) );
  AOI22X1 U33540 ( .A(reg_A[107]), .B(n25252), .C(reg_A[111]), .D(n25253), .Y(
        n38714) );
  OAI21X1 U33541 ( .A(n25041), .B(n25469), .C(n38715), .Y(n38712) );
  AOI22X1 U33542 ( .A(reg_A[126]), .B(n25257), .C(reg_A[106]), .D(n25135), .Y(
        n38715) );
  OAI21X1 U33543 ( .A(n25669), .B(n38716), .C(n36750), .Y(n38613) );
  NAND2X1 U33544 ( .A(n30792), .B(n29565), .Y(n36750) );
  NAND2X1 U33545 ( .A(n29315), .B(n38159), .Y(n38716) );
  NAND2X1 U33546 ( .A(n26151), .B(n25031), .Y(n29315) );
  AOI21X1 U33547 ( .A(n37984), .B(n25686), .C(n38717), .Y(n38685) );
  OAI22X1 U33548 ( .A(n26854), .B(n38556), .C(n38604), .D(n25672), .Y(n38717)
         );
  INVX1 U33549 ( .A(n38515), .Y(n38604) );
  OAI22X1 U33550 ( .A(n26151), .B(n38718), .C(n38719), .D(n26147), .Y(n38515)
         );
  NAND2X1 U33551 ( .A(n38720), .B(n38721), .Y(n38556) );
  AOI22X1 U33552 ( .A(n26859), .B(n25436), .C(n26860), .D(n25670), .Y(n38721)
         );
  AND2X1 U33553 ( .A(n26456), .B(n26863), .Y(n26860) );
  AND2X1 U33554 ( .A(n26456), .B(reg_B[4]), .Y(n26859) );
  AOI22X1 U33555 ( .A(n26455), .B(n25424), .C(n38349), .D(n26452), .Y(n38720)
         );
  OAI21X1 U33556 ( .A(reg_A[96]), .B(n26861), .C(n38722), .Y(n38349) );
  AOI22X1 U33557 ( .A(n38723), .B(n26863), .C(n26462), .D(n25298), .Y(n38722)
         );
  NOR2X1 U33558 ( .A(n26863), .B(reg_B[1]), .Y(n26462) );
  INVX1 U33559 ( .A(n38639), .Y(n38723) );
  MUX2X1 U33560 ( .B(n25296), .A(n25287), .S(reg_B[1]), .Y(n38639) );
  NAND2X1 U33561 ( .A(reg_B[1]), .B(reg_B[4]), .Y(n26861) );
  NOR2X1 U33562 ( .A(n26596), .B(n26452), .Y(n26455) );
  NAND2X1 U33563 ( .A(n30910), .B(n26030), .Y(n26854) );
  NAND3X1 U33564 ( .A(n38724), .B(n38725), .C(n38726), .Y(n38683) );
  NOR2X1 U33565 ( .A(n38727), .B(n38728), .Y(n38726) );
  OAI22X1 U33566 ( .A(n26881), .B(n38056), .C(n38729), .D(n38543), .Y(n38728)
         );
  INVX1 U33567 ( .A(n25687), .Y(n38729) );
  NAND2X1 U33568 ( .A(n27443), .B(n26262), .Y(n26881) );
  INVX1 U33569 ( .A(n25994), .Y(n26262) );
  NAND2X1 U33570 ( .A(reg_B[3]), .B(n30910), .Y(n25994) );
  OAI21X1 U33571 ( .A(n25793), .B(n38636), .C(n38730), .Y(n38727) );
  NAND3X1 U33572 ( .A(n25572), .B(n25188), .C(n38538), .Y(n38730) );
  NAND2X1 U33573 ( .A(reg_B[124]), .B(n25357), .Y(n38636) );
  OAI21X1 U33574 ( .A(n38731), .B(n38732), .C(n26480), .Y(n38725) );
  OAI22X1 U33575 ( .A(n38395), .B(n25546), .C(n38733), .D(n25549), .Y(n38732)
         );
  INVX1 U33576 ( .A(n37855), .Y(n38733) );
  OAI22X1 U33577 ( .A(n38734), .B(n36141), .C(n36479), .D(n38597), .Y(n38731)
         );
  INVX1 U33578 ( .A(n36911), .Y(n36479) );
  INVX1 U33579 ( .A(n36877), .Y(n38734) );
  AOI22X1 U33580 ( .A(n38602), .B(n25689), .C(reg_A[96]), .D(n32741), .Y(
        n38724) );
  NAND3X1 U33581 ( .A(n30913), .B(n31636), .C(n38735), .Y(n32741) );
  AOI22X1 U33582 ( .A(n38736), .B(n27676), .C(n25840), .D(n25629), .Y(n38735)
         );
  NOR2X1 U33583 ( .A(n26004), .B(n26596), .Y(n38736) );
  NAND2X1 U33584 ( .A(n27676), .B(reg_B[0]), .Y(n31636) );
  NAND2X1 U33585 ( .A(n37014), .B(reg_B[3]), .Y(n30913) );
  NOR2X1 U33586 ( .A(n38737), .B(n38738), .Y(n38681) );
  NAND3X1 U33587 ( .A(n38739), .B(n38740), .C(n38741), .Y(n38738) );
  AOI21X1 U33588 ( .A(n38514), .B(n25669), .C(n38742), .Y(n38741) );
  OAI21X1 U33589 ( .A(n38743), .B(n38083), .C(n38744), .Y(n38742) );
  OAI21X1 U33590 ( .A(n38745), .B(n38746), .C(n25119), .Y(n38744) );
  NAND2X1 U33591 ( .A(n38747), .B(n38748), .Y(n38746) );
  AOI22X1 U33592 ( .A(reg_A[101]), .B(n25074), .C(reg_A[100]), .D(n25123), .Y(
        n38748) );
  AOI22X1 U33593 ( .A(reg_A[97]), .B(n25124), .C(reg_A[105]), .D(n25125), .Y(
        n38747) );
  OR2X1 U33594 ( .A(n38749), .B(n38750), .Y(n38745) );
  OAI22X1 U33595 ( .A(n25030), .B(n25289), .C(n25033), .D(n25396), .Y(n38750)
         );
  OAI21X1 U33596 ( .A(n25040), .B(n25448), .C(n38751), .Y(n38749) );
  AOI22X1 U33597 ( .A(reg_A[104]), .B(n25135), .C(reg_A[102]), .D(n25136), .Y(
        n38751) );
  INVX1 U33598 ( .A(n38328), .Y(n38083) );
  INVX1 U33599 ( .A(n25673), .Y(n38743) );
  INVX1 U33600 ( .A(n38649), .Y(n38514) );
  INVX1 U33601 ( .A(n38647), .Y(n38740) );
  OAI21X1 U33602 ( .A(n38752), .B(n38753), .C(n38754), .Y(n38647) );
  INVX1 U33603 ( .A(n38480), .Y(n38754) );
  OAI21X1 U33604 ( .A(n27438), .B(n38050), .C(n38755), .Y(n38480) );
  NOR2X1 U33605 ( .A(n38326), .B(n38327), .Y(n38755) );
  INVX1 U33606 ( .A(n37927), .Y(n38327) );
  NAND2X1 U33607 ( .A(n37006), .B(n25932), .Y(n37927) );
  INVX1 U33608 ( .A(n37635), .Y(n37006) );
  NAND2X1 U33609 ( .A(reg_B[123]), .B(reg_A[96]), .Y(n37635) );
  AND2X1 U33610 ( .A(reg_B[109]), .B(n38756), .Y(n38326) );
  OAI21X1 U33611 ( .A(n25032), .B(n38752), .C(n38649), .Y(n38756) );
  NAND2X1 U33612 ( .A(reg_A[104]), .B(n26504), .Y(n38649) );
  NAND2X1 U33613 ( .A(n36240), .B(reg_A[96]), .Y(n38050) );
  NOR2X1 U33614 ( .A(n36291), .B(n36177), .Y(n36240) );
  NAND2X1 U33615 ( .A(reg_B[110]), .B(n25188), .Y(n38753) );
  AOI22X1 U33616 ( .A(n34606), .B(reg_A[104]), .C(n25918), .D(n38757), .Y(
        n38739) );
  NAND3X1 U33617 ( .A(n38758), .B(n38759), .C(n38760), .Y(n38757) );
  NOR2X1 U33618 ( .A(n38761), .B(n38762), .Y(n38760) );
  OAI22X1 U33619 ( .A(n26800), .B(n25436), .C(n26801), .D(n25670), .Y(n38762)
         );
  OAI21X1 U33620 ( .A(n25062), .B(n25448), .C(n38763), .Y(n38761) );
  AOI22X1 U33621 ( .A(reg_A[104]), .B(n26803), .C(reg_A[102]), .D(n26804), .Y(
        n38763) );
  AOI22X1 U33622 ( .A(reg_A[96]), .B(n25614), .C(reg_A[97]), .D(n25615), .Y(
        n38759) );
  INVX1 U33623 ( .A(n38764), .Y(n38758) );
  OAI21X1 U33624 ( .A(n25296), .B(n25736), .C(n38688), .Y(n38764) );
  AOI22X1 U33625 ( .A(n25613), .B(reg_A[98]), .C(n26878), .D(reg_A[99]), .Y(
        n38688) );
  NOR2X1 U33626 ( .A(n38559), .B(n38765), .Y(n34606) );
  OAI21X1 U33627 ( .A(n27358), .B(n26007), .C(n26943), .Y(n38765) );
  NAND2X1 U33628 ( .A(n25029), .B(n29565), .Y(n38559) );
  NAND3X1 U33629 ( .A(n38766), .B(n38767), .C(n38768), .Y(n38737) );
  AOI21X1 U33630 ( .A(n38769), .B(n26756), .C(n38770), .Y(n38768) );
  OAI22X1 U33631 ( .A(n38771), .B(n38131), .C(n38577), .D(n38479), .Y(n38770)
         );
  INVX1 U33632 ( .A(n38772), .Y(n38479) );
  OAI21X1 U33633 ( .A(n25820), .B(n25296), .C(n38773), .Y(n38772) );
  AOI22X1 U33634 ( .A(n38347), .B(reg_A[97]), .C(n38107), .D(reg_A[101]), .Y(
        n38773) );
  INVX1 U33635 ( .A(n38676), .Y(n38131) );
  OAI21X1 U33636 ( .A(n38774), .B(n36246), .C(n38775), .Y(n38769) );
  AOI22X1 U33637 ( .A(n25793), .B(n38671), .C(n25399), .D(n38776), .Y(n38775)
         );
  INVX1 U33638 ( .A(n38449), .Y(n38671) );
  AOI22X1 U33639 ( .A(n38012), .B(n36177), .C(n25405), .D(reg_A[101]), .Y(
        n38449) );
  OAI22X1 U33640 ( .A(n25287), .B(n36318), .C(n25296), .D(n36668), .Y(n38012)
         );
  AOI22X1 U33641 ( .A(reg_A[108]), .B(n25152), .C(n38383), .D(n25696), .Y(
        n38767) );
  INVX1 U33642 ( .A(n28570), .Y(n25152) );
  NAND2X1 U33643 ( .A(n25203), .B(n27241), .Y(n28570) );
  AOI22X1 U33644 ( .A(n25700), .B(n38536), .C(n37986), .D(n38677), .Y(n38766)
         );
  NAND3X1 U33645 ( .A(n38777), .B(n38778), .C(n38779), .Y(result[104]) );
  NOR2X1 U33646 ( .A(n38780), .B(n38781), .Y(n38779) );
  NAND3X1 U33647 ( .A(n38782), .B(n38783), .C(n38784), .Y(n38781) );
  AOI21X1 U33648 ( .A(n38785), .B(n28575), .C(n38786), .Y(n38784) );
  OAI21X1 U33649 ( .A(n32872), .B(n25424), .C(n38787), .Y(n38786) );
  OAI21X1 U33650 ( .A(n38788), .B(n38789), .C(n25730), .Y(n38787) );
  OAI21X1 U33651 ( .A(n26800), .B(n25474), .C(n38790), .Y(n38789) );
  AOI22X1 U33652 ( .A(reg_A[111]), .B(n25613), .C(reg_A[108]), .D(n25749), .Y(
        n38790) );
  NAND2X1 U33653 ( .A(n38791), .B(n38792), .Y(n38788) );
  AOI22X1 U33654 ( .A(reg_A[105]), .B(n26803), .C(reg_A[107]), .D(n26804), .Y(
        n38792) );
  AOI22X1 U33655 ( .A(reg_A[106]), .B(n26927), .C(reg_A[110]), .D(n26878), .Y(
        n38791) );
  INVX1 U33656 ( .A(n38793), .Y(n32872) );
  OAI21X1 U33657 ( .A(n26664), .B(n25835), .C(n38794), .Y(n38793) );
  AOI21X1 U33658 ( .A(n25840), .B(n25124), .C(n37014), .Y(n38794) );
  INVX1 U33659 ( .A(n26985), .Y(n37014) );
  NAND2X1 U33660 ( .A(reg_B[1]), .B(n30910), .Y(n26985) );
  INVX1 U33661 ( .A(n26420), .Y(n28575) );
  NAND2X1 U33662 ( .A(n26456), .B(n30910), .Y(n26420) );
  NOR2X1 U33663 ( .A(n26452), .B(reg_B[1]), .Y(n26456) );
  OAI21X1 U33664 ( .A(n38795), .B(n38796), .C(n26480), .Y(n38783) );
  OAI22X1 U33665 ( .A(n38416), .B(n25546), .C(n38490), .D(n25549), .Y(n38796)
         );
  INVX1 U33666 ( .A(n37882), .Y(n38490) );
  OAI22X1 U33667 ( .A(n36986), .B(n36141), .C(n38797), .D(n38597), .Y(n38795)
         );
  NAND2X1 U33668 ( .A(reg_B[123]), .B(n36355), .Y(n38597) );
  INVX1 U33669 ( .A(n36619), .Y(n38797) );
  NAND2X1 U33670 ( .A(reg_B[123]), .B(n36356), .Y(n36141) );
  INVX1 U33671 ( .A(n37883), .Y(n36986) );
  AOI22X1 U33672 ( .A(n38492), .B(n27008), .C(n38538), .D(n38798), .Y(n38782)
         );
  INVX1 U33673 ( .A(n26729), .Y(n27008) );
  NAND2X1 U33674 ( .A(n27443), .B(n30910), .Y(n26729) );
  INVX1 U33675 ( .A(n27857), .Y(n27443) );
  NAND2X1 U33676 ( .A(n26596), .B(n26452), .Y(n27857) );
  AND2X1 U33677 ( .A(n38799), .B(n38800), .Y(n38492) );
  AOI22X1 U33678 ( .A(n26601), .B(n25361), .C(n26602), .D(n25670), .Y(n38800)
         );
  AOI22X1 U33679 ( .A(n27012), .B(n25298), .C(n26597), .D(n25448), .Y(n38799)
         );
  NAND3X1 U33680 ( .A(n38801), .B(n38802), .C(n38803), .Y(n38780) );
  AOI21X1 U33681 ( .A(n38602), .B(n25825), .C(n38804), .Y(n38803) );
  OAI22X1 U33682 ( .A(n25810), .B(n38543), .C(n38719), .D(n38805), .Y(n38804)
         );
  AOI21X1 U33683 ( .A(reg_A[96]), .B(n38347), .C(n38538), .Y(n38719) );
  INVX1 U33684 ( .A(n38614), .Y(n38538) );
  NAND2X1 U33685 ( .A(n38467), .B(n38806), .Y(n38614) );
  OAI21X1 U33686 ( .A(n38159), .B(n25436), .C(n38718), .Y(n38806) );
  NAND2X1 U33687 ( .A(n25393), .B(n25382), .Y(n38543) );
  INVX1 U33688 ( .A(n38807), .Y(n25810) );
  NOR2X1 U33689 ( .A(n38544), .B(n38159), .Y(n38602) );
  OAI21X1 U33690 ( .A(n36973), .B(n38808), .C(reg_A[104]), .Y(n38802) );
  INVX1 U33691 ( .A(n32826), .Y(n38808) );
  NAND2X1 U33692 ( .A(n38809), .B(n25029), .Y(n32826) );
  AOI22X1 U33693 ( .A(n33724), .B(n26943), .C(n25279), .D(n25517), .Y(n38809)
         );
  INVX1 U33694 ( .A(n25372), .Y(n25517) );
  INVX1 U33695 ( .A(n29565), .Y(n25279) );
  NAND2X1 U33696 ( .A(n27523), .B(n31658), .Y(n29565) );
  AOI21X1 U33697 ( .A(n38810), .B(n38811), .C(n38812), .Y(n38801) );
  INVX1 U33698 ( .A(n38718), .Y(n38811) );
  NAND2X1 U33699 ( .A(reg_A[104]), .B(n38159), .Y(n38718) );
  NOR2X1 U33700 ( .A(n26151), .B(n25669), .Y(n38810) );
  NOR2X1 U33701 ( .A(n38813), .B(n38814), .Y(n38778) );
  OAI21X1 U33702 ( .A(n25198), .B(n38815), .C(n38816), .Y(n38814) );
  AOI22X1 U33703 ( .A(n38493), .B(n38677), .C(n38676), .D(n38817), .Y(n38816)
         );
  OAI21X1 U33704 ( .A(n26147), .B(n25671), .C(n25344), .Y(n38676) );
  NAND2X1 U33705 ( .A(n25696), .B(reg_B[110]), .Y(n25344) );
  INVX1 U33706 ( .A(n38179), .Y(n38493) );
  AOI22X1 U33707 ( .A(n26267), .B(n25559), .C(n25188), .D(n25572), .Y(n38179)
         );
  AOI21X1 U33708 ( .A(n25355), .B(n38818), .C(n38819), .Y(n38815) );
  OAI22X1 U33709 ( .A(n38774), .B(n36136), .C(n38669), .D(n25568), .Y(n38819)
         );
  INVX1 U33710 ( .A(n38776), .Y(n38669) );
  INVX1 U33711 ( .A(n38820), .Y(n38774) );
  OAI21X1 U33712 ( .A(n38771), .B(n38343), .C(n38821), .Y(n38813) );
  AOI22X1 U33713 ( .A(n37984), .B(n38822), .C(n25793), .D(n38536), .Y(n38821)
         );
  OAI21X1 U33714 ( .A(n38823), .B(n27438), .C(n38824), .Y(n38536) );
  OAI21X1 U33715 ( .A(n38825), .B(n38826), .C(n25699), .Y(n38824) );
  NOR2X1 U33716 ( .A(reg_B[125]), .B(n38109), .Y(n38825) );
  AOI22X1 U33717 ( .A(reg_A[96]), .B(n36686), .C(reg_A[104]), .D(n36338), .Y(
        n38109) );
  AOI21X1 U33718 ( .A(reg_A[104]), .B(n25427), .C(n38826), .Y(n38823) );
  NOR2X1 U33719 ( .A(n25436), .B(n25544), .Y(n38826) );
  INVX1 U33720 ( .A(n37986), .Y(n38343) );
  OAI22X1 U33721 ( .A(n26147), .B(n25668), .C(n25794), .D(n38635), .Y(n37986)
         );
  NOR2X1 U33722 ( .A(n38827), .B(n38828), .Y(n38777) );
  OAI21X1 U33723 ( .A(n25794), .B(n38752), .C(n38829), .Y(n38828) );
  AOI22X1 U33724 ( .A(n25918), .B(n38830), .C(n25310), .D(n38831), .Y(n38829)
         );
  NAND3X1 U33725 ( .A(n38832), .B(n38833), .C(n38834), .Y(n38831) );
  AND2X1 U33726 ( .A(n38835), .B(n38836), .Y(n38834) );
  NOR2X1 U33727 ( .A(n38837), .B(n38838), .Y(n38836) );
  OAI21X1 U33728 ( .A(n25050), .B(n25497), .C(n38839), .Y(n38838) );
  AOI22X1 U33729 ( .A(reg_A[122]), .B(n25241), .C(reg_A[126]), .D(n25242), .Y(
        n38839) );
  OAI21X1 U33730 ( .A(n25038), .B(n25321), .C(n38840), .Y(n38837) );
  AOI22X1 U33731 ( .A(reg_A[121]), .B(n25246), .C(reg_A[120]), .D(n25247), .Y(
        n38840) );
  NOR2X1 U33732 ( .A(n38841), .B(n38842), .Y(n38835) );
  OAI21X1 U33733 ( .A(n25033), .B(n25450), .C(n38843), .Y(n38842) );
  AOI22X1 U33734 ( .A(reg_A[107]), .B(n25136), .C(reg_A[106]), .D(n25252), .Y(
        n38843) );
  OAI21X1 U33735 ( .A(n25042), .B(n25296), .C(n38844), .Y(n38841) );
  AOI22X1 U33736 ( .A(reg_A[124]), .B(n25339), .C(reg_A[125]), .D(n25257), .Y(
        n38844) );
  NOR2X1 U33737 ( .A(n38845), .B(n38846), .Y(n38833) );
  OAI21X1 U33738 ( .A(n25027), .B(n25335), .C(n38847), .Y(n38846) );
  AOI22X1 U33739 ( .A(reg_A[113]), .B(n25629), .C(reg_A[112]), .D(n25124), .Y(
        n38847) );
  OAI21X1 U33740 ( .A(n25028), .B(n25474), .C(n38848), .Y(n38845) );
  AOI22X1 U33741 ( .A(reg_A[111]), .B(n25628), .C(reg_A[108]), .D(n25066), .Y(
        n38848) );
  NOR2X1 U33742 ( .A(n38849), .B(n38850), .Y(n38832) );
  OAI21X1 U33743 ( .A(n25043), .B(n25298), .C(n38851), .Y(n38850) );
  AOI22X1 U33744 ( .A(reg_A[116]), .B(n25635), .C(reg_A[117]), .D(n25325), .Y(
        n38851) );
  OAI21X1 U33745 ( .A(n25065), .B(n36140), .C(n38852), .Y(n38849) );
  AOI22X1 U33746 ( .A(reg_A[114]), .B(n25637), .C(reg_A[118]), .D(n25234), .Y(
        n38852) );
  NAND3X1 U33747 ( .A(n38853), .B(n38854), .C(n38855), .Y(n38830) );
  NOR2X1 U33748 ( .A(n38856), .B(n38857), .Y(n38855) );
  OAI22X1 U33749 ( .A(n26936), .B(n25287), .C(n25745), .D(n25289), .Y(n38857)
         );
  OAI21X1 U33750 ( .A(n25062), .B(n25361), .C(n38858), .Y(n38856) );
  AOI22X1 U33751 ( .A(reg_A[103]), .B(n26803), .C(reg_A[101]), .D(n26804), .Y(
        n38858) );
  AOI22X1 U33752 ( .A(reg_A[100]), .B(n25749), .C(reg_A[99]), .D(n25750), .Y(
        n38854) );
  AOI22X1 U33753 ( .A(reg_A[96]), .B(n25615), .C(reg_A[104]), .D(n26924), .Y(
        n38853) );
  NAND2X1 U33754 ( .A(n38859), .B(n38860), .Y(n38827) );
  OAI21X1 U33755 ( .A(n38861), .B(n38862), .C(n26928), .Y(n38860) );
  NAND2X1 U33756 ( .A(n38863), .B(n38864), .Y(n38862) );
  AOI22X1 U33757 ( .A(reg_A[111]), .B(n26002), .C(reg_A[108]), .D(n26003), .Y(
        n38864) );
  AOI22X1 U33758 ( .A(reg_A[109]), .B(n25751), .C(reg_A[104]), .D(n26004), .Y(
        n38863) );
  NAND2X1 U33759 ( .A(n38865), .B(n38866), .Y(n38861) );
  AOI22X1 U33760 ( .A(reg_A[105]), .B(n26007), .C(reg_A[107]), .D(n26008), .Y(
        n38866) );
  AOI22X1 U33761 ( .A(reg_A[106]), .B(n26009), .C(reg_A[110]), .D(n26010), .Y(
        n38865) );
  AOI22X1 U33762 ( .A(n38867), .B(n25119), .C(n38328), .D(n25803), .Y(n38859)
         );
  NOR2X1 U33763 ( .A(n38544), .B(reg_B[109]), .Y(n38328) );
  NAND2X1 U33764 ( .A(n25382), .B(n38084), .Y(n38544) );
  OAI21X1 U33765 ( .A(reg_B[108]), .B(n25415), .C(n26999), .Y(n38084) );
  NAND3X1 U33766 ( .A(n38868), .B(n38869), .C(n38870), .Y(n38867) );
  NOR2X1 U33767 ( .A(n38871), .B(n38872), .Y(n38870) );
  OAI22X1 U33768 ( .A(n25033), .B(n25289), .C(n25040), .D(n25361), .Y(n38872)
         );
  OAI22X1 U33769 ( .A(n25041), .B(n25670), .C(n25042), .D(n25448), .Y(n38871)
         );
  AOI22X1 U33770 ( .A(reg_A[97]), .B(n25628), .C(reg_A[100]), .D(n25066), .Y(
        n38869) );
  AOI22X1 U33771 ( .A(reg_A[99]), .B(n25123), .C(reg_A[104]), .D(n25125), .Y(
        n38868) );
  OR2X1 U33772 ( .A(n38873), .B(n38874), .Y(result[103]) );
  NAND3X1 U33773 ( .A(n38875), .B(n38876), .C(n38877), .Y(n38874) );
  NOR2X1 U33774 ( .A(n38878), .B(n38879), .Y(n38877) );
  OAI21X1 U33775 ( .A(n38880), .B(n27438), .C(n38881), .Y(n38879) );
  AOI22X1 U33776 ( .A(reg_A[110]), .B(n25293), .C(n25170), .D(n38882), .Y(
        n38881) );
  NAND3X1 U33777 ( .A(n38883), .B(n38884), .C(n38885), .Y(n38882) );
  AOI21X1 U33778 ( .A(n25379), .B(n38886), .C(n38887), .Y(n38885) );
  OAI22X1 U33779 ( .A(n38888), .B(n25656), .C(n25448), .D(n25711), .Y(n38887)
         );
  INVX1 U33780 ( .A(n38677), .Y(n38888) );
  AOI22X1 U33781 ( .A(n38889), .B(n38890), .C(n25097), .D(n38891), .Y(n38884)
         );
  OAI21X1 U33782 ( .A(n38892), .B(n36246), .C(n38880), .Y(n38891) );
  INVX1 U33783 ( .A(n38893), .Y(n38890) );
  AOI22X1 U33784 ( .A(reg_A[99]), .B(n38894), .C(reg_A[97]), .D(n38895), .Y(
        n38893) );
  AOI22X1 U33785 ( .A(n25604), .B(n38896), .C(n25822), .D(reg_A[101]), .Y(
        n38883) );
  INVX1 U33786 ( .A(n38897), .Y(n25822) );
  OAI21X1 U33787 ( .A(n38898), .B(n25671), .C(n38899), .Y(n38896) );
  AOI22X1 U33788 ( .A(n25559), .B(n38900), .C(n25562), .D(n38817), .Y(n38899)
         );
  OAI22X1 U33789 ( .A(n25030), .B(n26990), .C(n26936), .D(n27152), .Y(n25293)
         );
  INVX1 U33790 ( .A(n38901), .Y(n38880) );
  OAI21X1 U33791 ( .A(n38902), .B(n36136), .C(n38903), .Y(n38901) );
  AOI22X1 U33792 ( .A(n25793), .B(n38776), .C(n25700), .D(n38820), .Y(n38903)
         );
  OAI22X1 U33793 ( .A(n25396), .B(n25544), .C(n25356), .D(n25448), .Y(n38776)
         );
  OAI21X1 U33794 ( .A(n25295), .B(n25474), .C(n38904), .Y(n38878) );
  AOI22X1 U33795 ( .A(reg_A[107]), .B(n29029), .C(reg_A[108]), .D(n29030), .Y(
        n38904) );
  OAI22X1 U33796 ( .A(n25028), .B(n26990), .C(n26800), .D(n27152), .Y(n29030)
         );
  OAI22X1 U33797 ( .A(n26431), .B(n26990), .C(n26801), .D(n27152), .Y(n29029)
         );
  INVX1 U33798 ( .A(n29031), .Y(n25295) );
  OAI22X1 U33799 ( .A(n25033), .B(n26990), .C(n25745), .D(n27152), .Y(n29031)
         );
  NOR2X1 U33800 ( .A(n38905), .B(n38906), .Y(n38876) );
  OAI21X1 U33801 ( .A(n29036), .B(n25298), .C(n38907), .Y(n38906) );
  OAI21X1 U33802 ( .A(n38908), .B(n38909), .C(n25310), .Y(n38907) );
  NAND3X1 U33803 ( .A(n38910), .B(n38911), .C(n38912), .Y(n38909) );
  NOR2X1 U33804 ( .A(n38913), .B(n38914), .Y(n38912) );
  OAI22X1 U33805 ( .A(n25036), .B(n25483), .C(n25473), .D(n25771), .Y(n38914)
         );
  OAI22X1 U33806 ( .A(n25037), .B(n25476), .C(n25320), .D(n25497), .Y(n38913)
         );
  AOI22X1 U33807 ( .A(reg_A[117]), .B(n25234), .C(reg_A[118]), .D(n25235), .Y(
        n38911) );
  AOI22X1 U33808 ( .A(reg_A[115]), .B(n25635), .C(reg_A[116]), .D(n25325), .Y(
        n38910) );
  NAND3X1 U33809 ( .A(n38915), .B(n38916), .C(n38917), .Y(n38908) );
  NOR2X1 U33810 ( .A(n38918), .B(n38919), .Y(n38917) );
  OAI22X1 U33811 ( .A(n25331), .B(n25490), .C(n25038), .D(n25494), .Y(n38919)
         );
  OAI22X1 U33812 ( .A(n25334), .B(n36140), .C(n25336), .D(n25493), .Y(n38918)
         );
  INVX1 U33813 ( .A(reg_A[120]), .Y(n25493) );
  INVX1 U33814 ( .A(reg_A[119]), .Y(n36140) );
  AOI22X1 U33815 ( .A(reg_A[125]), .B(n25242), .C(reg_A[126]), .D(n25338), .Y(
        n38916) );
  AOI22X1 U33816 ( .A(reg_A[123]), .B(n25339), .C(reg_A[124]), .D(n25257), .Y(
        n38915) );
  INVX1 U33817 ( .A(n27940), .Y(n29036) );
  OAI22X1 U33818 ( .A(n25042), .B(n26990), .C(n25748), .D(n27152), .Y(n27940)
         );
  OAI22X1 U33819 ( .A(n25945), .B(n38920), .C(n27964), .D(n25448), .Y(n38905)
         );
  INVX1 U33820 ( .A(n33034), .Y(n27964) );
  OAI21X1 U33821 ( .A(n26943), .B(n37184), .C(n32946), .Y(n33034) );
  INVX1 U33822 ( .A(n25283), .Y(n32946) );
  NAND2X1 U33823 ( .A(n35065), .B(n33195), .Y(n25283) );
  AOI21X1 U33824 ( .A(n25125), .B(n25310), .C(n29546), .Y(n35065) );
  INVX1 U33825 ( .A(n25795), .Y(n29546) );
  NAND2X1 U33826 ( .A(n30427), .B(reg_B[3]), .Y(n25945) );
  AOI21X1 U33827 ( .A(reg_A[106]), .B(n29051), .C(n38921), .Y(n38875) );
  OAI22X1 U33828 ( .A(n27938), .B(n25296), .C(n27512), .D(n25452), .Y(n38921)
         );
  INVX1 U33829 ( .A(n25302), .Y(n27512) );
  OAI22X1 U33830 ( .A(n25034), .B(n26990), .C(n27252), .D(n27152), .Y(n25302)
         );
  INVX1 U33831 ( .A(n37015), .Y(n27938) );
  OAI22X1 U33832 ( .A(n25040), .B(n26990), .C(n25746), .D(n27152), .Y(n37015)
         );
  INVX1 U33833 ( .A(n27968), .Y(n29051) );
  AOI22X1 U33834 ( .A(n25136), .B(n25310), .C(n26804), .D(n25730), .Y(n27968)
         );
  NAND3X1 U33835 ( .A(n38922), .B(n38923), .C(n38924), .Y(n38873) );
  NOR2X1 U33836 ( .A(n38925), .B(n38926), .Y(n38924) );
  OAI21X1 U33837 ( .A(n28053), .B(n38056), .C(n38927), .Y(n38926) );
  AOI22X1 U33838 ( .A(reg_A[100]), .B(n38928), .C(n38929), .D(n37958), .Y(
        n38927) );
  OAI21X1 U33839 ( .A(n25519), .B(n38387), .C(n27095), .Y(n38928) );
  NAND2X1 U33840 ( .A(n25999), .B(n26008), .Y(n27095) );
  MUX2X1 U33841 ( .B(reg_A[102]), .A(reg_A[103]), .S(n26863), .Y(n38056) );
  NAND2X1 U33842 ( .A(n30427), .B(n26032), .Y(n28053) );
  NAND3X1 U33843 ( .A(n38930), .B(n38931), .C(n38932), .Y(n38925) );
  AOI21X1 U33844 ( .A(n38933), .B(reg_B[125]), .C(n38812), .Y(n38932) );
  NOR2X1 U33845 ( .A(n38934), .B(n36246), .Y(n38933) );
  OAI21X1 U33846 ( .A(n38935), .B(n38936), .C(n27067), .Y(n38931) );
  NAND2X1 U33847 ( .A(n26864), .B(n30990), .Y(n27067) );
  OAI21X1 U33848 ( .A(n25060), .B(n25448), .C(n38937), .Y(n38936) );
  AOI22X1 U33849 ( .A(reg_A[99]), .B(n25749), .C(reg_A[98]), .D(n25750), .Y(
        n38937) );
  NAND2X1 U33850 ( .A(n38938), .B(n38939), .Y(n38935) );
  AOI22X1 U33851 ( .A(reg_A[102]), .B(n26803), .C(reg_A[100]), .D(n26804), .Y(
        n38939) );
  AOI22X1 U33852 ( .A(reg_A[101]), .B(n26927), .C(reg_A[97]), .D(n26878), .Y(
        n38938) );
  OAI21X1 U33853 ( .A(n38940), .B(n38941), .C(n25119), .Y(n38930) );
  NAND2X1 U33854 ( .A(n25835), .B(n30951), .Y(n25119) );
  OAI21X1 U33855 ( .A(n25043), .B(n25448), .C(n38942), .Y(n38941) );
  AOI22X1 U33856 ( .A(reg_A[99]), .B(n25075), .C(reg_A[98]), .D(n25123), .Y(
        n38942) );
  NAND2X1 U33857 ( .A(n38943), .B(n38944), .Y(n38940) );
  AOI22X1 U33858 ( .A(reg_A[102]), .B(n25135), .C(reg_A[100]), .D(n25136), .Y(
        n38944) );
  AOI22X1 U33859 ( .A(reg_A[101]), .B(n25252), .C(reg_A[97]), .D(n25253), .Y(
        n38943) );
  NOR2X1 U33860 ( .A(n38945), .B(n38946), .Y(n38923) );
  OAI21X1 U33861 ( .A(n25289), .B(n27108), .C(n38947), .Y(n38946) );
  NAND2X1 U33862 ( .A(n25999), .B(n38948), .Y(n38947) );
  OAI21X1 U33863 ( .A(n25754), .B(n25287), .C(n38949), .Y(n38948) );
  AOI22X1 U33864 ( .A(reg_A[102]), .B(n26007), .C(reg_A[101]), .D(n26009), .Y(
        n38949) );
  INVX1 U33865 ( .A(n37184), .Y(n25999) );
  NAND2X1 U33866 ( .A(n25751), .B(n38950), .Y(n27108) );
  OAI21X1 U33867 ( .A(n38951), .B(n25342), .C(n38952), .Y(n38945) );
  OAI21X1 U33868 ( .A(n38953), .B(n38954), .C(n25188), .Y(n38952) );
  OAI21X1 U33869 ( .A(n38955), .B(n25671), .C(n38752), .Y(n38954) );
  OAI21X1 U33870 ( .A(n38956), .B(n38635), .C(n38957), .Y(n38953) );
  AOI22X1 U33871 ( .A(n25572), .B(n38900), .C(n25709), .D(n38677), .Y(n38957)
         );
  OAI22X1 U33872 ( .A(n25396), .B(n38003), .C(n25820), .D(n25448), .Y(n38677)
         );
  NOR2X1 U33873 ( .A(n38958), .B(reg_B[110]), .Y(n25572) );
  NAND2X1 U33874 ( .A(n38959), .B(reg_B[110]), .Y(n38635) );
  AOI21X1 U33875 ( .A(n38960), .B(reg_B[102]), .C(n38961), .Y(n38951) );
  MUX2X1 U33876 ( .B(n38962), .A(n38963), .S(reg_B[103]), .Y(n38961) );
  AOI22X1 U33877 ( .A(n38894), .B(reg_A[99]), .C(reg_A[103]), .D(n25574), .Y(
        n38962) );
  AOI21X1 U33878 ( .A(reg_A[96]), .B(n28055), .C(n38964), .Y(n38922) );
  OAI21X1 U33879 ( .A(n25396), .B(n27995), .C(n38965), .Y(n38964) );
  OAI21X1 U33880 ( .A(n38966), .B(n38967), .C(n25382), .Y(n38965) );
  OAI21X1 U33881 ( .A(n25448), .B(n25711), .C(n38968), .Y(n38967) );
  AOI22X1 U33882 ( .A(n25393), .B(n25404), .C(n25571), .D(n25389), .Y(n38968)
         );
  NAND2X1 U33883 ( .A(n38969), .B(n38970), .Y(n25389) );
  AOI22X1 U33884 ( .A(reg_A[104]), .B(n25559), .C(reg_A[106]), .D(n25560), .Y(
        n38970) );
  AOI22X1 U33885 ( .A(reg_A[103]), .B(n25561), .C(reg_A[105]), .D(n25562), .Y(
        n38969) );
  INVX1 U33886 ( .A(n38971), .Y(n25571) );
  NAND2X1 U33887 ( .A(n38972), .B(n38973), .Y(n25404) );
  AOI22X1 U33888 ( .A(reg_A[106]), .B(n25355), .C(reg_A[105]), .D(n25399), .Y(
        n38973) );
  AOI22X1 U33889 ( .A(n25793), .B(reg_A[103]), .C(reg_A[104]), .D(n25700), .Y(
        n38972) );
  OAI21X1 U33890 ( .A(n38974), .B(n25558), .C(n38975), .Y(n38966) );
  AOI22X1 U33891 ( .A(n38976), .B(n38347), .C(n25097), .D(n38977), .Y(n38975)
         );
  NAND2X1 U33892 ( .A(n38978), .B(n38979), .Y(n38977) );
  AOI22X1 U33893 ( .A(n25405), .B(n25408), .C(n25407), .D(n37655), .Y(n38979)
         );
  NAND2X1 U33894 ( .A(n38980), .B(n38981), .Y(n37655) );
  AOI22X1 U33895 ( .A(n25355), .B(reg_A[118]), .C(n25399), .D(reg_A[117]), .Y(
        n38981) );
  AOI22X1 U33896 ( .A(n25793), .B(reg_A[115]), .C(n25700), .D(reg_A[116]), .Y(
        n38980) );
  NAND2X1 U33897 ( .A(n38982), .B(n38983), .Y(n25408) );
  AOI22X1 U33898 ( .A(n25355), .B(reg_A[110]), .C(n25399), .D(reg_A[109]), .Y(
        n38983) );
  AOI22X1 U33899 ( .A(n25793), .B(reg_A[107]), .C(reg_A[108]), .D(n25700), .Y(
        n38982) );
  AOI22X1 U33900 ( .A(reg_B[123]), .B(n37135), .C(n25409), .D(n25406), .Y(
        n38978) );
  NAND2X1 U33901 ( .A(n38984), .B(n38985), .Y(n25406) );
  AOI22X1 U33902 ( .A(n25355), .B(reg_A[114]), .C(n25399), .D(reg_A[113]), .Y(
        n38985) );
  AOI22X1 U33903 ( .A(n25793), .B(reg_A[111]), .C(n25700), .D(reg_A[112]), .Y(
        n38984) );
  INVX1 U33904 ( .A(n25549), .Y(n25409) );
  OAI21X1 U33905 ( .A(n37653), .B(n36236), .C(n38986), .Y(n37135) );
  AOI22X1 U33906 ( .A(n36355), .B(n38002), .C(n36148), .D(n36241), .Y(n38986)
         );
  INVX1 U33907 ( .A(n36170), .Y(n36148) );
  NAND2X1 U33908 ( .A(n25793), .B(reg_A[127]), .Y(n36170) );
  INVX1 U33909 ( .A(n38506), .Y(n38002) );
  NOR2X1 U33910 ( .A(n38987), .B(n38988), .Y(n38506) );
  OAI22X1 U33911 ( .A(n25323), .B(n25568), .C(n25317), .D(n36136), .Y(n38988)
         );
  OAI21X1 U33912 ( .A(n25319), .B(n36246), .C(n36131), .Y(n38987) );
  NAND2X1 U33913 ( .A(n25793), .B(reg_A[123]), .Y(n36131) );
  AND2X1 U33914 ( .A(n38989), .B(n38990), .Y(n37653) );
  AOI22X1 U33915 ( .A(n25355), .B(reg_A[122]), .C(n25399), .D(reg_A[121]), .Y(
        n38990) );
  AOI22X1 U33916 ( .A(n25793), .B(reg_A[119]), .C(n25700), .D(reg_A[120]), .Y(
        n38989) );
  NOR2X1 U33917 ( .A(n25452), .B(n25656), .Y(n38976) );
  INVX1 U33918 ( .A(n38548), .Y(n38974) );
  NAND2X1 U33919 ( .A(n38991), .B(n38992), .Y(n38548) );
  AOI22X1 U33920 ( .A(reg_A[108]), .B(n25559), .C(reg_A[110]), .D(n25560), .Y(
        n38992) );
  AOI22X1 U33921 ( .A(reg_A[107]), .B(n25561), .C(reg_A[109]), .D(n25562), .Y(
        n38991) );
  NAND2X1 U33922 ( .A(n26003), .B(n38950), .Y(n27995) );
  NAND2X1 U33923 ( .A(n29998), .B(n37184), .Y(n38950) );
  INVX1 U33924 ( .A(n29082), .Y(n28055) );
  NOR2X1 U33925 ( .A(n34282), .B(n38993), .Y(n29082) );
  OAI21X1 U33926 ( .A(n25753), .B(n37184), .C(n38994), .Y(n38993) );
  OAI22X1 U33927 ( .A(n27676), .B(n37186), .C(n26002), .D(n26036), .Y(n38994)
         );
  AOI21X1 U33928 ( .A(n26596), .B(n25753), .C(n26864), .Y(n37186) );
  NAND2X1 U33929 ( .A(n26045), .B(n25029), .Y(n37184) );
  OAI21X1 U33930 ( .A(n25030), .B(n30951), .C(n28562), .Y(n34282) );
  NAND2X1 U33931 ( .A(n25613), .B(n25918), .Y(n28562) );
  INVX1 U33932 ( .A(n30990), .Y(n25918) );
  NAND2X1 U33933 ( .A(n26045), .B(n25604), .Y(n30990) );
  NAND2X1 U33934 ( .A(n26045), .B(n25044), .Y(n30951) );
  NAND3X1 U33935 ( .A(n38995), .B(n38996), .C(n38997), .Y(result[102]) );
  NOR2X1 U33936 ( .A(n38998), .B(n38999), .Y(n38997) );
  NAND2X1 U33937 ( .A(n39000), .B(n39001), .Y(n38999) );
  AOI21X1 U33938 ( .A(n26480), .B(n39002), .C(n39003), .Y(n39001) );
  OAI22X1 U33939 ( .A(n27190), .B(n38193), .C(n25525), .D(n39004), .Y(n39003)
         );
  INVX1 U33940 ( .A(n39005), .Y(n39004) );
  NAND2X1 U33941 ( .A(n39006), .B(n39007), .Y(n25525) );
  MUX2X1 U33942 ( .B(n25361), .A(n25448), .S(reg_B[103]), .Y(n39006) );
  NAND2X1 U33943 ( .A(n39008), .B(n39009), .Y(n38193) );
  AOI22X1 U33944 ( .A(n26601), .B(n25436), .C(n26602), .D(n25396), .Y(n39009)
         );
  AOI22X1 U33945 ( .A(n27012), .B(n25361), .C(n26597), .D(n25670), .Y(n39008)
         );
  OAI21X1 U33946 ( .A(n25545), .B(n25549), .C(n39010), .Y(n39002) );
  AOI22X1 U33947 ( .A(n25407), .B(n37681), .C(reg_B[123]), .D(n37298), .Y(
        n39010) );
  OAI21X1 U33948 ( .A(n38190), .B(n36236), .C(n39011), .Y(n37298) );
  AOI22X1 U33949 ( .A(n36355), .B(n36790), .C(n36241), .D(n36362), .Y(n39011)
         );
  INVX1 U33950 ( .A(n38596), .Y(n36362) );
  AOI21X1 U33951 ( .A(reg_A[127]), .B(n25700), .C(n36331), .Y(n38596) );
  NOR2X1 U33952 ( .A(n25397), .B(n25319), .Y(n36331) );
  INVX1 U33953 ( .A(n38595), .Y(n36790) );
  NOR2X1 U33954 ( .A(n39012), .B(n39013), .Y(n38595) );
  OAI22X1 U33955 ( .A(n25321), .B(n25568), .C(n25323), .D(n36136), .Y(n39013)
         );
  INVX1 U33956 ( .A(reg_A[124]), .Y(n25323) );
  OAI21X1 U33957 ( .A(n25317), .B(n36246), .C(n36743), .Y(n39012) );
  NAND2X1 U33958 ( .A(n25793), .B(reg_A[122]), .Y(n36743) );
  INVX1 U33959 ( .A(n37682), .Y(n38190) );
  NAND2X1 U33960 ( .A(n39014), .B(n39015), .Y(n37682) );
  AOI22X1 U33961 ( .A(n25355), .B(reg_A[121]), .C(n25399), .D(reg_A[120]), .Y(
        n39015) );
  AOI22X1 U33962 ( .A(n25793), .B(reg_A[118]), .C(n25700), .D(reg_A[119]), .Y(
        n39014) );
  NAND2X1 U33963 ( .A(n39016), .B(n39017), .Y(n37681) );
  AOI22X1 U33964 ( .A(n25355), .B(reg_A[117]), .C(n25399), .D(reg_A[116]), .Y(
        n39017) );
  AOI22X1 U33965 ( .A(n25793), .B(reg_A[114]), .C(n25700), .D(reg_A[115]), .Y(
        n39016) );
  INVX1 U33966 ( .A(n38108), .Y(n25545) );
  NAND2X1 U33967 ( .A(n39018), .B(n39019), .Y(n38108) );
  AOI22X1 U33968 ( .A(n25355), .B(reg_A[113]), .C(n25399), .D(reg_A[112]), .Y(
        n39019) );
  AOI22X1 U33969 ( .A(n25793), .B(reg_A[110]), .C(reg_A[111]), .D(n25700), .Y(
        n39018) );
  AOI21X1 U33970 ( .A(n37984), .B(n25552), .C(n39020), .Y(n39000) );
  OAI21X1 U33971 ( .A(n39021), .B(n25794), .C(n39022), .Y(n39020) );
  OAI21X1 U33972 ( .A(n39023), .B(n39024), .C(n25382), .Y(n39022) );
  OAI21X1 U33973 ( .A(n38095), .B(n25674), .C(n39025), .Y(n39024) );
  AOI22X1 U33974 ( .A(n25393), .B(n25547), .C(n25388), .D(n25535), .Y(n39025)
         );
  NAND2X1 U33975 ( .A(n39026), .B(n39027), .Y(n25535) );
  AOI22X1 U33976 ( .A(reg_A[107]), .B(n25559), .C(reg_A[109]), .D(n25560), .Y(
        n39027) );
  AOI22X1 U33977 ( .A(reg_A[106]), .B(n25561), .C(n25562), .D(reg_A[108]), .Y(
        n39026) );
  NAND2X1 U33978 ( .A(n39028), .B(n39029), .Y(n25547) );
  AOI22X1 U33979 ( .A(reg_A[105]), .B(n25355), .C(reg_A[104]), .D(n25399), .Y(
        n39029) );
  AOI22X1 U33980 ( .A(reg_A[102]), .B(n25793), .C(reg_A[103]), .D(n25700), .Y(
        n39028) );
  INVX1 U33981 ( .A(n25554), .Y(n38095) );
  OAI21X1 U33982 ( .A(n25452), .B(n25672), .C(n38145), .Y(n25554) );
  NAND2X1 U33983 ( .A(reg_A[110]), .B(n25561), .Y(n38145) );
  NAND2X1 U33984 ( .A(n39030), .B(n39031), .Y(n39023) );
  AOI22X1 U33985 ( .A(n39032), .B(reg_A[102]), .C(n25801), .D(reg_A[103]), .Y(
        n39031) );
  AOI22X1 U33986 ( .A(n25821), .B(reg_A[104]), .C(n25816), .D(reg_A[105]), .Y(
        n39030) );
  AOI21X1 U33987 ( .A(reg_B[110]), .B(n25692), .C(n39033), .Y(n39021) );
  OAI21X1 U33988 ( .A(n25436), .B(n39034), .C(n38752), .Y(n39033) );
  NAND2X1 U33989 ( .A(n38383), .B(n39035), .Y(n38752) );
  NAND2X1 U33990 ( .A(n38959), .B(n39036), .Y(n39034) );
  INVX1 U33991 ( .A(n25519), .Y(n39036) );
  NAND2X1 U33992 ( .A(n39037), .B(n39038), .Y(n25552) );
  AOI22X1 U33993 ( .A(n25355), .B(reg_A[109]), .C(n25399), .D(reg_A[108]), .Y(
        n39038) );
  AOI22X1 U33994 ( .A(reg_A[106]), .B(n25793), .C(reg_A[107]), .D(n25700), .Y(
        n39037) );
  NAND3X1 U33995 ( .A(n39039), .B(n39040), .C(n39041), .Y(n38998) );
  NOR2X1 U33996 ( .A(n39042), .B(n39043), .Y(n39041) );
  OAI21X1 U33997 ( .A(n25031), .B(n39044), .C(n39045), .Y(n39043) );
  OAI21X1 U33998 ( .A(n25352), .B(n25696), .C(n39046), .Y(n39045) );
  INVX1 U33999 ( .A(n39047), .Y(n39044) );
  MUX2X1 U34000 ( .B(n38963), .A(n39048), .S(reg_B[103]), .Y(n39047) );
  OAI21X1 U34001 ( .A(n25198), .B(n39049), .C(n39050), .Y(n39042) );
  NAND3X1 U34002 ( .A(n26267), .B(n39051), .C(n25562), .Y(n39050) );
  AOI22X1 U34003 ( .A(n25793), .B(n38820), .C(reg_B[127]), .D(n39052), .Y(
        n39049) );
  OAI22X1 U34004 ( .A(n25356), .B(n25361), .C(n25289), .D(n25544), .Y(n38820)
         );
  INVX1 U34005 ( .A(n26756), .Y(n25198) );
  NAND2X1 U34006 ( .A(n26610), .B(n25024), .Y(n26756) );
  OAI21X1 U34007 ( .A(n39053), .B(n29220), .C(reg_A[100]), .Y(n39040) );
  OAI21X1 U34008 ( .A(n25040), .B(n25835), .C(n39054), .Y(n29220) );
  NOR2X1 U34009 ( .A(n29394), .B(n27183), .Y(n39054) );
  INVX1 U34010 ( .A(n31351), .Y(n27183) );
  NAND2X1 U34011 ( .A(n26927), .B(n30910), .Y(n31351) );
  AOI22X1 U34012 ( .A(n25399), .B(n39055), .C(n25170), .D(n39056), .Y(n39039)
         );
  OAI22X1 U34013 ( .A(n39048), .B(n25802), .C(n39057), .D(n25373), .Y(n39056)
         );
  INVX1 U34014 ( .A(n38886), .Y(n39057) );
  NAND2X1 U34015 ( .A(n39058), .B(n38963), .Y(n38886) );
  AOI22X1 U34016 ( .A(n25574), .B(reg_A[102]), .C(reg_A[98]), .D(n38894), .Y(
        n38963) );
  AOI22X1 U34017 ( .A(n38895), .B(reg_A[96]), .C(reg_A[100]), .D(n25575), .Y(
        n39058) );
  OAI22X1 U34018 ( .A(n38892), .B(n26610), .C(n27438), .D(n39059), .Y(n39055)
         );
  NOR2X1 U34019 ( .A(n39060), .B(n39061), .Y(n38996) );
  OAI21X1 U34020 ( .A(n33194), .B(n25361), .C(n39062), .Y(n39061) );
  AOI22X1 U34021 ( .A(reg_A[101]), .B(n29291), .C(reg_A[99]), .D(n29155), .Y(
        n39062) );
  OAI21X1 U34022 ( .A(n25041), .B(n25835), .C(n39063), .Y(n29155) );
  NOR2X1 U34023 ( .A(n29439), .B(n27204), .Y(n39063) );
  INVX1 U34024 ( .A(n33975), .Y(n27204) );
  NAND2X1 U34025 ( .A(n26804), .B(n30910), .Y(n33975) );
  INVX1 U34026 ( .A(n30636), .Y(n29439) );
  OAI21X1 U34027 ( .A(n25042), .B(n25835), .C(n39064), .Y(n29291) );
  NOR2X1 U34028 ( .A(n29502), .B(n27188), .Y(n39064) );
  INVX1 U34029 ( .A(n33978), .Y(n27188) );
  NAND2X1 U34030 ( .A(n30910), .B(n26803), .Y(n33978) );
  INVX1 U34031 ( .A(n29366), .Y(n29502) );
  NOR2X1 U34032 ( .A(n29393), .B(n39065), .Y(n33194) );
  OAI21X1 U34033 ( .A(n25043), .B(n25835), .C(n34999), .Y(n39065) );
  NAND2X1 U34034 ( .A(n26924), .B(n30910), .Y(n34999) );
  INVX1 U34035 ( .A(n26864), .Y(n30910) );
  OAI21X1 U34036 ( .A(n38771), .B(n38577), .C(n39066), .Y(n39060) );
  AOI22X1 U34037 ( .A(n36280), .B(n25357), .C(n25310), .D(n39067), .Y(n39066)
         );
  NAND3X1 U34038 ( .A(n39068), .B(n39069), .C(n39070), .Y(n39067) );
  NOR2X1 U34039 ( .A(n39071), .B(n39072), .Y(n39070) );
  OR2X1 U34040 ( .A(n39073), .B(n39074), .Y(n39072) );
  OAI21X1 U34041 ( .A(n25043), .B(n25361), .C(n39075), .Y(n39074) );
  AOI22X1 U34042 ( .A(reg_A[114]), .B(n25635), .C(reg_A[115]), .D(n25325), .Y(
        n39075) );
  OAI21X1 U34043 ( .A(n25065), .B(n25332), .C(n39076), .Y(n39073) );
  AOI22X1 U34044 ( .A(reg_A[112]), .B(n25637), .C(reg_A[116]), .D(n25234), .Y(
        n39076) );
  INVX1 U34045 ( .A(reg_A[117]), .Y(n25332) );
  NAND3X1 U34046 ( .A(n39077), .B(n39078), .C(n39079), .Y(n39071) );
  AOI21X1 U34047 ( .A(reg_A[113]), .B(n25222), .C(n39080), .Y(n39079) );
  OAI22X1 U34048 ( .A(n25034), .B(n25450), .C(n25223), .D(n25452), .Y(n39080)
         );
  AOI22X1 U34049 ( .A(reg_A[108]), .B(n25253), .C(reg_A[109]), .D(n25628), .Y(
        n39078) );
  AOI22X1 U34050 ( .A(reg_A[106]), .B(n25075), .C(reg_A[107]), .D(n25123), .Y(
        n39077) );
  NOR2X1 U34051 ( .A(n39081), .B(n39082), .Y(n39069) );
  OAI21X1 U34052 ( .A(n25238), .B(n25494), .C(n39083), .Y(n39082) );
  AOI22X1 U34053 ( .A(reg_A[124]), .B(n25242), .C(reg_A[125]), .D(n25338), .Y(
        n39083) );
  NAND2X1 U34054 ( .A(n39084), .B(n39085), .Y(n39081) );
  AOI22X1 U34055 ( .A(reg_A[119]), .B(n25246), .C(reg_A[118]), .D(n25247), .Y(
        n39085) );
  AOI22X1 U34056 ( .A(reg_A[121]), .B(n25487), .C(reg_A[120]), .D(n25241), .Y(
        n39084) );
  NOR2X1 U34057 ( .A(n39086), .B(n39087), .Y(n39068) );
  OAI21X1 U34058 ( .A(n25040), .B(n25298), .C(n39088), .Y(n39087) );
  AOI22X1 U34059 ( .A(reg_A[103]), .B(n25135), .C(reg_A[105]), .D(n25136), .Y(
        n39088) );
  OAI21X1 U34060 ( .A(n25057), .B(n25319), .C(n39089), .Y(n39086) );
  AOI22X1 U34061 ( .A(reg_A[123]), .B(n25257), .C(reg_A[127]), .D(n25857), .Y(
        n39089) );
  INVX1 U34062 ( .A(n36439), .Y(n36280) );
  NAND2X1 U34063 ( .A(reg_B[125]), .B(reg_B[126]), .Y(n36439) );
  INVX1 U34064 ( .A(n38031), .Y(n38577) );
  NAND2X1 U34065 ( .A(n38004), .B(n38805), .Y(n38031) );
  INVX1 U34066 ( .A(n38461), .Y(n38805) );
  NOR2X1 U34067 ( .A(n25656), .B(n25697), .Y(n38461) );
  NAND2X1 U34068 ( .A(n25561), .B(n25604), .Y(n25656) );
  INVX1 U34069 ( .A(n38900), .Y(n38771) );
  OAI22X1 U34070 ( .A(n25289), .B(n38003), .C(n25820), .D(n25361), .Y(n38900)
         );
  NOR2X1 U34071 ( .A(n39090), .B(n39091), .Y(n38995) );
  NAND2X1 U34072 ( .A(n39092), .B(n39093), .Y(n39091) );
  AOI22X1 U34073 ( .A(n25730), .B(n39094), .C(n27402), .D(reg_A[103]), .Y(
        n39092) );
  NAND3X1 U34074 ( .A(n39095), .B(n39096), .C(n39097), .Y(n39094) );
  NOR2X1 U34075 ( .A(n39098), .B(n39099), .Y(n39097) );
  OAI22X1 U34076 ( .A(n26936), .B(n25474), .C(n25745), .D(n25469), .Y(n39099)
         );
  OAI21X1 U34077 ( .A(n25062), .B(n25298), .C(n39100), .Y(n39098) );
  AOI22X1 U34078 ( .A(reg_A[103]), .B(n26803), .C(reg_A[105]), .D(n26804), .Y(
        n39100) );
  AOI21X1 U34079 ( .A(reg_A[111]), .B(n25614), .C(n39101), .Y(n39096) );
  OAI22X1 U34080 ( .A(n26800), .B(n25470), .C(n26801), .D(n25468), .Y(n39101)
         );
  AOI22X1 U34081 ( .A(reg_A[110]), .B(n25615), .C(reg_A[102]), .D(n26924), .Y(
        n39095) );
  OAI21X1 U34082 ( .A(n29248), .B(n25287), .C(n39102), .Y(n39090) );
  AOI22X1 U34083 ( .A(reg_A[98]), .B(n29250), .C(reg_A[96]), .D(n29127), .Y(
        n39102) );
  OR2X1 U34084 ( .A(n27192), .B(n39103), .Y(n29127) );
  OAI21X1 U34085 ( .A(n26894), .B(n27523), .C(n39104), .Y(n39103) );
  OAI21X1 U34086 ( .A(n26530), .B(n25063), .C(n27676), .Y(n39104) );
  INVX1 U34087 ( .A(n25835), .Y(n27676) );
  INVX1 U34088 ( .A(n34598), .Y(n26894) );
  OAI21X1 U34089 ( .A(n25403), .B(n25131), .C(n27219), .Y(n34598) );
  INVX1 U34090 ( .A(n25211), .Y(n27219) );
  NAND2X1 U34091 ( .A(n30179), .B(n28311), .Y(n25211) );
  NAND2X1 U34092 ( .A(n26878), .B(n25604), .Y(n28311) );
  NAND2X1 U34093 ( .A(n26010), .B(n25029), .Y(n30179) );
  OAI21X1 U34094 ( .A(n39105), .B(n26864), .C(n28434), .Y(n27192) );
  NAND2X1 U34095 ( .A(n30427), .B(n26530), .Y(n28434) );
  NOR2X1 U34096 ( .A(n26530), .B(reg_B[1]), .Y(n39105) );
  INVX1 U34097 ( .A(n29129), .Y(n29250) );
  NOR2X1 U34098 ( .A(n31307), .B(n39106), .Y(n29129) );
  OAI21X1 U34099 ( .A(n26431), .B(n25835), .C(n29397), .Y(n39106) );
  INVX1 U34100 ( .A(n29507), .Y(n29397) );
  INVX1 U34101 ( .A(n27173), .Y(n31307) );
  NOR2X1 U34102 ( .A(n25721), .B(n25948), .Y(n27173) );
  INVX1 U34103 ( .A(n28122), .Y(n25948) );
  NAND2X1 U34104 ( .A(n30427), .B(n26003), .Y(n28122) );
  NOR2X1 U34105 ( .A(n26801), .B(n26864), .Y(n25721) );
  NOR2X1 U34106 ( .A(n27256), .B(n39107), .Y(n29248) );
  OAI21X1 U34107 ( .A(n25028), .B(n25835), .C(n30649), .Y(n39107) );
  NAND2X1 U34108 ( .A(n27358), .B(n25044), .Y(n25835) );
  OAI21X1 U34109 ( .A(n26864), .B(n26800), .C(n32117), .Y(n27256) );
  NAND2X1 U34110 ( .A(n30427), .B(n25751), .Y(n32117) );
  NAND3X1 U34111 ( .A(n39108), .B(n39109), .C(n39110), .Y(result[101]) );
  NOR2X1 U34112 ( .A(n39111), .B(n39112), .Y(n39110) );
  NAND3X1 U34113 ( .A(n39113), .B(n39093), .C(n39114), .Y(n39112) );
  NOR2X1 U34114 ( .A(n39115), .B(n39116), .Y(n39114) );
  OAI22X1 U34115 ( .A(n39117), .B(n37301), .C(n39048), .D(n25273), .Y(n39116)
         );
  INVX1 U34116 ( .A(n39118), .Y(n39048) );
  OAI21X1 U34117 ( .A(n25590), .B(n25670), .C(n39119), .Y(n39118) );
  AOI22X1 U34118 ( .A(n38894), .B(reg_A[97]), .C(reg_A[99]), .D(n25575), .Y(
        n39119) );
  OAI21X1 U34119 ( .A(n39120), .B(n27152), .C(n39121), .Y(n39115) );
  OAI21X1 U34120 ( .A(n39122), .B(n39123), .C(n27358), .Y(n39121) );
  OAI21X1 U34121 ( .A(n29339), .B(n25670), .C(n39124), .Y(n39123) );
  AOI22X1 U34122 ( .A(reg_A[97]), .B(n25650), .C(reg_A[100]), .D(n29341), .Y(
        n39124) );
  OAI21X1 U34123 ( .A(n25403), .B(n26431), .C(n25438), .Y(n25650) );
  NAND2X1 U34124 ( .A(n39125), .B(n39126), .Y(n39122) );
  AOI22X1 U34125 ( .A(n39127), .B(n29345), .C(reg_A[98]), .D(n29346), .Y(
        n39126) );
  NAND2X1 U34126 ( .A(n25599), .B(n36451), .Y(n29346) );
  INVX1 U34127 ( .A(n27374), .Y(n29345) );
  NAND2X1 U34128 ( .A(n25029), .B(n26030), .Y(n27374) );
  INVX1 U34129 ( .A(n38920), .Y(n39127) );
  NAND2X1 U34130 ( .A(n39128), .B(n39129), .Y(n38920) );
  AOI22X1 U34131 ( .A(n26292), .B(n25287), .C(n26293), .D(n25670), .Y(n39129)
         );
  NOR2X1 U34132 ( .A(reg_B[2]), .B(reg_B[4]), .Y(n26293) );
  NOR2X1 U34133 ( .A(n26452), .B(reg_B[4]), .Y(n26292) );
  AOI22X1 U34134 ( .A(n26294), .B(n25424), .C(n26295), .D(n25436), .Y(n39128)
         );
  NOR2X1 U34135 ( .A(n26863), .B(reg_B[2]), .Y(n26295) );
  AOI22X1 U34136 ( .A(reg_A[99]), .B(n29349), .C(reg_A[96]), .D(n29350), .Y(
        n39125) );
  NAND2X1 U34137 ( .A(n39130), .B(n39131), .Y(n29350) );
  OAI21X1 U34138 ( .A(n25063), .B(n38398), .C(n25044), .Y(n39131) );
  INVX1 U34139 ( .A(n37451), .Y(n39130) );
  NAND2X1 U34140 ( .A(n35069), .B(n27375), .Y(n37451) );
  NAND2X1 U34141 ( .A(n26530), .B(n25029), .Y(n27375) );
  OAI21X1 U34142 ( .A(reg_B[1]), .B(n38398), .C(n25604), .Y(n35069) );
  OR2X1 U34143 ( .A(n26530), .B(n26294), .Y(n38398) );
  NOR2X1 U34144 ( .A(n26452), .B(n26863), .Y(n26294) );
  NAND2X1 U34145 ( .A(n25598), .B(n38413), .Y(n29349) );
  AND2X1 U34146 ( .A(n39132), .B(n39133), .Y(n39120) );
  NOR2X1 U34147 ( .A(n39134), .B(n39135), .Y(n39133) );
  OAI21X1 U34148 ( .A(n26801), .B(n25296), .C(n39136), .Y(n39135) );
  AOI22X1 U34149 ( .A(reg_A[107]), .B(n26878), .C(reg_A[108]), .D(n25613), .Y(
        n39136) );
  OAI21X1 U34150 ( .A(n25062), .B(n25448), .C(n39137), .Y(n39134) );
  AOI22X1 U34151 ( .A(reg_A[102]), .B(n26803), .C(reg_A[104]), .D(n26804), .Y(
        n39137) );
  NOR2X1 U34152 ( .A(n39138), .B(n39139), .Y(n39132) );
  OAI22X1 U34153 ( .A(n25736), .B(n25670), .C(n31398), .D(n25452), .Y(n39139)
         );
  OAI21X1 U34154 ( .A(n27252), .B(n25474), .C(n39140), .Y(n39138) );
  AOI22X1 U34155 ( .A(reg_A[106]), .B(n25750), .C(reg_A[110]), .D(n25614), .Y(
        n39140) );
  AOI21X1 U34156 ( .A(n38895), .B(n39141), .C(n38812), .Y(n39093) );
  NOR2X1 U34157 ( .A(n38934), .B(n36338), .Y(n38812) );
  INVX1 U34158 ( .A(n36668), .Y(n36338) );
  NAND2X1 U34159 ( .A(n25551), .B(n36291), .Y(n36668) );
  NOR2X1 U34160 ( .A(n25424), .B(n25031), .Y(n39141) );
  NOR2X1 U34161 ( .A(n25343), .B(n39007), .Y(n38895) );
  AOI22X1 U34162 ( .A(n27402), .B(reg_A[102]), .C(n29361), .D(reg_A[103]), .Y(
        n39113) );
  INVX1 U34163 ( .A(n25717), .Y(n29361) );
  INVX1 U34164 ( .A(n25719), .Y(n27402) );
  NAND3X1 U34165 ( .A(n39142), .B(n39143), .C(n39144), .Y(n39111) );
  NOR2X1 U34166 ( .A(n39145), .B(n39146), .Y(n39144) );
  OAI21X1 U34167 ( .A(n25436), .B(n29366), .C(n39147), .Y(n39146) );
  OAI21X1 U34168 ( .A(n39148), .B(n39149), .C(n25382), .Y(n39147) );
  OAI21X1 U34169 ( .A(n39150), .B(n25674), .C(n39151), .Y(n39149) );
  AOI22X1 U34170 ( .A(n25393), .B(n25685), .C(n25388), .D(n25673), .Y(n39151)
         );
  NAND2X1 U34171 ( .A(n39152), .B(n39153), .Y(n25673) );
  AOI22X1 U34172 ( .A(reg_A[106]), .B(n25559), .C(n25560), .D(reg_A[108]), .Y(
        n39153) );
  AOI22X1 U34173 ( .A(reg_A[105]), .B(n25561), .C(n25562), .D(reg_A[107]), .Y(
        n39152) );
  NAND2X1 U34174 ( .A(n39154), .B(n39155), .Y(n25685) );
  AOI22X1 U34175 ( .A(reg_A[104]), .B(n25355), .C(n25399), .D(reg_A[103]), .Y(
        n39155) );
  AOI22X1 U34176 ( .A(reg_A[101]), .B(n25793), .C(reg_A[102]), .D(n25700), .Y(
        n39154) );
  INVX1 U34177 ( .A(n25689), .Y(n39150) );
  OAI21X1 U34178 ( .A(n25452), .B(n25668), .C(n39156), .Y(n25689) );
  AOI22X1 U34179 ( .A(reg_A[110]), .B(n25559), .C(reg_A[109]), .D(n25561), .Y(
        n39156) );
  NAND2X1 U34180 ( .A(n39157), .B(n39158), .Y(n39148) );
  AOI22X1 U34181 ( .A(n39032), .B(reg_A[101]), .C(n25801), .D(reg_A[102]), .Y(
        n39158) );
  AOI22X1 U34182 ( .A(n25821), .B(reg_A[103]), .C(n25816), .D(reg_A[104]), .Y(
        n39157) );
  OAI21X1 U34183 ( .A(n25424), .B(n30649), .C(n39159), .Y(n39145) );
  OAI21X1 U34184 ( .A(n39160), .B(n39161), .C(reg_A[98]), .Y(n39159) );
  OAI21X1 U34185 ( .A(n39162), .B(n39163), .C(n30636), .Y(n39161) );
  NAND2X1 U34186 ( .A(reg_B[103]), .B(n26504), .Y(n39163) );
  AND2X1 U34187 ( .A(n25427), .B(n37958), .Y(n39160) );
  NOR2X1 U34188 ( .A(n36246), .B(n25024), .Y(n37958) );
  NAND2X1 U34189 ( .A(n26045), .B(n34599), .Y(n30649) );
  OAI21X1 U34190 ( .A(n25403), .B(n26703), .C(n25207), .Y(n34599) );
  INVX1 U34191 ( .A(n28355), .Y(n25207) );
  NAND2X1 U34192 ( .A(n30355), .B(n25449), .Y(n28355) );
  NAND2X1 U34193 ( .A(n25750), .B(n25604), .Y(n25449) );
  NAND2X1 U34194 ( .A(n25751), .B(n25029), .Y(n30355) );
  OAI21X1 U34195 ( .A(n39164), .B(n39165), .C(n25310), .Y(n39143) );
  NAND3X1 U34196 ( .A(n39166), .B(n39167), .C(n39168), .Y(n39165) );
  NOR2X1 U34197 ( .A(n39169), .B(n39170), .Y(n39168) );
  OAI21X1 U34198 ( .A(n25043), .B(n25670), .C(n39171), .Y(n39170) );
  AOI22X1 U34199 ( .A(reg_A[113]), .B(n25635), .C(reg_A[114]), .D(n25325), .Y(
        n39171) );
  OAI21X1 U34200 ( .A(n25065), .B(n25337), .C(n39172), .Y(n39169) );
  AOI22X1 U34201 ( .A(reg_A[111]), .B(n25637), .C(reg_A[115]), .D(n25234), .Y(
        n39172) );
  NOR2X1 U34202 ( .A(n39173), .B(n39174), .Y(n39167) );
  OAI22X1 U34203 ( .A(n25028), .B(n25468), .C(n26431), .D(n25296), .Y(n39174)
         );
  INVX1 U34204 ( .A(reg_A[106]), .Y(n25468) );
  OAI22X1 U34205 ( .A(n25030), .B(n25469), .C(n25131), .D(n25470), .Y(n39173)
         );
  INVX1 U34206 ( .A(reg_A[107]), .Y(n25470) );
  AOI21X1 U34207 ( .A(reg_A[112]), .B(n25222), .C(n39175), .Y(n39166) );
  OAI22X1 U34208 ( .A(n25034), .B(n25474), .C(n25037), .D(n25450), .Y(n39175)
         );
  INVX1 U34209 ( .A(reg_A[110]), .Y(n25450) );
  NAND3X1 U34210 ( .A(n39176), .B(n39177), .C(n39178), .Y(n39164) );
  NOR2X1 U34211 ( .A(n39179), .B(n39180), .Y(n39178) );
  OAI21X1 U34212 ( .A(n25046), .B(n25490), .C(n39181), .Y(n39180) );
  AOI22X1 U34213 ( .A(reg_A[123]), .B(n25242), .C(reg_A[124]), .D(n25338), .Y(
        n39181) );
  NAND2X1 U34214 ( .A(n39182), .B(n39183), .Y(n39179) );
  AOI22X1 U34215 ( .A(reg_A[118]), .B(n25246), .C(reg_A[117]), .D(n25247), .Y(
        n39183) );
  AOI22X1 U34216 ( .A(reg_A[120]), .B(n25487), .C(reg_A[119]), .D(n25241), .Y(
        n39182) );
  NOR2X1 U34217 ( .A(n39184), .B(n39185), .Y(n39177) );
  OAI22X1 U34218 ( .A(n25059), .B(n25497), .C(n25320), .D(n25317), .Y(n39185)
         );
  INVX1 U34219 ( .A(reg_A[125]), .Y(n25317) );
  INVX1 U34220 ( .A(reg_A[127]), .Y(n25497) );
  OAI22X1 U34221 ( .A(n25322), .B(n25319), .C(n26719), .D(n25494), .Y(n39184)
         );
  AOI21X1 U34222 ( .A(reg_A[103]), .B(n25252), .C(n39186), .Y(n39176) );
  OAI22X1 U34223 ( .A(n25041), .B(n25298), .C(n25042), .D(n25361), .Y(n39186)
         );
  AOI22X1 U34224 ( .A(n37984), .B(n25687), .C(reg_A[101]), .D(n29393), .Y(
        n39142) );
  NAND2X1 U34225 ( .A(n39187), .B(n39188), .Y(n25687) );
  AOI22X1 U34226 ( .A(n25355), .B(reg_A[108]), .C(n25399), .D(reg_A[107]), .Y(
        n39188) );
  AOI22X1 U34227 ( .A(reg_A[105]), .B(n25793), .C(reg_A[106]), .D(n25700), .Y(
        n39187) );
  NOR2X1 U34228 ( .A(n39189), .B(n39190), .Y(n39109) );
  OAI21X1 U34229 ( .A(n39191), .B(n39192), .C(n39193), .Y(n39190) );
  AOI22X1 U34230 ( .A(n39005), .B(n25691), .C(n39194), .D(n25669), .Y(n39193)
         );
  INVX1 U34231 ( .A(n25348), .Y(n39194) );
  NAND2X1 U34232 ( .A(n25692), .B(n25188), .Y(n25348) );
  INVX1 U34233 ( .A(n38955), .Y(n25692) );
  INVX1 U34234 ( .A(n39195), .Y(n25691) );
  MUX2X1 U34235 ( .B(n39196), .A(n39197), .S(reg_B[103]), .Y(n39195) );
  NOR2X1 U34236 ( .A(reg_B[102]), .B(n25361), .Y(n39197) );
  INVX1 U34237 ( .A(n25350), .Y(n39192) );
  NAND3X1 U34238 ( .A(n39198), .B(n39199), .C(n39200), .Y(n39189) );
  AOI22X1 U34239 ( .A(n39201), .B(n38468), .C(n39202), .D(n38960), .Y(n39200)
         );
  MUX2X1 U34240 ( .B(n39203), .A(n39204), .S(reg_B[103]), .Y(n38960) );
  MUX2X1 U34241 ( .B(reg_A[100]), .A(reg_A[96]), .S(reg_B[101]), .Y(n39204) );
  MUX2X1 U34242 ( .B(reg_A[101]), .A(reg_A[97]), .S(reg_B[101]), .Y(n39203) );
  NOR2X1 U34243 ( .A(reg_B[102]), .B(n25031), .Y(n39202) );
  NOR2X1 U34244 ( .A(n25820), .B(n38387), .Y(n39201) );
  INVX1 U34245 ( .A(n25696), .Y(n38387) );
  NOR2X1 U34246 ( .A(n38958), .B(n25032), .Y(n25696) );
  OAI21X1 U34247 ( .A(n36329), .B(n25277), .C(n39052), .Y(n39199) );
  OAI22X1 U34248 ( .A(reg_B[126]), .B(n38902), .C(n25396), .D(n25425), .Y(
        n39052) );
  INVX1 U34249 ( .A(n38818), .Y(n38902) );
  OAI22X1 U34250 ( .A(n25356), .B(n25670), .C(n25287), .D(n25544), .Y(n38818)
         );
  INVX1 U34251 ( .A(n37303), .Y(n25277) );
  INVX1 U34252 ( .A(n36838), .Y(n36329) );
  NAND2X1 U34253 ( .A(n25932), .B(n36172), .Y(n36838) );
  OAI21X1 U34254 ( .A(n39053), .B(n29394), .C(reg_A[99]), .Y(n39198) );
  INVX1 U34255 ( .A(n29513), .Y(n29394) );
  INVX1 U34256 ( .A(n39205), .Y(n39053) );
  NAND3X1 U34257 ( .A(n26504), .B(n39206), .C(n25575), .Y(n39205) );
  NAND2X1 U34258 ( .A(n25029), .B(n25372), .Y(n25342) );
  NOR2X1 U34259 ( .A(n39207), .B(n39208), .Y(n39108) );
  OAI21X1 U34260 ( .A(n39209), .B(n39210), .C(n39211), .Y(n39208) );
  AOI22X1 U34261 ( .A(n38383), .B(n38798), .C(n26480), .D(n39212), .Y(n39211)
         );
  OAI21X1 U34262 ( .A(n38324), .B(n25549), .C(n39213), .Y(n39212) );
  AOI22X1 U34263 ( .A(n25407), .B(n37855), .C(reg_B[123]), .D(n37456), .Y(
        n39213) );
  OAI21X1 U34264 ( .A(n38395), .B(n36236), .C(n39214), .Y(n37456) );
  AOI22X1 U34265 ( .A(n36355), .B(n36877), .C(n36241), .D(n36911), .Y(n39214)
         );
  OAI21X1 U34266 ( .A(n25319), .B(n25568), .C(n39215), .Y(n36911) );
  AOI22X1 U34267 ( .A(n25399), .B(reg_A[127]), .C(n25793), .D(reg_A[125]), .Y(
        n39215) );
  NAND2X1 U34268 ( .A(n39216), .B(n39217), .Y(n36877) );
  AOI22X1 U34269 ( .A(n25355), .B(reg_A[124]), .C(n25399), .D(reg_A[123]), .Y(
        n39217) );
  AOI22X1 U34270 ( .A(n25793), .B(reg_A[121]), .C(n25700), .D(reg_A[122]), .Y(
        n39216) );
  INVX1 U34271 ( .A(n37856), .Y(n38395) );
  NAND2X1 U34272 ( .A(n39218), .B(n39219), .Y(n37856) );
  AOI22X1 U34273 ( .A(n25355), .B(reg_A[120]), .C(n25399), .D(reg_A[119]), .Y(
        n39219) );
  AOI22X1 U34274 ( .A(n25793), .B(reg_A[117]), .C(n25700), .D(reg_A[118]), .Y(
        n39218) );
  NAND2X1 U34275 ( .A(n39220), .B(n39221), .Y(n37855) );
  AOI22X1 U34276 ( .A(n25355), .B(reg_A[116]), .C(n25399), .D(reg_A[115]), .Y(
        n39221) );
  AOI22X1 U34277 ( .A(n25793), .B(reg_A[113]), .C(n25700), .D(reg_A[114]), .Y(
        n39220) );
  INVX1 U34278 ( .A(n25686), .Y(n38324) );
  NAND2X1 U34279 ( .A(n39222), .B(n39223), .Y(n25686) );
  AOI22X1 U34280 ( .A(n25355), .B(reg_A[112]), .C(n25399), .D(reg_A[111]), .Y(
        n39223) );
  AOI22X1 U34281 ( .A(n25793), .B(reg_A[109]), .C(reg_A[110]), .D(n25700), .Y(
        n39222) );
  INVX1 U34282 ( .A(n38004), .Y(n38798) );
  NAND2X1 U34283 ( .A(n25709), .B(n25188), .Y(n38004) );
  NOR2X1 U34284 ( .A(n39224), .B(reg_B[110]), .Y(n25709) );
  NOR2X1 U34285 ( .A(n38467), .B(n25424), .Y(n38383) );
  INVX1 U34286 ( .A(n39046), .Y(n39210) );
  OAI22X1 U34287 ( .A(n25519), .B(n25396), .C(reg_B[110]), .D(n38956), .Y(
        n39046) );
  INVX1 U34288 ( .A(n38817), .Y(n38956) );
  OAI22X1 U34289 ( .A(n25287), .B(n38003), .C(n25820), .D(n25670), .Y(n38817)
         );
  INVX1 U34290 ( .A(n25345), .Y(n39209) );
  NAND2X1 U34291 ( .A(n25513), .B(n38152), .Y(n25345) );
  NAND2X1 U34292 ( .A(n38959), .B(n25188), .Y(n38152) );
  INVX1 U34293 ( .A(n39224), .Y(n38959) );
  NAND2X1 U34294 ( .A(n39225), .B(n39226), .Y(n39207) );
  AOI22X1 U34295 ( .A(n38929), .B(n37920), .C(n29507), .D(reg_A[97]), .Y(
        n39226) );
  NOR2X1 U34296 ( .A(n25568), .B(n25024), .Y(n37920) );
  AOI22X1 U34297 ( .A(n25352), .B(n39227), .C(n36437), .D(n25357), .Y(n39225)
         );
  INVX1 U34298 ( .A(n38934), .Y(n25357) );
  NOR2X1 U34299 ( .A(n36177), .B(n25793), .Y(n36437) );
  INVX1 U34300 ( .A(n39228), .Y(n25352) );
  NAND3X1 U34301 ( .A(n39229), .B(n39230), .C(n39231), .Y(result[100]) );
  NOR2X1 U34302 ( .A(n39232), .B(n39233), .Y(n39231) );
  NAND3X1 U34303 ( .A(n39234), .B(n39235), .C(n39236), .Y(n39233) );
  AOI21X1 U34304 ( .A(reg_A[98]), .B(n31793), .C(n39237), .Y(n39236) );
  OAI21X1 U34305 ( .A(n33307), .B(n25396), .C(n39238), .Y(n39237) );
  OAI21X1 U34306 ( .A(n39239), .B(n39240), .C(n25730), .Y(n39238) );
  NAND2X1 U34307 ( .A(n39241), .B(n39242), .Y(n39240) );
  AOI22X1 U34308 ( .A(reg_A[109]), .B(n25614), .C(reg_A[108]), .D(n25615), .Y(
        n39242) );
  AOI22X1 U34309 ( .A(reg_A[111]), .B(n25616), .C(reg_A[110]), .D(n25607), .Y(
        n39241) );
  NAND2X1 U34310 ( .A(n39243), .B(n39244), .Y(n39239) );
  AOI22X1 U34311 ( .A(reg_A[106]), .B(n26878), .C(reg_A[107]), .D(n25613), .Y(
        n39244) );
  AOI22X1 U34312 ( .A(reg_A[104]), .B(n25749), .C(reg_A[105]), .D(n25750), .Y(
        n39243) );
  INVX1 U34313 ( .A(n31769), .Y(n33307) );
  OAI21X1 U34314 ( .A(n29467), .B(n31658), .C(n29366), .Y(n31769) );
  NAND2X1 U34315 ( .A(n26045), .B(n29568), .Y(n29366) );
  OAI21X1 U34316 ( .A(n25403), .B(n25784), .C(n27218), .Y(n29568) );
  INVX1 U34317 ( .A(n25441), .Y(n27218) );
  NAND2X1 U34318 ( .A(n28303), .B(n30791), .Y(n25441) );
  NAND2X1 U34319 ( .A(n26007), .B(n25029), .Y(n30791) );
  INVX1 U34320 ( .A(n29341), .Y(n29467) );
  OAI21X1 U34321 ( .A(n25403), .B(n25784), .C(n28303), .Y(n29341) );
  NAND2X1 U34322 ( .A(n26803), .B(n25604), .Y(n28303) );
  OAI21X1 U34323 ( .A(n25598), .B(n31658), .C(n29513), .Y(n31793) );
  NAND2X1 U34324 ( .A(n26045), .B(n29569), .Y(n29513) );
  OAI21X1 U34325 ( .A(n25403), .B(n25133), .C(n28353), .Y(n29569) );
  INVX1 U34326 ( .A(n27243), .Y(n28353) );
  NAND2X1 U34327 ( .A(n25437), .B(n38413), .Y(n27243) );
  NAND2X1 U34328 ( .A(n26009), .B(n25589), .Y(n38413) );
  INVX1 U34329 ( .A(n27637), .Y(n25598) );
  OAI21X1 U34330 ( .A(n25403), .B(n25133), .C(n25437), .Y(n27637) );
  NAND2X1 U34331 ( .A(n26927), .B(n25604), .Y(n25437) );
  OAI21X1 U34332 ( .A(n39245), .B(n39246), .C(n25382), .Y(n39235) );
  OAI21X1 U34333 ( .A(n39247), .B(n25674), .C(n39248), .Y(n39246) );
  AOI22X1 U34334 ( .A(n25393), .B(n25809), .C(n25388), .D(n25803), .Y(n39248)
         );
  NAND2X1 U34335 ( .A(n39249), .B(n39250), .Y(n25803) );
  AOI22X1 U34336 ( .A(reg_A[105]), .B(n25559), .C(reg_A[107]), .D(n25560), .Y(
        n39250) );
  AOI22X1 U34337 ( .A(reg_A[104]), .B(n25561), .C(reg_A[106]), .D(n25562), .Y(
        n39249) );
  INVX1 U34338 ( .A(n25558), .Y(n25388) );
  NAND2X1 U34339 ( .A(n38107), .B(n25604), .Y(n25558) );
  INVX1 U34340 ( .A(n38003), .Y(n38107) );
  NAND2X1 U34341 ( .A(n39251), .B(n39252), .Y(n25809) );
  AOI22X1 U34342 ( .A(n25355), .B(reg_A[103]), .C(reg_A[102]), .D(n25399), .Y(
        n39252) );
  AOI22X1 U34343 ( .A(reg_A[100]), .B(n25793), .C(reg_A[101]), .D(n25700), .Y(
        n39251) );
  INVX1 U34344 ( .A(n25569), .Y(n25393) );
  NAND2X1 U34345 ( .A(n38347), .B(n25604), .Y(n25674) );
  INVX1 U34346 ( .A(n38032), .Y(n38347) );
  NAND2X1 U34347 ( .A(reg_B[108]), .B(n38159), .Y(n38032) );
  INVX1 U34348 ( .A(n25825), .Y(n39247) );
  NAND2X1 U34349 ( .A(n39253), .B(n39254), .Y(n25825) );
  AOI22X1 U34350 ( .A(reg_A[109]), .B(n25559), .C(n25560), .D(reg_A[111]), .Y(
        n39254) );
  INVX1 U34351 ( .A(n25671), .Y(n25560) );
  INVX1 U34352 ( .A(n25672), .Y(n25559) );
  AOI22X1 U34353 ( .A(reg_A[108]), .B(n25561), .C(n25562), .D(reg_A[110]), .Y(
        n39253) );
  INVX1 U34354 ( .A(n25668), .Y(n25562) );
  INVX1 U34355 ( .A(n25669), .Y(n25561) );
  NAND2X1 U34356 ( .A(n39255), .B(n39256), .Y(n39245) );
  AOI22X1 U34357 ( .A(n39032), .B(reg_A[100]), .C(n25801), .D(reg_A[101]), .Y(
        n39256) );
  NOR2X1 U34358 ( .A(n25672), .B(n38971), .Y(n25801) );
  NAND2X1 U34359 ( .A(reg_B[111]), .B(n25521), .Y(n25672) );
  NOR2X1 U34360 ( .A(n25669), .B(n38971), .Y(n39032) );
  NAND2X1 U34361 ( .A(n25521), .B(n37993), .Y(n25669) );
  AOI22X1 U34362 ( .A(n25821), .B(reg_A[102]), .C(n25816), .D(reg_A[103]), .Y(
        n39255) );
  NOR2X1 U34363 ( .A(n25671), .B(n38971), .Y(n25816) );
  NAND2X1 U34364 ( .A(reg_B[110]), .B(reg_B[111]), .Y(n25671) );
  NOR2X1 U34365 ( .A(n25668), .B(n38971), .Y(n25821) );
  NAND2X1 U34366 ( .A(reg_B[110]), .B(n37993), .Y(n25668) );
  AOI22X1 U34367 ( .A(n26480), .B(n39257), .C(n25053), .D(n39258), .Y(n39234)
         );
  NAND3X1 U34368 ( .A(n39259), .B(n39260), .C(n39261), .Y(n39258) );
  INVX1 U34369 ( .A(n39262), .Y(n39261) );
  OAI21X1 U34370 ( .A(n37229), .B(n25374), .C(n39263), .Y(n39262) );
  AOI22X1 U34371 ( .A(n25376), .B(n25379), .C(reg_A[96]), .D(n25690), .Y(
        n39263) );
  NOR2X1 U34372 ( .A(n25343), .B(n26999), .Y(n25690) );
  INVX1 U34373 ( .A(n25802), .Y(n25379) );
  NAND2X1 U34374 ( .A(reg_B[103]), .B(n25589), .Y(n25802) );
  NAND2X1 U34375 ( .A(reg_B[127]), .B(n25044), .Y(n37229) );
  AOI22X1 U34376 ( .A(n39264), .B(n38468), .C(n25604), .D(n39265), .Y(n39260)
         );
  OAI21X1 U34377 ( .A(n39266), .B(n38958), .C(n38955), .Y(n39265) );
  NAND3X1 U34378 ( .A(n39035), .B(n25820), .C(reg_A[96]), .Y(n38955) );
  NAND2X1 U34379 ( .A(reg_B[111]), .B(n39035), .Y(n38958) );
  MUX2X1 U34380 ( .B(n25436), .A(n25289), .S(reg_B[110]), .Y(n38468) );
  NOR2X1 U34381 ( .A(n39224), .B(n38971), .Y(n39264) );
  NAND2X1 U34382 ( .A(n25522), .B(n25604), .Y(n38971) );
  NAND2X1 U34383 ( .A(n39035), .B(n37993), .Y(n39224) );
  INVX1 U34384 ( .A(n25591), .Y(n39035) );
  NAND3X1 U34385 ( .A(n39267), .B(n39268), .C(n39269), .Y(n25591) );
  NOR2X1 U34386 ( .A(n39270), .B(n39271), .Y(n39269) );
  NAND2X1 U34387 ( .A(n39272), .B(n25574), .Y(n39271) );
  NOR2X1 U34388 ( .A(reg_B[100]), .B(n26377), .Y(n39272) );
  NAND2X1 U34389 ( .A(n25984), .B(n26275), .Y(n26377) );
  INVX1 U34390 ( .A(n26067), .Y(n26275) );
  NAND2X1 U34391 ( .A(n26063), .B(n26197), .Y(n26067) );
  INVX1 U34392 ( .A(reg_B[93]), .Y(n26197) );
  INVX1 U34393 ( .A(reg_B[92]), .Y(n26063) );
  NAND2X1 U34394 ( .A(n25950), .B(n25976), .Y(n25972) );
  INVX1 U34395 ( .A(reg_B[95]), .Y(n25976) );
  INVX1 U34396 ( .A(reg_B[94]), .Y(n25950) );
  NAND2X1 U34397 ( .A(n39273), .B(n39206), .Y(n39270) );
  NOR2X1 U34398 ( .A(reg_B[105]), .B(reg_B[104]), .Y(n39273) );
  NOR2X1 U34399 ( .A(reg_B[97]), .B(n39274), .Y(n39268) );
  OR2X1 U34400 ( .A(reg_B[99]), .B(reg_B[98]), .Y(n39274) );
  NOR2X1 U34401 ( .A(reg_B[106]), .B(n39275), .Y(n39267) );
  OR2X1 U34402 ( .A(reg_B[96]), .B(reg_B[107]), .Y(n39275) );
  AOI22X1 U34403 ( .A(reg_A[100]), .B(n39276), .C(reg_A[98]), .D(n39277), .Y(
        n39259) );
  OAI21X1 U34404 ( .A(n25569), .B(n36136), .C(n38897), .Y(n39277) );
  NAND2X1 U34405 ( .A(n38889), .B(n25575), .Y(n38897) );
  OAI21X1 U34406 ( .A(n25569), .B(n25397), .C(n25711), .Y(n39276) );
  NAND2X1 U34407 ( .A(n38889), .B(n25574), .Y(n25711) );
  INVX1 U34408 ( .A(n25590), .Y(n25574) );
  INVX1 U34409 ( .A(n25373), .Y(n38889) );
  NAND2X1 U34410 ( .A(n25029), .B(n39206), .Y(n25373) );
  NAND2X1 U34411 ( .A(n25427), .B(n25044), .Y(n25569) );
  OAI21X1 U34412 ( .A(n25808), .B(n25549), .C(n39278), .Y(n39257) );
  AOI22X1 U34413 ( .A(n25407), .B(n37882), .C(reg_B[123]), .D(n37474), .Y(
        n39278) );
  OAI21X1 U34414 ( .A(n38416), .B(n36236), .C(n39279), .Y(n37474) );
  AOI22X1 U34415 ( .A(n36355), .B(n37883), .C(n36241), .D(n36619), .Y(n39279)
         );
  NAND2X1 U34416 ( .A(n39280), .B(n39281), .Y(n36619) );
  AOI22X1 U34417 ( .A(n25355), .B(reg_A[127]), .C(n25399), .D(reg_A[126]), .Y(
        n39281) );
  AOI22X1 U34418 ( .A(n25793), .B(reg_A[124]), .C(n25700), .D(reg_A[125]), .Y(
        n39280) );
  INVX1 U34419 ( .A(n36288), .Y(n36241) );
  NAND2X1 U34420 ( .A(reg_B[124]), .B(n36177), .Y(n36288) );
  NAND2X1 U34421 ( .A(n39282), .B(n39283), .Y(n37883) );
  AOI22X1 U34422 ( .A(n25355), .B(reg_A[123]), .C(n25399), .D(reg_A[122]), .Y(
        n39283) );
  AOI22X1 U34423 ( .A(n25793), .B(reg_A[120]), .C(n25700), .D(reg_A[121]), .Y(
        n39282) );
  INVX1 U34424 ( .A(n37884), .Y(n38416) );
  NAND2X1 U34425 ( .A(n39284), .B(n39285), .Y(n37884) );
  AOI22X1 U34426 ( .A(n25355), .B(reg_A[119]), .C(n25399), .D(reg_A[118]), .Y(
        n39285) );
  AOI22X1 U34427 ( .A(n25793), .B(reg_A[116]), .C(n25700), .D(reg_A[117]), .Y(
        n39284) );
  NAND2X1 U34428 ( .A(n39286), .B(n39287), .Y(n37882) );
  AOI22X1 U34429 ( .A(n25355), .B(reg_A[115]), .C(n25399), .D(reg_A[114]), .Y(
        n39287) );
  AOI22X1 U34430 ( .A(n25793), .B(reg_A[112]), .C(n25700), .D(reg_A[113]), .Y(
        n39286) );
  INVX1 U34431 ( .A(n25546), .Y(n25407) );
  NAND2X1 U34432 ( .A(n36686), .B(reg_B[125]), .Y(n25546) );
  NAND2X1 U34433 ( .A(n36686), .B(n36177), .Y(n25549) );
  INVX1 U34434 ( .A(n36318), .Y(n36686) );
  NAND2X1 U34435 ( .A(reg_B[124]), .B(n25551), .Y(n36318) );
  INVX1 U34436 ( .A(n38822), .Y(n25808) );
  NAND2X1 U34437 ( .A(n39288), .B(n39289), .Y(n38822) );
  AOI22X1 U34438 ( .A(n25355), .B(reg_A[111]), .C(n25399), .D(reg_A[110]), .Y(
        n39289) );
  AOI22X1 U34439 ( .A(n25793), .B(reg_A[108]), .C(reg_A[109]), .D(n25700), .Y(
        n39288) );
  OR2X1 U34440 ( .A(n39290), .B(n39291), .Y(n39232) );
  OAI21X1 U34441 ( .A(n39266), .B(n39228), .C(n39292), .Y(n39291) );
  AOI22X1 U34442 ( .A(n25350), .B(n25376), .C(n38785), .D(n29209), .Y(n39292)
         );
  INVX1 U34443 ( .A(n27190), .Y(n29209) );
  NAND2X1 U34444 ( .A(n30427), .B(n26452), .Y(n27190) );
  INVX1 U34445 ( .A(n38411), .Y(n38785) );
  NAND2X1 U34446 ( .A(n39293), .B(n39294), .Y(n38411) );
  AOI22X1 U34447 ( .A(n26601), .B(n25289), .C(n26602), .D(n25287), .Y(n39294)
         );
  AOI22X1 U34448 ( .A(n27012), .B(n25436), .C(n26597), .D(n25396), .Y(n39293)
         );
  NAND2X1 U34449 ( .A(reg_B[4]), .B(n26030), .Y(n27454) );
  NAND2X1 U34450 ( .A(n26030), .B(n26863), .Y(n26599) );
  OAI22X1 U34451 ( .A(n25590), .B(n25396), .C(n39162), .D(n25287), .Y(n25376)
         );
  NOR2X1 U34452 ( .A(n39206), .B(n26151), .Y(n25350) );
  NAND2X1 U34453 ( .A(reg_B[111]), .B(n26267), .Y(n39228) );
  INVX1 U34454 ( .A(n25346), .Y(n39266) );
  OAI21X1 U34455 ( .A(n25519), .B(n25287), .C(n39295), .Y(n25346) );
  NAND3X1 U34456 ( .A(n25522), .B(n25521), .C(reg_A[99]), .Y(n39295) );
  INVX1 U34457 ( .A(reg_B[110]), .Y(n25521) );
  OAI21X1 U34458 ( .A(n39296), .B(n25513), .C(n39297), .Y(n39290) );
  AOI22X1 U34459 ( .A(reg_A[100]), .B(n39298), .C(n39005), .D(n25826), .Y(
        n39297) );
  INVX1 U34460 ( .A(n39299), .Y(n25826) );
  MUX2X1 U34461 ( .B(n39300), .A(n39196), .S(reg_B[103]), .Y(n39299) );
  MUX2X1 U34462 ( .B(n25448), .A(n25670), .S(n39007), .Y(n39196) );
  MUX2X1 U34463 ( .B(n25436), .A(n25361), .S(reg_B[102]), .Y(n39300) );
  NOR2X1 U34464 ( .A(n25523), .B(reg_B[101]), .Y(n39005) );
  NAND2X1 U34465 ( .A(n25382), .B(n25589), .Y(n25523) );
  OAI21X1 U34466 ( .A(n29339), .B(n31658), .C(n29532), .Y(n39298) );
  NOR2X1 U34467 ( .A(n29393), .B(n36973), .Y(n29532) );
  INVX1 U34468 ( .A(n33195), .Y(n36973) );
  NAND2X1 U34469 ( .A(n25730), .B(n26924), .Y(n33195) );
  NAND2X1 U34470 ( .A(n33358), .B(n25795), .Y(n29393) );
  NAND2X1 U34471 ( .A(n26928), .B(n26004), .Y(n25795) );
  INVX1 U34472 ( .A(n29466), .Y(n29339) );
  OAI21X1 U34473 ( .A(n25403), .B(n25228), .C(n27442), .Y(n29466) );
  NAND2X1 U34474 ( .A(n26267), .B(n37993), .Y(n25513) );
  INVX1 U34475 ( .A(reg_B[111]), .Y(n37993) );
  NAND2X1 U34476 ( .A(n25170), .B(n25604), .Y(n26147) );
  INVX1 U34477 ( .A(n39227), .Y(n39296) );
  OAI22X1 U34478 ( .A(n25289), .B(n25519), .C(reg_B[110]), .D(n38898), .Y(
        n39227) );
  INVX1 U34479 ( .A(n39051), .Y(n38898) );
  OAI22X1 U34480 ( .A(n25424), .B(n38003), .C(n25820), .D(n25436), .Y(n39051)
         );
  NAND2X1 U34481 ( .A(reg_B[109]), .B(n38467), .Y(n38003) );
  NAND2X1 U34482 ( .A(reg_B[110]), .B(n25522), .Y(n25519) );
  INVX1 U34483 ( .A(n25820), .Y(n25522) );
  NAND2X1 U34484 ( .A(n38467), .B(n38159), .Y(n25820) );
  INVX1 U34485 ( .A(reg_B[109]), .Y(n38159) );
  INVX1 U34486 ( .A(reg_B[108]), .Y(n38467) );
  NOR2X1 U34487 ( .A(n39301), .B(n39302), .Y(n39230) );
  OAI21X1 U34488 ( .A(n31797), .B(n25424), .C(n39303), .Y(n39302) );
  AOI22X1 U34489 ( .A(n25310), .B(n39304), .C(reg_A[103]), .D(n26739), .Y(
        n39303) );
  OAI21X1 U34490 ( .A(n25747), .B(n27152), .C(n25718), .Y(n26739) );
  INVX1 U34491 ( .A(n29547), .Y(n25718) );
  NOR2X1 U34492 ( .A(n25726), .B(n30090), .Y(n29547) );
  NAND3X1 U34493 ( .A(n39305), .B(n39306), .C(n39307), .Y(n39304) );
  NOR2X1 U34494 ( .A(n39308), .B(n39309), .Y(n39307) );
  NAND3X1 U34495 ( .A(n39310), .B(n39311), .C(n39312), .Y(n39309) );
  AOI21X1 U34496 ( .A(reg_A[103]), .B(n25136), .C(n39313), .Y(n39312) );
  OAI22X1 U34497 ( .A(n25042), .B(n25670), .C(n25319), .D(n25316), .Y(n39313)
         );
  INVX1 U34498 ( .A(reg_A[126]), .Y(n25319) );
  INVX1 U34499 ( .A(reg_A[101]), .Y(n25670) );
  AOI22X1 U34500 ( .A(reg_A[121]), .B(n25257), .C(reg_A[125]), .D(n25857), .Y(
        n39311) );
  INVX1 U34501 ( .A(n25322), .Y(n25857) );
  AOI22X1 U34502 ( .A(n25647), .B(reg_A[124]), .C(reg_A[127]), .D(n25648), .Y(
        n39310) );
  INVX1 U34503 ( .A(n25318), .Y(n25648) );
  NAND3X1 U34504 ( .A(n39314), .B(n39315), .C(n39316), .Y(n39308) );
  AOI21X1 U34505 ( .A(reg_A[120]), .B(n25339), .C(n39317), .Y(n39316) );
  OAI22X1 U34506 ( .A(n25491), .B(n25321), .C(n25492), .D(n25494), .Y(n39317)
         );
  INVX1 U34507 ( .A(reg_A[122]), .Y(n25494) );
  INVX1 U34508 ( .A(reg_A[123]), .Y(n25321) );
  AOI22X1 U34509 ( .A(reg_A[117]), .B(n25246), .C(reg_A[116]), .D(n25247), .Y(
        n39315) );
  AOI22X1 U34510 ( .A(reg_A[119]), .B(n25487), .C(reg_A[118]), .D(n25241), .Y(
        n39314) );
  NOR2X1 U34511 ( .A(n39318), .B(n39319), .Y(n39306) );
  OAI21X1 U34512 ( .A(n25034), .B(n25469), .C(n39320), .Y(n39319) );
  AOI22X1 U34513 ( .A(reg_A[105]), .B(n25123), .C(reg_A[109]), .D(n25629), .Y(
        n39320) );
  INVX1 U34514 ( .A(reg_A[108]), .Y(n25469) );
  NAND2X1 U34515 ( .A(n39321), .B(n39322), .Y(n39318) );
  AOI22X1 U34516 ( .A(reg_A[102]), .B(n25252), .C(reg_A[106]), .D(n25253), .Y(
        n39322) );
  AOI22X1 U34517 ( .A(reg_A[107]), .B(n25628), .C(reg_A[104]), .D(n25066), .Y(
        n39321) );
  NOR2X1 U34518 ( .A(n39323), .B(n39324), .Y(n39305) );
  OAI21X1 U34519 ( .A(n25043), .B(n25436), .C(n39325), .Y(n39324) );
  AOI22X1 U34520 ( .A(reg_A[112]), .B(n25635), .C(reg_A[113]), .D(n25325), .Y(
        n39325) );
  NAND2X1 U34521 ( .A(n39326), .B(n39327), .Y(n39323) );
  AOI22X1 U34522 ( .A(reg_A[111]), .B(n25222), .C(reg_A[110]), .D(n25637), .Y(
        n39327) );
  AOI22X1 U34523 ( .A(reg_A[114]), .B(n25234), .C(reg_A[115]), .D(n25235), .Y(
        n39326) );
  INVX1 U34524 ( .A(reg_A[96]), .Y(n25424) );
  INVX1 U34525 ( .A(n39328), .Y(n31797) );
  OAI21X1 U34526 ( .A(n29473), .B(n31658), .C(n39329), .Y(n39328) );
  AOI21X1 U34527 ( .A(n30427), .B(reg_B[2]), .C(n29507), .Y(n39329) );
  NOR2X1 U34528 ( .A(n27523), .B(n26895), .Y(n29507) );
  AOI21X1 U34529 ( .A(n25044), .B(n25075), .C(n27242), .Y(n26895) );
  NAND2X1 U34530 ( .A(n25438), .B(n31058), .Y(n27242) );
  NAND2X1 U34531 ( .A(n26003), .B(n25589), .Y(n31058) );
  NAND2X1 U34532 ( .A(n25749), .B(n25604), .Y(n25438) );
  INVX1 U34533 ( .A(n29998), .Y(n30427) );
  NAND2X1 U34534 ( .A(n27358), .B(n25589), .Y(n29998) );
  AND2X1 U34535 ( .A(n34070), .B(n39330), .Y(n29473) );
  OAI21X1 U34536 ( .A(n25044), .B(n25604), .C(reg_B[2]), .Y(n39330) );
  INVX1 U34537 ( .A(n32943), .Y(n34070) );
  OAI21X1 U34538 ( .A(n26664), .B(n25403), .C(n35476), .Y(n32943) );
  NAND2X1 U34539 ( .A(reg_B[1]), .B(n25604), .Y(n35476) );
  INVX1 U34540 ( .A(n26036), .Y(n26664) );
  NAND2X1 U34541 ( .A(n27677), .B(n26596), .Y(n26036) );
  OAI21X1 U34542 ( .A(n25427), .B(n38934), .C(n39331), .Y(n39301) );
  AOI22X1 U34543 ( .A(reg_A[97]), .B(n31770), .C(n37984), .D(n38807), .Y(
        n39331) );
  NAND2X1 U34544 ( .A(n39332), .B(n39333), .Y(n38807) );
  AOI22X1 U34545 ( .A(n25355), .B(reg_A[107]), .C(reg_A[106]), .D(n25399), .Y(
        n39333) );
  NAND2X1 U34546 ( .A(reg_B[126]), .B(n36172), .Y(n36136) );
  NAND2X1 U34547 ( .A(reg_B[127]), .B(reg_B[126]), .Y(n36246) );
  AOI22X1 U34548 ( .A(reg_A[104]), .B(n25793), .C(reg_A[105]), .D(n25700), .Y(
        n39332) );
  NAND2X1 U34549 ( .A(reg_B[127]), .B(n25428), .Y(n25568) );
  NAND2X1 U34550 ( .A(n25428), .B(n36172), .Y(n25397) );
  INVX1 U34551 ( .A(n36960), .Y(n37984) );
  NAND2X1 U34552 ( .A(n26480), .B(n25405), .Y(n36960) );
  NAND2X1 U34553 ( .A(n25382), .B(n25044), .Y(n26996) );
  OAI21X1 U34554 ( .A(n25599), .B(n31658), .C(n30636), .Y(n31770) );
  NAND2X1 U34555 ( .A(n26045), .B(n36883), .Y(n30636) );
  OAI21X1 U34556 ( .A(n25403), .B(n25254), .C(n39334), .Y(n36883) );
  INVX1 U34557 ( .A(n27241), .Y(n39334) );
  NAND2X1 U34558 ( .A(n30437), .B(n36451), .Y(n27241) );
  NAND2X1 U34559 ( .A(n26008), .B(n25029), .Y(n36451) );
  INVX1 U34560 ( .A(n27358), .Y(n31658) );
  INVX1 U34561 ( .A(n27740), .Y(n25599) );
  OAI21X1 U34562 ( .A(n25403), .B(n25254), .C(n30437), .Y(n27740) );
  NAND2X1 U34563 ( .A(n26804), .B(n25604), .Y(n30437) );
  NAND2X1 U34564 ( .A(reg_A[96]), .B(n25932), .Y(n38934) );
  NAND2X1 U34565 ( .A(n25372), .B(n25044), .Y(n27438) );
  NOR2X1 U34566 ( .A(n39335), .B(n39336), .Y(n39229) );
  OAI22X1 U34567 ( .A(n25374), .B(n37301), .C(n39191), .D(n25273), .Y(n39336)
         );
  NAND2X1 U34568 ( .A(n26186), .B(n39206), .Y(n25273) );
  INVX1 U34569 ( .A(reg_B[103]), .Y(n39206) );
  NAND2X1 U34570 ( .A(n25170), .B(n25589), .Y(n26151) );
  INVX1 U34571 ( .A(n39337), .Y(n39191) );
  OAI21X1 U34572 ( .A(n25590), .B(n25436), .C(n39338), .Y(n39337) );
  AOI22X1 U34573 ( .A(n38894), .B(reg_A[96]), .C(reg_A[98]), .D(n25575), .Y(
        n39338) );
  INVX1 U34574 ( .A(n39162), .Y(n25575) );
  NAND2X1 U34575 ( .A(reg_B[102]), .B(n25343), .Y(n39162) );
  INVX1 U34576 ( .A(n25413), .Y(n38894) );
  NAND2X1 U34577 ( .A(reg_B[101]), .B(n39007), .Y(n25413) );
  NAND2X1 U34578 ( .A(n25343), .B(n39007), .Y(n25590) );
  INVX1 U34579 ( .A(reg_B[102]), .Y(n39007) );
  INVX1 U34580 ( .A(reg_B[101]), .Y(n25343) );
  NAND2X1 U34581 ( .A(reg_B[127]), .B(n25699), .Y(n37301) );
  INVX1 U34582 ( .A(n25278), .Y(n25374) );
  OAI21X1 U34583 ( .A(n25287), .B(n25425), .C(n39339), .Y(n25278) );
  NAND3X1 U34584 ( .A(n25427), .B(n25428), .C(reg_A[99]), .Y(n39339) );
  INVX1 U34585 ( .A(reg_B[126]), .Y(n25428) );
  OAI21X1 U34586 ( .A(n39117), .B(n37303), .C(n39340), .Y(n39335) );
  AOI22X1 U34587 ( .A(reg_A[102]), .B(n26783), .C(reg_A[101]), .D(n28923), .Y(
        n39340) );
  OAI21X1 U34588 ( .A(n25748), .B(n27152), .C(n25719), .Y(n28923) );
  NAND2X1 U34589 ( .A(n26928), .B(n26007), .Y(n25719) );
  OAI21X1 U34590 ( .A(n25062), .B(n27152), .C(n25717), .Y(n26783) );
  NAND2X1 U34591 ( .A(n26928), .B(n26009), .Y(n25717) );
  NAND2X1 U34592 ( .A(n25699), .B(n36172), .Y(n37303) );
  INVX1 U34593 ( .A(reg_B[127]), .Y(n36172) );
  INVX1 U34594 ( .A(n26610), .Y(n25699) );
  INVX1 U34595 ( .A(n39341), .Y(n39117) );
  OAI22X1 U34596 ( .A(reg_B[126]), .B(n38892), .C(n25289), .D(n25425), .Y(
        n39341) );
  NAND2X1 U34597 ( .A(n25427), .B(reg_B[126]), .Y(n25425) );
  AOI21X1 U34598 ( .A(reg_A[96]), .B(n25405), .C(n38929), .Y(n38892) );
  INVX1 U34599 ( .A(n39059), .Y(n38929) );
  NAND2X1 U34600 ( .A(reg_A[100]), .B(n25427), .Y(n39059) );
  INVX1 U34601 ( .A(n25356), .Y(n25427) );
  NAND2X1 U34602 ( .A(n36356), .B(n25551), .Y(n25356) );
  INVX1 U34603 ( .A(n36236), .Y(n36356) );
  NAND2X1 U34604 ( .A(n36291), .B(n36177), .Y(n36236) );
  INVX1 U34605 ( .A(reg_B[125]), .Y(n36177) );
  INVX1 U34606 ( .A(n25544), .Y(n25405) );
  NAND2X1 U34607 ( .A(n36355), .B(n25551), .Y(n25544) );
  INVX1 U34608 ( .A(reg_B[123]), .Y(n25551) );
  INVX1 U34609 ( .A(n36247), .Y(n36355) );
  NAND2X1 U34610 ( .A(reg_B[125]), .B(n36291), .Y(n36247) );
  INVX1 U34611 ( .A(reg_B[124]), .Y(n36291) );
  NAND2X1 U34612 ( .A(n39342), .B(n39343), .Y(result[0]) );
  AOI21X1 U34613 ( .A(n25310), .B(n39344), .C(n39345), .Y(n39343) );
  NAND2X1 U34614 ( .A(n39346), .B(n39347), .Y(n39345) );
  OAI21X1 U34615 ( .A(n39348), .B(n39349), .C(n25730), .Y(n39347) );
  INVX1 U34616 ( .A(n27152), .Y(n25730) );
  NAND2X1 U34617 ( .A(n25203), .B(n25604), .Y(n27152) );
  NAND3X1 U34618 ( .A(n39350), .B(n39351), .C(n39352), .Y(n39349) );
  NOR2X1 U34619 ( .A(n39353), .B(n39354), .Y(n39352) );
  OAI22X1 U34620 ( .A(n26742), .B(n25736), .C(n25206), .D(n25737), .Y(n39354)
         );
  OAI22X1 U34621 ( .A(n25255), .B(n25738), .C(n29279), .D(n25739), .Y(n39353)
         );
  AOI22X1 U34622 ( .A(n25615), .B(reg_A[8]), .C(n25616), .D(reg_A[11]), .Y(
        n39351) );
  AOI22X1 U34623 ( .A(n25607), .B(reg_A[10]), .C(n25608), .D(reg_A[14]), .Y(
        n39350) );
  NAND3X1 U34624 ( .A(n39355), .B(n39356), .C(n39357), .Y(n39348) );
  NOR2X1 U34625 ( .A(n39358), .B(n39359), .Y(n39357) );
  OAI22X1 U34626 ( .A(n26677), .B(n25745), .C(n25128), .D(n25746), .Y(n39359)
         );
  OAI22X1 U34627 ( .A(n25130), .B(n25747), .C(n25748), .D(n25177), .Y(n39358)
         );
  AOI22X1 U34628 ( .A(n25613), .B(reg_A[7]), .C(n25749), .D(reg_A[4]), .Y(
        n39356) );
  AOI22X1 U34629 ( .A(n25750), .B(reg_A[5]), .C(n25614), .D(reg_A[9]), .Y(
        n39355) );
  OAI21X1 U34630 ( .A(n39360), .B(n39361), .C(reg_A[0]), .Y(n39346) );
  OAI21X1 U34631 ( .A(n33394), .B(n33724), .C(n35222), .Y(n39361) );
  AOI21X1 U34632 ( .A(n28040), .B(n25170), .C(n39362), .Y(n35222) );
  OAI21X1 U34633 ( .A(n33911), .B(n26610), .C(n33358), .Y(n39362) );
  NAND2X1 U34634 ( .A(n26045), .B(n25284), .Y(n33358) );
  OAI21X1 U34635 ( .A(n25403), .B(n25043), .C(n25204), .Y(n25284) );
  NOR2X1 U34636 ( .A(n27389), .B(n30792), .Y(n25204) );
  NOR2X1 U34637 ( .A(n26943), .B(n26999), .Y(n30792) );
  INVX1 U34638 ( .A(n25589), .Y(n26999) );
  INVX1 U34639 ( .A(n27442), .Y(n27389) );
  NAND2X1 U34640 ( .A(n26924), .B(n25604), .Y(n27442) );
  NAND3X1 U34641 ( .A(n39363), .B(alu_op[2]), .C(alu_op[4]), .Y(n27523) );
  NAND2X1 U34642 ( .A(n25170), .B(n25044), .Y(n26610) );
  NAND3X1 U34643 ( .A(alu_op[2]), .B(n39364), .C(n39363), .Y(n25697) );
  INVX1 U34644 ( .A(n34088), .Y(n28040) );
  NOR2X1 U34645 ( .A(n25372), .B(n27358), .Y(n33724) );
  NOR2X1 U34646 ( .A(n25589), .B(n25044), .Y(n33394) );
  NAND2X1 U34647 ( .A(n26864), .B(n25032), .Y(n39360) );
  NAND2X1 U34648 ( .A(n25604), .B(n25372), .Y(n25794) );
  NOR2X1 U34649 ( .A(n39365), .B(alu_op[4]), .Y(n25372) );
  NAND2X1 U34650 ( .A(n27358), .B(n25604), .Y(n26864) );
  NOR2X1 U34651 ( .A(n39364), .B(n39365), .Y(n27358) );
  NAND3X1 U34652 ( .A(alu_op[3]), .B(alu_op[2]), .C(n39366), .Y(n39365) );
  NOR2X1 U34653 ( .A(alu_op[1]), .B(n39367), .Y(n39366) );
  NAND2X1 U34654 ( .A(n39368), .B(n39369), .Y(n39344) );
  NOR2X1 U34655 ( .A(n39370), .B(n39371), .Y(n39369) );
  NAND3X1 U34656 ( .A(n39372), .B(n39373), .C(n39374), .Y(n39371) );
  NOR2X1 U34657 ( .A(n39375), .B(n39376), .Y(n39374) );
  OAI22X1 U34658 ( .A(n27961), .B(n25316), .C(n32918), .D(n25318), .Y(n39376)
         );
  NAND2X1 U34659 ( .A(n25616), .B(reg_B[0]), .Y(n25318) );
  INVX1 U34660 ( .A(reg_A[27]), .Y(n32918) );
  NAND2X1 U34661 ( .A(n25607), .B(reg_B[0]), .Y(n25316) );
  INVX1 U34662 ( .A(reg_A[26]), .Y(n27961) );
  OAI22X1 U34663 ( .A(n27962), .B(n25320), .C(n27960), .D(n25322), .Y(n39375)
         );
  NAND2X1 U34664 ( .A(n25614), .B(reg_B[0]), .Y(n25322) );
  INVX1 U34665 ( .A(reg_A[25]), .Y(n27960) );
  NAND2X1 U34666 ( .A(n25615), .B(reg_B[0]), .Y(n25320) );
  INVX1 U34667 ( .A(reg_A[24]), .Y(n27962) );
  AOI22X1 U34668 ( .A(n25631), .B(reg_A[30]), .C(n25764), .D(reg_A[31]), .Y(
        n39373) );
  INVX1 U34669 ( .A(n25852), .Y(n25764) );
  NAND2X1 U34670 ( .A(n37982), .B(reg_B[0]), .Y(n25852) );
  INVX1 U34671 ( .A(n25854), .Y(n25631) );
  NAND2X1 U34672 ( .A(n25608), .B(reg_B[0]), .Y(n25854) );
  AOI22X1 U34673 ( .A(n25324), .B(reg_A[28]), .C(n25765), .D(reg_A[29]), .Y(
        n39372) );
  INVX1 U34674 ( .A(n25498), .Y(n25765) );
  NAND2X1 U34675 ( .A(n25610), .B(reg_B[0]), .Y(n25498) );
  INVX1 U34676 ( .A(n25499), .Y(n25324) );
  NAND2X1 U34677 ( .A(n25609), .B(reg_B[0]), .Y(n25499) );
  NAND3X1 U34678 ( .A(n39377), .B(n39378), .C(n39379), .Y(n39370) );
  NOR2X1 U34679 ( .A(n39380), .B(n39381), .Y(n39379) );
  OAI22X1 U34680 ( .A(n25051), .B(n25224), .C(n25243), .D(n25220), .Y(n39381)
         );
  NAND2X1 U34681 ( .A(n26804), .B(reg_B[0]), .Y(n25243) );
  NAND2X1 U34682 ( .A(n26927), .B(reg_B[0]), .Y(n25331) );
  OAI22X1 U34683 ( .A(n25334), .B(n25250), .C(n25336), .D(n27953), .Y(n39380)
         );
  NAND2X1 U34684 ( .A(reg_B[0]), .B(n26803), .Y(n25336) );
  NAND2X1 U34685 ( .A(n26924), .B(reg_B[0]), .Y(n25334) );
  AOI22X1 U34686 ( .A(reg_A[22]), .B(n25242), .C(n25338), .D(reg_A[23]), .Y(
        n39378) );
  NAND2X1 U34687 ( .A(n25613), .B(reg_B[0]), .Y(n25491) );
  NAND2X1 U34688 ( .A(reg_B[0]), .B(n26878), .Y(n25492) );
  AOI22X1 U34689 ( .A(reg_A[20]), .B(n25339), .C(reg_A[21]), .D(n25257), .Y(
        n39377) );
  NAND2X1 U34690 ( .A(n25750), .B(reg_B[0]), .Y(n26719) );
  NAND2X1 U34691 ( .A(n25749), .B(reg_B[0]), .Y(n25238) );
  NOR2X1 U34692 ( .A(n39382), .B(n39383), .Y(n39368) );
  NAND3X1 U34693 ( .A(n39384), .B(n39385), .C(n39386), .Y(n39383) );
  NOR2X1 U34694 ( .A(n39387), .B(n39388), .Y(n39386) );
  OAI22X1 U34695 ( .A(n26742), .B(n25228), .C(n25206), .D(n25229), .Y(n39388)
         );
  NAND2X1 U34696 ( .A(n25610), .B(n27677), .Y(n25229) );
  INVX1 U34697 ( .A(n25737), .Y(n25610) );
  NAND2X1 U34698 ( .A(reg_B[1]), .B(n25751), .Y(n25737) );
  NAND2X1 U34699 ( .A(n26924), .B(n27677), .Y(n25228) );
  INVX1 U34700 ( .A(n25736), .Y(n26924) );
  NAND2X1 U34701 ( .A(n26004), .B(n26596), .Y(n25736) );
  OAI22X1 U34702 ( .A(n25255), .B(n25231), .C(n29279), .D(n25482), .Y(n39387)
         );
  NAND2X1 U34703 ( .A(n37982), .B(n27677), .Y(n25482) );
  INVX1 U34704 ( .A(n25739), .Y(n37982) );
  NAND2X1 U34705 ( .A(reg_B[1]), .B(n26002), .Y(n25739) );
  NAND2X1 U34706 ( .A(n25609), .B(n27677), .Y(n25231) );
  INVX1 U34707 ( .A(n25738), .Y(n25609) );
  NAND2X1 U34708 ( .A(reg_B[1]), .B(n26003), .Y(n25738) );
  INVX1 U34709 ( .A(reg_A[12]), .Y(n25255) );
  AOI22X1 U34710 ( .A(n25124), .B(reg_A[8]), .C(n25222), .D(reg_A[11]), .Y(
        n39385) );
  NAND2X1 U34711 ( .A(n25616), .B(n27677), .Y(n25473) );
  NAND2X1 U34712 ( .A(reg_B[1]), .B(n26008), .Y(n29558) );
  NAND2X1 U34713 ( .A(n25615), .B(n27677), .Y(n25467) );
  NAND2X1 U34714 ( .A(reg_B[1]), .B(n26004), .Y(n27252) );
  INVX1 U34715 ( .A(n26943), .Y(n26004) );
  AOI22X1 U34716 ( .A(n25637), .B(reg_A[10]), .C(n25234), .D(reg_A[14]), .Y(
        n39384) );
  NAND2X1 U34717 ( .A(n25608), .B(n27677), .Y(n25475) );
  NAND2X1 U34718 ( .A(reg_B[1]), .B(n26010), .Y(n32194) );
  NAND2X1 U34719 ( .A(n25607), .B(n27677), .Y(n25219) );
  NAND2X1 U34720 ( .A(reg_B[1]), .B(n26009), .Y(n31398) );
  NAND3X1 U34721 ( .A(n39389), .B(n39390), .C(n39391), .Y(n39382) );
  NOR2X1 U34722 ( .A(n39392), .B(n39393), .Y(n39391) );
  OAI22X1 U34723 ( .A(n26677), .B(n25131), .C(n25128), .D(n25133), .Y(n39393)
         );
  NAND2X1 U34724 ( .A(n26927), .B(n27677), .Y(n25133) );
  INVX1 U34725 ( .A(n25746), .Y(n26927) );
  NAND2X1 U34726 ( .A(n26009), .B(n26596), .Y(n25746) );
  NAND2X1 U34727 ( .A(n26878), .B(n27677), .Y(n25131) );
  NAND2X1 U34728 ( .A(n26010), .B(n26596), .Y(n25745) );
  OAI22X1 U34729 ( .A(n25130), .B(n25254), .C(n25177), .D(n25784), .Y(n39392)
         );
  NAND2X1 U34730 ( .A(n26803), .B(n27677), .Y(n25784) );
  NAND2X1 U34731 ( .A(n26007), .B(n26596), .Y(n25748) );
  NAND2X1 U34732 ( .A(n26804), .B(n27677), .Y(n25254) );
  NAND2X1 U34733 ( .A(n26008), .B(n26596), .Y(n25747) );
  AOI22X1 U34734 ( .A(n25628), .B(reg_A[7]), .C(n25070), .D(reg_A[4]), .Y(
        n39390) );
  INVX1 U34735 ( .A(n26431), .Y(n25122) );
  NAND2X1 U34736 ( .A(n25749), .B(n27677), .Y(n26431) );
  NAND2X1 U34737 ( .A(n26003), .B(n26596), .Y(n26801) );
  INVX1 U34738 ( .A(n26945), .Y(n26003) );
  NAND2X1 U34739 ( .A(n25613), .B(n27677), .Y(n25129) );
  NAND2X1 U34740 ( .A(n26002), .B(n26596), .Y(n26936) );
  INVX1 U34741 ( .A(n25753), .Y(n26002) );
  AOI22X1 U34742 ( .A(n25123), .B(reg_A[5]), .C(n25629), .D(reg_A[9]), .Y(
        n39389) );
  NAND2X1 U34743 ( .A(n25614), .B(n27677), .Y(n25223) );
  NAND2X1 U34744 ( .A(reg_B[1]), .B(n26007), .Y(n27253) );
  NAND2X1 U34745 ( .A(n25750), .B(n27677), .Y(n26703) );
  INVX1 U34746 ( .A(reg_B[0]), .Y(n27677) );
  NAND2X1 U34747 ( .A(n25751), .B(n26596), .Y(n26800) );
  INVX1 U34748 ( .A(reg_B[1]), .Y(n26596) );
  INVX1 U34749 ( .A(n26944), .Y(n25751) );
  NAND2X1 U34750 ( .A(n25203), .B(n25044), .Y(n26990) );
  AOI22X1 U34751 ( .A(n25382), .B(n39394), .C(n26928), .D(n39395), .Y(n39342)
         );
  NAND3X1 U34752 ( .A(n39396), .B(n39397), .C(n39398), .Y(n39395) );
  NOR2X1 U34753 ( .A(n39399), .B(n39400), .Y(n39398) );
  OAI22X1 U34754 ( .A(n26742), .B(n26943), .C(n29265), .D(n26944), .Y(n39400)
         );
  NAND2X1 U34755 ( .A(n25025), .B(reg_B[4]), .Y(n26944) );
  INVX1 U34756 ( .A(reg_A[5]), .Y(n29265) );
  NAND2X1 U34757 ( .A(n26032), .B(n26863), .Y(n26943) );
  OAI22X1 U34758 ( .A(n30569), .B(n26945), .C(n25132), .D(n25753), .Y(n39399)
         );
  NAND2X1 U34759 ( .A(n26530), .B(reg_B[4]), .Y(n25753) );
  NAND2X1 U34760 ( .A(n25025), .B(n26863), .Y(n26945) );
  NOR2X1 U34761 ( .A(n26452), .B(reg_B[3]), .Y(n26034) );
  INVX1 U34762 ( .A(reg_A[4]), .Y(n30569) );
  AOI22X1 U34763 ( .A(reg_A[1]), .B(n26007), .C(n26008), .D(reg_A[3]), .Y(
        n39397) );
  INVX1 U34764 ( .A(n30090), .Y(n26008) );
  NAND2X1 U34765 ( .A(n26602), .B(n26452), .Y(n30090) );
  NAND2X1 U34766 ( .A(reg_B[3]), .B(reg_B[4]), .Y(n27455) );
  INVX1 U34767 ( .A(n27925), .Y(n26007) );
  NAND2X1 U34768 ( .A(reg_B[4]), .B(n26032), .Y(n27925) );
  NAND2X1 U34769 ( .A(n26452), .B(n26030), .Y(n35474) );
  INVX1 U34770 ( .A(reg_B[3]), .Y(n26030) );
  AOI22X1 U34771 ( .A(n26009), .B(reg_A[2]), .C(n26010), .D(reg_A[6]), .Y(
        n39396) );
  INVX1 U34772 ( .A(n25754), .Y(n26010) );
  NAND2X1 U34773 ( .A(n26530), .B(n26863), .Y(n25754) );
  NAND2X1 U34774 ( .A(reg_B[2]), .B(reg_B[3]), .Y(n26208) );
  INVX1 U34775 ( .A(n31144), .Y(n26009) );
  NAND2X1 U34776 ( .A(n26601), .B(n26452), .Y(n31144) );
  INVX1 U34777 ( .A(reg_B[2]), .Y(n26452) );
  NAND2X1 U34778 ( .A(reg_B[3]), .B(n26863), .Y(n27575) );
  INVX1 U34779 ( .A(reg_B[4]), .Y(n26863) );
  INVX1 U34780 ( .A(n25726), .Y(n26928) );
  NAND2X1 U34781 ( .A(n25203), .B(n25029), .Y(n25726) );
  NAND3X1 U34782 ( .A(n39363), .B(n39401), .C(alu_op[4]), .Y(n30931) );
  NAND3X1 U34783 ( .A(n39402), .B(n39403), .C(n39404), .Y(n39394) );
  NOR2X1 U34784 ( .A(n39405), .B(n39406), .Y(n39404) );
  OAI21X1 U34785 ( .A(n34088), .B(n26742), .C(n39407), .Y(n39406) );
  OAI21X1 U34786 ( .A(n39408), .B(n39409), .C(n25044), .Y(n39407) );
  NOR2X1 U34787 ( .A(n39410), .B(ctrl_ww[1]), .Y(n25097) );
  OAI21X1 U34788 ( .A(n26742), .B(n33911), .C(n39411), .Y(n39409) );
  AOI22X1 U34789 ( .A(reg_B[27]), .B(n35612), .C(n30644), .D(n31783), .Y(
        n39411) );
  NAND2X1 U34790 ( .A(n39412), .B(n39413), .Y(n31783) );
  AOI22X1 U34791 ( .A(n25156), .B(reg_A[8]), .C(n25142), .D(reg_A[9]), .Y(
        n39413) );
  AOI22X1 U34792 ( .A(reg_A[10]), .B(n25258), .C(reg_A[11]), .D(n26761), .Y(
        n39412) );
  INVX1 U34793 ( .A(n25099), .Y(n30644) );
  NAND2X1 U34794 ( .A(n33919), .B(n33955), .Y(n25099) );
  NAND2X1 U34795 ( .A(n39414), .B(n39415), .Y(n35612) );
  AOI22X1 U34796 ( .A(n34188), .B(n26777), .C(n34180), .D(n26778), .Y(n39415)
         );
  NAND2X1 U34797 ( .A(n39416), .B(n39417), .Y(n26778) );
  AOI22X1 U34798 ( .A(reg_A[24]), .B(n25156), .C(n25142), .D(reg_A[25]), .Y(
        n39417) );
  AOI22X1 U34799 ( .A(reg_A[26]), .B(n25258), .C(reg_A[27]), .D(n26761), .Y(
        n39416) );
  INVX1 U34800 ( .A(n33957), .Y(n34180) );
  NAND2X1 U34801 ( .A(reg_B[28]), .B(n33955), .Y(n33957) );
  NAND2X1 U34802 ( .A(n39418), .B(n39419), .Y(n26777) );
  AOI22X1 U34803 ( .A(reg_A[28]), .B(n25156), .C(n25142), .D(reg_A[29]), .Y(
        n39419) );
  AOI22X1 U34804 ( .A(reg_A[30]), .B(n25258), .C(reg_A[31]), .D(n26761), .Y(
        n39418) );
  NOR2X1 U34805 ( .A(n34493), .B(n33955), .Y(n34188) );
  AOI22X1 U34806 ( .A(n34189), .B(n36037), .C(n34190), .D(n26773), .Y(n39414)
         );
  NAND2X1 U34807 ( .A(n39420), .B(n39421), .Y(n26773) );
  AOI22X1 U34808 ( .A(reg_A[20]), .B(n25156), .C(n25142), .D(reg_A[21]), .Y(
        n39421) );
  AOI22X1 U34809 ( .A(reg_A[22]), .B(n25258), .C(reg_A[23]), .D(n26761), .Y(
        n39420) );
  INVX1 U34810 ( .A(n34009), .Y(n34190) );
  NAND2X1 U34811 ( .A(reg_B[29]), .B(n34493), .Y(n34009) );
  NAND2X1 U34812 ( .A(n39422), .B(n39423), .Y(n36037) );
  AOI22X1 U34813 ( .A(reg_A[16]), .B(n25156), .C(n25142), .D(reg_A[17]), .Y(
        n39423) );
  AOI22X1 U34814 ( .A(reg_A[18]), .B(n25258), .C(reg_A[19]), .D(n26761), .Y(
        n39422) );
  INVX1 U34815 ( .A(n34230), .Y(n34189) );
  NAND2X1 U34816 ( .A(n34493), .B(n33955), .Y(n34230) );
  NAND2X1 U34817 ( .A(n33890), .B(n32933), .Y(n33911) );
  INVX1 U34818 ( .A(n33915), .Y(n33890) );
  NAND2X1 U34819 ( .A(n32934), .B(n33865), .Y(n33915) );
  NAND2X1 U34820 ( .A(n39424), .B(n39425), .Y(n39408) );
  AOI22X1 U34821 ( .A(n25110), .B(n39426), .C(reg_A[1]), .D(n32984), .Y(n39425) );
  INVX1 U34822 ( .A(n32950), .Y(n32984) );
  NAND2X1 U34823 ( .A(n32933), .B(n34405), .Y(n32950) );
  INVX1 U34824 ( .A(n33977), .Y(n34405) );
  NAND2X1 U34825 ( .A(reg_B[31]), .B(n32934), .Y(n33977) );
  NAND2X1 U34826 ( .A(n33955), .B(n34176), .Y(n34012) );
  OAI22X1 U34827 ( .A(n25130), .B(n25264), .C(n25128), .D(n29305), .Y(n39426)
         );
  INVX1 U34828 ( .A(n26775), .Y(n25110) );
  NAND2X1 U34829 ( .A(n32933), .B(n33955), .Y(n26775) );
  INVX1 U34830 ( .A(reg_B[29]), .Y(n33955) );
  AOI22X1 U34831 ( .A(n25101), .B(n31831), .C(n26772), .D(n26771), .Y(n39424)
         );
  NAND2X1 U34832 ( .A(n39427), .B(n39428), .Y(n26771) );
  AOI22X1 U34833 ( .A(reg_A[12]), .B(n25156), .C(n25142), .D(reg_A[13]), .Y(
        n39428) );
  AOI22X1 U34834 ( .A(reg_A[14]), .B(n25258), .C(reg_A[15]), .D(n26761), .Y(
        n39427) );
  INVX1 U34835 ( .A(n25106), .Y(n26772) );
  NAND2X1 U34836 ( .A(n33919), .B(reg_B[29]), .Y(n25106) );
  INVX1 U34837 ( .A(n34465), .Y(n33919) );
  NAND2X1 U34838 ( .A(reg_B[28]), .B(n31782), .Y(n34465) );
  NAND2X1 U34839 ( .A(n39429), .B(n39430), .Y(n31831) );
  AOI22X1 U34840 ( .A(n25156), .B(reg_A[4]), .C(n25142), .D(reg_A[5]), .Y(
        n39430) );
  NAND2X1 U34841 ( .A(reg_B[31]), .B(n34176), .Y(n26758) );
  NAND2X1 U34842 ( .A(n34176), .B(n33865), .Y(n25262) );
  INVX1 U34843 ( .A(reg_B[30]), .Y(n34176) );
  AOI22X1 U34844 ( .A(n25258), .B(reg_A[6]), .C(n26761), .D(reg_A[7]), .Y(
        n39429) );
  NAND2X1 U34845 ( .A(reg_B[30]), .B(reg_B[31]), .Y(n25264) );
  NAND2X1 U34846 ( .A(reg_B[30]), .B(n33865), .Y(n29305) );
  INVX1 U34847 ( .A(reg_B[31]), .Y(n33865) );
  INVX1 U34848 ( .A(n28033), .Y(n25101) );
  NAND2X1 U34849 ( .A(n32933), .B(reg_B[29]), .Y(n28033) );
  INVX1 U34850 ( .A(n33807), .Y(n32933) );
  NAND2X1 U34851 ( .A(n31782), .B(n34493), .Y(n33807) );
  INVX1 U34852 ( .A(reg_B[28]), .Y(n34493) );
  INVX1 U34853 ( .A(reg_B[27]), .Y(n31782) );
  INVX1 U34854 ( .A(reg_A[0]), .Y(n26742) );
  NOR2X1 U34855 ( .A(n31809), .B(n27980), .Y(n34088) );
  NOR2X1 U34856 ( .A(n31786), .B(n29235), .Y(n27980) );
  NOR2X1 U34857 ( .A(n30631), .B(n26692), .Y(n31809) );
  OAI22X1 U34858 ( .A(n34076), .B(n25130), .C(n32947), .D(n25177), .Y(n39405)
         );
  AOI22X1 U34859 ( .A(n25172), .B(n28023), .C(n27984), .D(n28009), .Y(n32947)
         );
  INVX1 U34860 ( .A(n33000), .Y(n34076) );
  OAI21X1 U34861 ( .A(n25194), .B(n30631), .C(n39431), .Y(n33000) );
  NAND3X1 U34862 ( .A(reg_B[7]), .B(reg_B[6]), .C(n27984), .Y(n39431) );
  AOI21X1 U34863 ( .A(n32997), .B(n31803), .C(n39432), .Y(n39403) );
  OAI22X1 U34864 ( .A(n35295), .B(n25128), .C(n26780), .D(n28026), .Y(n39432)
         );
  NAND2X1 U34865 ( .A(n35865), .B(n25604), .Y(n28026) );
  INVX1 U34866 ( .A(n35728), .Y(n35865) );
  NAND2X1 U34867 ( .A(reg_B[12]), .B(n26723), .Y(n35728) );
  INVX1 U34868 ( .A(n31802), .Y(n26780) );
  NAND2X1 U34869 ( .A(n39433), .B(n39434), .Y(n31802) );
  AOI22X1 U34870 ( .A(reg_A[10]), .B(n26733), .C(reg_A[9]), .D(n25172), .Y(
        n39434) );
  AOI22X1 U34871 ( .A(reg_A[11]), .B(n26734), .C(n25116), .D(reg_A[8]), .Y(
        n39433) );
  AOI22X1 U34872 ( .A(n26733), .B(n28023), .C(n27984), .D(n27985), .Y(n35295)
         );
  INVX1 U34873 ( .A(n29235), .Y(n27984) );
  NAND2X1 U34874 ( .A(n25029), .B(n31789), .Y(n29235) );
  INVX1 U34875 ( .A(reg_B[5]), .Y(n31789) );
  INVX1 U34876 ( .A(n30631), .Y(n28023) );
  NAND2X1 U34877 ( .A(n25604), .B(n31796), .Y(n30631) );
  NOR2X1 U34878 ( .A(reg_B[12]), .B(reg_B[13]), .Y(n31796) );
  NAND2X1 U34879 ( .A(n39435), .B(n39436), .Y(n31803) );
  AOI22X1 U34880 ( .A(n39437), .B(reg_B[7]), .C(n28009), .D(reg_A[5]), .Y(
        n39436) );
  NOR2X1 U34881 ( .A(n28041), .B(reg_B[6]), .Y(n28009) );
  NOR2X1 U34882 ( .A(n25132), .B(n28005), .Y(n39437) );
  AOI22X1 U34883 ( .A(n27985), .B(reg_A[6]), .C(n27986), .D(reg_A[4]), .Y(
        n39435) );
  INVX1 U34884 ( .A(n31786), .Y(n27986) );
  NAND2X1 U34885 ( .A(n28005), .B(n28041), .Y(n31786) );
  INVX1 U34886 ( .A(reg_B[7]), .Y(n28041) );
  NOR2X1 U34887 ( .A(n28005), .B(reg_B[7]), .Y(n27985) );
  INVX1 U34888 ( .A(reg_B[6]), .Y(n28005) );
  INVX1 U34889 ( .A(n27982), .Y(n32997) );
  NAND2X1 U34890 ( .A(reg_B[5]), .B(n25029), .Y(n27982) );
  NOR2X1 U34891 ( .A(ctrl_ww[0]), .B(ctrl_ww[1]), .Y(n25589) );
  AOI22X1 U34892 ( .A(n34083), .B(n26779), .C(n28038), .D(n31804), .Y(n39402)
         );
  NAND2X1 U34893 ( .A(n39438), .B(n39439), .Y(n31804) );
  AOI22X1 U34894 ( .A(reg_A[6]), .B(n26733), .C(reg_A[5]), .D(n25172), .Y(
        n39439) );
  AOI22X1 U34895 ( .A(n26734), .B(reg_A[7]), .C(n25116), .D(reg_A[4]), .Y(
        n39438) );
  INVX1 U34896 ( .A(n32976), .Y(n28038) );
  NAND2X1 U34897 ( .A(n25604), .B(n26691), .Y(n32976) );
  NOR2X1 U34898 ( .A(n26723), .B(reg_B[12]), .Y(n26691) );
  INVX1 U34899 ( .A(reg_B[13]), .Y(n26723) );
  NAND2X1 U34900 ( .A(n39440), .B(n39441), .Y(n26779) );
  AOI22X1 U34901 ( .A(reg_A[14]), .B(n26733), .C(reg_A[13]), .D(n25172), .Y(
        n39441) );
  INVX1 U34902 ( .A(n26731), .Y(n25172) );
  NAND2X1 U34903 ( .A(reg_B[15]), .B(n29256), .Y(n26731) );
  INVX1 U34904 ( .A(n25189), .Y(n26733) );
  NAND2X1 U34905 ( .A(reg_B[14]), .B(n29302), .Y(n25189) );
  AOI22X1 U34906 ( .A(reg_A[15]), .B(n26734), .C(n25116), .D(reg_A[12]), .Y(
        n39440) );
  INVX1 U34907 ( .A(n26692), .Y(n25116) );
  NAND2X1 U34908 ( .A(n29256), .B(n29302), .Y(n26692) );
  INVX1 U34909 ( .A(reg_B[15]), .Y(n29302) );
  INVX1 U34910 ( .A(reg_B[14]), .Y(n29256) );
  INVX1 U34911 ( .A(n25194), .Y(n26734) );
  NAND2X1 U34912 ( .A(reg_B[14]), .B(reg_B[15]), .Y(n25194) );
  INVX1 U34913 ( .A(n35274), .Y(n34083) );
  NAND2X1 U34914 ( .A(n35864), .B(n25604), .Y(n35274) );
  NAND2X1 U34915 ( .A(ctrl_ww[1]), .B(n39410), .Y(n25415) );
  INVX1 U34916 ( .A(ctrl_ww[0]), .Y(n39410) );
  AND2X1 U34917 ( .A(reg_B[12]), .B(reg_B[13]), .Y(n35864) );
  NAND3X1 U34918 ( .A(n39401), .B(n39364), .C(n39363), .Y(n25087) );
  NOR3X1 U34919 ( .A(alu_op[1]), .B(alu_op[3]), .C(n39367), .Y(n39363) );
  INVX1 U34920 ( .A(alu_op[0]), .Y(n39367) );
  INVX1 U34921 ( .A(alu_op[4]), .Y(n39364) );
  INVX1 U34922 ( .A(alu_op[2]), .Y(n39401) );
endmodule

