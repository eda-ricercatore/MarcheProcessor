/**
 * This is written by Zhiyang Ong 
 * and Andrew Mattheisen 
 * for EE577b Troy WideWord Processor Project
 */
 
/**
 * Reference:
 * Nestoras Tzartzanis, EE 577B Verilog Example, Jan 25, 1996
 * http://www-scf.usc.edu/~ee577/tutorial/verilog/alu.v
 */

/**
 * Note that all instructions are 32-bits, and that Big-Endian
 * byte and bit labeling is used. Hence, a[0] is the most
 * significant bit, and a[31] is the least significant bit.
 *
 * Use of casex and casez may affect functionality, and produce
 * larger and slower designs that omit the full_case directive
 *
 * Reference:
 * Don Mills and Clifford E. Cummings, "RTL Coding Styles That
 * Yield Simulation and Synthesis Mismatches", SNUG 1999
 *
 * ALU is a combinational logic block without clock signals
 */

`include "control.h"
// ncverilog only
//`include "~/ee577b/syn/src/control.h"
// synthesis only


// Behavioral model for the ALU
module alu(reg_A,reg_B,ctrl_ppp,ctrl_ww,alu_op,result);

	// Output signals...
	// Result from copmputing an arithmetic or logical operation
	output [0:127] result;
	
	
	
	
	// ===============================================================
	// Input signals
	// Input register A
	input [0:127] reg_A;
	// Input register B
	input [0:127] reg_B;
	// Clock signal
	//input clock;
	// Control signal bits - ppp
	input [0:2] ctrl_ppp;
	// Control signal bits - ww
	input [0:1] ctrl_ww;
	/**
	 * Control signal bits - determine which arithmetic or logic
	 * operation to perform
	 */
	input [0:4] alu_op;
	/**
	 * May also include: branch_offset[n:0], is_branch
	 * Size of branch offset is specified in the Instruction Set
	 * Architecture
	 *
	 * The reset signal for the ALU is ignored
	 */
	
	// PARAMETERS
	parameter zero = 1'b0;
	parameter one = 1'b1;

	
	
	
	// ===============================================================
	// Declare "wire" signals:
	//wire FSM_OUTPUT;
	



	
	// ===============================================================
	// Declare "reg" signals: 
	reg [0:127] result;		// Output signals

	
	
	
	// ===============================================================
	
	always @(reg_A or reg_B or ctrl_ppp or ctrl_ww or alu_op)
	begin
		/**
		 * Based on the assigned arithmetic or logic instruction,
		 * carry out the appropriate function on the operands
		 */
		case(alu_op)


//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
			// ================================================
			
			// SLLI instruction
			
			`aluwslli:
			begin
				case(ctrl_ppp)
					`aa:	// aluwslli SLLI `aa
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:15]<={reg_A[9:15],{1'b0}};
								result[16:23]<={reg_A[17:23],{1'b0}};
								result[24:31]<={reg_A[25:31],{1'b0}};
								result[32:39]<={reg_A[33:39],{1'b0}};
								result[40:47]<={reg_A[41:47],{1'b0}};
								result[48:55]<={reg_A[49:55],{1'b0}};
								result[56:63]<={reg_A[57:63],{1'b0}};
								result[64:71]<={reg_A[65:71],{1'b0}};
								result[72:79]<={reg_A[73:79],{1'b0}};
								result[80:87]<={reg_A[81:87],{1'b0}};
								result[88:95]<={reg_A[89:95],{1'b0}};
								result[96:103]<={reg_A[97:103],{1'b0}};
								result[104:111]<={reg_A[105:111],{1'b0}};
								result[112:119]<={reg_A[113:119],{1'b0}};
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:15]<={reg_A[10:15],{2{1'b0}}};
								result[16:23]<={reg_A[18:23],{2{1'b0}}};
								result[24:31]<={reg_A[26:31],{2{1'b0}}};
								result[32:39]<={reg_A[34:39],{2{1'b0}}};
								result[40:47]<={reg_A[42:47],{2{1'b0}}};
								result[48:55]<={reg_A[50:55],{2{1'b0}}};
								result[56:63]<={reg_A[58:63],{2{1'b0}}};
								result[64:71]<={reg_A[66:71],{2{1'b0}}};
								result[72:79]<={reg_A[74:79],{2{1'b0}}};
								result[80:87]<={reg_A[82:87],{2{1'b0}}};
								result[88:95]<={reg_A[90:95],{2{1'b0}}};
								result[96:103]<={reg_A[98:103],{2{1'b0}}};
								result[104:111]<={reg_A[106:111],{2{1'b0}}};
								result[112:119]<={reg_A[114:119],{2{1'b0}}};
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:15]<={reg_A[11:15],{3{1'b0}}};
								result[16:23]<={reg_A[19:23],{3{1'b0}}};
								result[24:31]<={reg_A[27:31],{3{1'b0}}};
								result[32:39]<={reg_A[35:39],{3{1'b0}}};
								result[40:47]<={reg_A[43:47],{3{1'b0}}};
								result[48:55]<={reg_A[51:55],{3{1'b0}}};
								result[56:63]<={reg_A[59:63],{3{1'b0}}};
								result[64:71]<={reg_A[67:71],{3{1'b0}}};
								result[72:79]<={reg_A[75:79],{3{1'b0}}};
								result[80:87]<={reg_A[83:87],{3{1'b0}}};
								result[88:95]<={reg_A[91:95],{3{1'b0}}};
								result[96:103]<={reg_A[99:103],{3{1'b0}}};
								result[104:111]<={reg_A[107:111],{3{1'b0}}};
								result[112:119]<={reg_A[115:119],{3{1'b0}}};
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:15]<={reg_A[12:15],{4{1'b0}}};
								result[16:23]<={reg_A[20:23],{4{1'b0}}};
								result[24:31]<={reg_A[28:31],{4{1'b0}}};
								result[32:39]<={reg_A[36:39],{4{1'b0}}};
								result[40:47]<={reg_A[44:47],{4{1'b0}}};
								result[48:55]<={reg_A[52:55],{4{1'b0}}};
								result[56:63]<={reg_A[60:63],{4{1'b0}}};
								result[64:71]<={reg_A[68:71],{4{1'b0}}};
								result[72:79]<={reg_A[76:79],{4{1'b0}}};
								result[80:87]<={reg_A[84:87],{4{1'b0}}};
								result[88:95]<={reg_A[92:95],{4{1'b0}}};
								result[96:103]<={reg_A[100:103],{4{1'b0}}};
								result[104:111]<={reg_A[108:111],{4{1'b0}}};
								result[112:119]<={reg_A[116:119],{4{1'b0}}};
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:15]<={reg_A[13:15],{5{1'b0}}};
								result[16:23]<={reg_A[21:23],{5{1'b0}}};
								result[24:31]<={reg_A[29:31],{5{1'b0}}};
								result[32:39]<={reg_A[37:39],{5{1'b0}}};
								result[40:47]<={reg_A[45:47],{5{1'b0}}};
								result[48:55]<={reg_A[53:55],{5{1'b0}}};
								result[56:63]<={reg_A[61:63],{5{1'b0}}};
								result[64:71]<={reg_A[69:71],{5{1'b0}}};
								result[72:79]<={reg_A[77:79],{5{1'b0}}};
								result[80:87]<={reg_A[85:87],{5{1'b0}}};
								result[88:95]<={reg_A[93:95],{5{1'b0}}};
								result[96:103]<={reg_A[101:103],{5{1'b0}}};
								result[104:111]<={reg_A[109:111],{5{1'b0}}};
								result[112:119]<={reg_A[117:119],{5{1'b0}}};
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:15]<={reg_A[14:15],{6{1'b0}}};
								result[16:23]<={reg_A[22:23],{6{1'b0}}};
								result[24:31]<={reg_A[30:31],{6{1'b0}}};
								result[32:39]<={reg_A[38:39],{6{1'b0}}};
								result[40:47]<={reg_A[46:47],{6{1'b0}}};
								result[48:55]<={reg_A[54:55],{6{1'b0}}};
								result[56:63]<={reg_A[62:63],{6{1'b0}}};
								result[64:71]<={reg_A[70:71],{6{1'b0}}};
								result[72:79]<={reg_A[78:79],{6{1'b0}}};
								result[80:87]<={reg_A[86:87],{6{1'b0}}};
								result[88:95]<={reg_A[94:95],{6{1'b0}}};
								result[96:103]<={reg_A[102:103],{6{1'b0}}};
								result[104:111]<={reg_A[110:111],{6{1'b0}}};
								result[112:119]<={reg_A[118:119],{6{1'b0}}};
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:15]<={reg_A[15],{7{1'b0}}};
								result[16:23]<={reg_A[23],{7{1'b0}}};
								result[24:31]<={reg_A[31],{7{1'b0}}};
								result[32:39]<={reg_A[39],{7{1'b0}}};
								result[40:47]<={reg_A[47],{7{1'b0}}};
								result[48:55]<={reg_A[55],{7{1'b0}}};
								result[56:63]<={reg_A[63],{7{1'b0}}};
								result[64:71]<={reg_A[71],{7{1'b0}}};
								result[72:79]<={reg_A[79],{7{1'b0}}};
								result[80:87]<={reg_A[87],{7{1'b0}}};
								result[88:95]<={reg_A[95],{7{1'b0}}};
								result[96:103]<={reg_A[103],{7{1'b0}}};
								result[104:111]<={reg_A[111],{7{1'b0}}};
								result[112:119]<={reg_A[119],{7{1'b0}}};
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:31]<={reg_A[17:31],{1'b0}};
								result[32:47]<={reg_A[33:47],{1'b0}};
								result[48:63]<={reg_A[49:63],{1'b0}};
								result[64:79]<={reg_A[65:79],{1'b0}};
								result[80:95]<={reg_A[81:95],{1'b0}};
								result[96:111]<={reg_A[97:111],{1'b0}};
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:31]<={reg_A[18:31],{2{1'b0}}};
								result[32:47]<={reg_A[34:47],{2{1'b0}}};
								result[48:63]<={reg_A[50:63],{2{1'b0}}};
								result[64:79]<={reg_A[66:79],{2{1'b0}}};
								result[80:95]<={reg_A[82:95],{2{1'b0}}};
								result[96:111]<={reg_A[98:111],{2{1'b0}}};
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:31]<={reg_A[19:31],{3{1'b0}}};
								result[32:47]<={reg_A[35:47],{3{1'b0}}};
								result[48:63]<={reg_A[51:63],{3{1'b0}}};
								result[64:79]<={reg_A[67:79],{3{1'b0}}};
								result[80:95]<={reg_A[83:95],{3{1'b0}}};
								result[96:111]<={reg_A[99:111],{3{1'b0}}};
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:31]<={reg_A[20:31],{4{1'b0}}};
								result[32:47]<={reg_A[36:47],{4{1'b0}}};
								result[48:63]<={reg_A[52:63],{4{1'b0}}};
								result[64:79]<={reg_A[68:79],{4{1'b0}}};
								result[80:95]<={reg_A[84:95],{4{1'b0}}};
								result[96:111]<={reg_A[100:111],{4{1'b0}}};
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:31]<={reg_A[21:31],{5{1'b0}}};
								result[32:47]<={reg_A[37:47],{5{1'b0}}};
								result[48:63]<={reg_A[52:63],{5{1'b0}}};
								result[64:79]<={reg_A[69:79],{5{1'b0}}};
								result[80:95]<={reg_A[85:95],{5{1'b0}}};
								result[96:111]<={reg_A[101:111],{5{1'b0}}};
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:31]<={reg_A[22:31],{6{1'b0}}};
								result[32:47]<={reg_A[38:47],{6{1'b0}}};
								result[48:63]<={reg_A[53:63],{6{1'b0}}};
								result[64:79]<={reg_A[70:79],{6{1'b0}}};
								result[80:95]<={reg_A[86:95],{6{1'b0}}};
								result[96:111]<={reg_A[102:111],{6{1'b0}}};
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:31]<={reg_A[23:31],{7{1'b0}}};
								result[32:47]<={reg_A[39:47],{7{1'b0}}};
								result[48:63]<={reg_A[54:63],{7{1'b0}}};
								result[64:79]<={reg_A[71:79],{7{1'b0}}};
								result[80:95]<={reg_A[87:95],{7{1'b0}}};
								result[96:111]<={reg_A[103:111],{7{1'b0}}};
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:31]<={reg_A[24:31],{8{1'b0}}};
								result[32:47]<={reg_A[40:47],{8{1'b0}}};
								result[48:63]<={reg_A[55:63],{8{1'b0}}};
								result[64:79]<={reg_A[72:79],{8{1'b0}}};
								result[80:95]<={reg_A[88:95],{8{1'b0}}};
								result[96:111]<={reg_A[104:111],{8{1'b0}}};
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:31]<={reg_A[25:31],{9{1'b0}}};
								result[32:47]<={reg_A[41:47],{9{1'b0}}};
								result[48:63]<={reg_A[56:63],{9{1'b0}}};
								result[64:79]<={reg_A[73:79],{9{1'b0}}};
								result[80:95]<={reg_A[89:95],{9{1'b0}}};
								result[96:111]<={reg_A[105:111],{9{1'b0}}};
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:31]<={reg_A[26:31],{10{1'b0}}};
								result[32:47]<={reg_A[42:47],{10{1'b0}}};
								result[48:63]<={reg_A[58:63],{10{1'b0}}};
								result[64:79]<={reg_A[74:79],{10{1'b0}}};
								result[80:95]<={reg_A[90:95],{10{1'b0}}};
								result[96:111]<={reg_A[106:111],{10{1'b0}}};
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:31]<={reg_A[27:31],{11{1'b0}}};
								result[32:47]<={reg_A[43:47],{11{1'b0}}};
								result[48:63]<={reg_A[59:63],{11{1'b0}}};
								result[64:79]<={reg_A[75:79],{11{1'b0}}};
								result[80:95]<={reg_A[91:95],{11{1'b0}}};
								result[96:111]<={reg_A[107:111],{11{1'b0}}};
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:31]<={reg_A[28:31],{12{1'b0}}};
								result[32:47]<={reg_A[44:47],{12{1'b0}}};
								result[48:63]<={reg_A[60:63],{12{1'b0}}};
								result[64:79]<={reg_A[76:79],{12{1'b0}}};
								result[80:95]<={reg_A[92:95],{12{1'b0}}};
								result[96:111]<={reg_A[108:111],{12{1'b0}}};
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:31]<={reg_A[29:31],{13{1'b0}}};
								result[32:47]<={reg_A[45:47],{13{1'b0}}};
								result[48:63]<={reg_A[61:63],{13{1'b0}}};
								result[64:79]<={reg_A[77:79],{13{1'b0}}};
								result[80:95]<={reg_A[93:95],{13{1'b0}}};
								result[96:111]<={reg_A[109:111],{13{1'b0}}};
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:31]<={reg_A[30:31],{14{1'b0}}};
								result[32:47]<={reg_A[46:47],{14{1'b0}}};
								result[48:63]<={reg_A[62:63],{14{1'b0}}};
								result[64:79]<={reg_A[78:79],{14{1'b0}}};
								result[80:95]<={reg_A[94:95],{14{1'b0}}};
								result[96:111]<={reg_A[110:111],{14{1'b0}}};
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:31]<={reg_A[31],{15{1'b0}}};
								result[32:47]<={reg_A[47],{15{1'b0}}};
								result[48:63]<={reg_A[63],{15{1'b0}}};
								result[64:79]<={reg_A[79],{15{1'b0}}};
								result[80:95]<={reg_A[95],{15{1'b0}}};
								result[96:111]<={reg_A[111],{15{1'b0}}};
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:63]<={reg_A[33:63],{1'b0}};
								result[64:95]<={reg_A[65:95],{1'b0}};
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:63]<={reg_A[34:63],{2{1'b0}}};
								result[64:95]<={reg_A[66:95],{2{1'b0}}};
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:63]<={reg_A[35:63],{3{1'b0}}};
								result[64:95]<={reg_A[67:95],{3{1'b0}}};
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:63]<={reg_A[36:63],{4{1'b0}}};
								result[64:95]<={reg_A[68:95],{4{1'b0}}};
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:63]<={reg_A[37:63],{5{1'b0}}};
								result[64:95]<={reg_A[69:95],{5{1'b0}}};
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:63]<={reg_A[38:63],{6{1'b0}}};
								result[64:95]<={reg_A[70:95],{6{1'b0}}};
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:63]<={reg_A[39:63],{7{1'b0}}};
								result[64:95]<={reg_A[71:95],{7{1'b0}}};
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:63]<={reg_A[40:63],{8{1'b0}}};
								result[64:95]<={reg_A[72:95],{8{1'b0}}};
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:63]<={reg_A[41:63],{9{1'b0}}};
								result[64:95]<={reg_A[73:95],{9{1'b0}}};
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:63]<={reg_A[42:63],{10{1'b0}}};
								result[64:95]<={reg_A[74:95],{10{1'b0}}};
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:63]<={reg_A[43:63],{11{1'b0}}};
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:63]<={reg_A[44:63],{12{1'b0}}};
								result[64:95]<={reg_A[76:95],{12{1'b0}}};
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:63]<={reg_A[45:63],{13{1'b0}}};
								result[64:95]<={reg_A[77:95],{13{1'b0}}};
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:63]<={reg_A[46:63],{14{1'b0}}};
								result[64:95]<={reg_A[78:95],{14{1'b0}}};
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:63]<={reg_A[47:63],{15{1'b0}}};
								result[64:95]<={reg_A[79:95],{15{1'b0}}};
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:63]<={reg_A[48:63],{16{1'b0}}};
								result[64:95]<={reg_A[80:95],{16{1'b0}}};
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:63]<={reg_A[49:63],{17{1'b0}}};
								result[64:95]<={reg_A[81:95],{17{1'b0}}};
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:63]<={reg_A[50:63],{18{1'b0}}};
								result[64:95]<={reg_A[82:95],{18{1'b0}}};
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:63]<={reg_A[51:63],{19{1'b0}}};
								result[64:95]<={reg_A[83:95],{19{1'b0}}};
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:63]<={reg_A[52:63],{20{1'b0}}};
								result[64:95]<={reg_A[84:95],{20{1'b0}}};
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:63]<={reg_A[53:63],{21{1'b0}}};
								result[64:95]<={reg_A[85:95],{21{1'b0}}};
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:63]<={reg_A[54:63],{22{1'b0}}};
								result[64:95]<={reg_A[86:95],{22{1'b0}}};
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:63]<={reg_A[55:63],{23{1'b0}}};
								result[64:95]<={reg_A[87:95],{23{1'b0}}};
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:63]<={reg_A[56:63],{24{1'b0}}};
								result[64:95]<={reg_A[88:95],{24{1'b0}}};
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:63]<={reg_A[57:63],{25{1'b0}}};
								result[64:95]<={reg_A[89:95],{25{1'b0}}};
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:63]<={reg_A[58:63],{26{1'b0}}};
								result[64:95]<={reg_A[90:95],{26{1'b0}}};
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:63]<={reg_A[59:63],{27{1'b0}}};
								result[64:95]<={reg_A[91:95],{27{1'b0}}};
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:63]<={reg_A[60:63],{28{1'b0}}};
								result[64:95]<={reg_A[92:95],{28{1'b0}}};
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:63]<={reg_A[61:63],{29{1'b0}}};
								result[64:95]<={reg_A[93:95],{29{1'b0}}};
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:63]<={reg_A[62:63],{30{1'b0}}};
								result[64:95]<={reg_A[94:95],{30{1'b0}}};
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:63]<={reg_A[63],{31{1'b0}}};
								result[64:95]<={reg_A[95],{31{1'b0}}};
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end
					

					`uu:	// aluwslli SLLI `uu
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:63]<=reg_A[0:63];
								result[64:127]<=64'd0;
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:15]<={reg_A[9:15],{1'b0}};
								result[16:23]<={reg_A[17:23],{1'b0}};
								result[24:31]<={reg_A[25:31],{1'b0}};
								result[32:39]<={reg_A[33:39],{1'b0}};
								result[40:47]<={reg_A[41:47],{1'b0}};
								result[48:55]<={reg_A[49:55],{1'b0}};
								result[56:63]<={reg_A[57:63],{1'b0}};
								result[64:127]<=64'd0;
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:15]<={reg_A[10:15],{2{1'b0}}};
								result[16:23]<={reg_A[18:23],{2{1'b0}}};
								result[24:31]<={reg_A[26:31],{2{1'b0}}};
								result[32:39]<={reg_A[34:39],{2{1'b0}}};
								result[40:47]<={reg_A[42:47],{2{1'b0}}};
								result[48:55]<={reg_A[50:55],{2{1'b0}}};
								result[56:63]<={reg_A[58:63],{2{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:15]<={reg_A[11:15],{3{1'b0}}};
								result[16:23]<={reg_A[19:23],{3{1'b0}}};
								result[24:31]<={reg_A[27:31],{3{1'b0}}};
								result[32:39]<={reg_A[35:39],{3{1'b0}}};
								result[40:47]<={reg_A[43:47],{3{1'b0}}};
								result[48:55]<={reg_A[51:55],{3{1'b0}}};
								result[56:63]<={reg_A[59:63],{3{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:15]<={reg_A[12:15],{4{1'b0}}};
								result[16:23]<={reg_A[20:23],{4{1'b0}}};
								result[24:31]<={reg_A[28:31],{4{1'b0}}};
								result[32:39]<={reg_A[36:39],{4{1'b0}}};
								result[40:47]<={reg_A[44:47],{4{1'b0}}};
								result[48:55]<={reg_A[52:55],{4{1'b0}}};
								result[56:63]<={reg_A[60:63],{4{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:15]<={reg_A[13:15],{5{1'b0}}};
								result[16:23]<={reg_A[21:23],{5{1'b0}}};
								result[24:31]<={reg_A[29:31],{5{1'b0}}};
								result[32:39]<={reg_A[37:39],{5{1'b0}}};
								result[40:47]<={reg_A[45:47],{5{1'b0}}};
								result[48:55]<={reg_A[53:55],{5{1'b0}}};
								result[56:63]<={reg_A[61:63],{5{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:15]<={reg_A[14:15],{6{1'b0}}};
								result[16:23]<={reg_A[22:23],{6{1'b0}}};
								result[24:31]<={reg_A[30:31],{6{1'b0}}};
								result[32:39]<={reg_A[38:39],{6{1'b0}}};
								result[40:47]<={reg_A[46:47],{6{1'b0}}};
								result[48:55]<={reg_A[54:55],{6{1'b0}}};
								result[56:63]<={reg_A[62:63],{6{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:15]<={reg_A[15],{7{1'b0}}};
								result[16:23]<={reg_A[23],{7{1'b0}}};
								result[24:31]<={reg_A[31],{7{1'b0}}};
								result[32:39]<={reg_A[39],{7{1'b0}}};
								result[40:47]<={reg_A[47],{7{1'b0}}};
								result[48:55]<={reg_A[55],{7{1'b0}}};
								result[56:63]<={reg_A[63],{7{1'b0}}};
								result[64:127]<=64'd0;
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:63]<=reg_A[0:63];
								result[64:127]<=64'd0;
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:31]<={reg_A[17:31],{1'b0}};
								result[32:47]<={reg_A[33:47],{1'b0}};
								result[48:63]<={reg_A[49:63],{1'b0}};
								result[64:127]<=64'd0;
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:31]<={reg_A[18:31],{2{1'b0}}};
								result[32:47]<={reg_A[34:47],{2{1'b0}}};
								result[48:63]<={reg_A[50:63],{2{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:31]<={reg_A[19:31],{3{1'b0}}};
								result[32:47]<={reg_A[35:47],{3{1'b0}}};
								result[48:63]<={reg_A[51:63],{3{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:31]<={reg_A[20:31],{4{1'b0}}};
								result[32:47]<={reg_A[36:47],{4{1'b0}}};
								result[48:63]<={reg_A[52:63],{4{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:31]<={reg_A[21:31],{5{1'b0}}};
								result[32:47]<={reg_A[37:47],{5{1'b0}}};
								result[48:63]<={reg_A[52:63],{5{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:31]<={reg_A[22:31],{6{1'b0}}};
								result[32:47]<={reg_A[38:47],{6{1'b0}}};
								result[48:63]<={reg_A[53:63],{6{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:31]<={reg_A[23:31],{7{1'b0}}};
								result[32:47]<={reg_A[39:47],{7{1'b0}}};
								result[48:63]<={reg_A[54:63],{7{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:31]<={reg_A[24:31],{8{1'b0}}};
								result[32:47]<={reg_A[40:47],{8{1'b0}}};
								result[48:63]<={reg_A[55:63],{8{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:31]<={reg_A[25:31],{9{1'b0}}};
								result[32:47]<={reg_A[41:47],{9{1'b0}}};
								result[48:63]<={reg_A[56:63],{9{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:31]<={reg_A[26:31],{10{1'b0}}};
								result[32:47]<={reg_A[42:47],{10{1'b0}}};
								result[48:63]<={reg_A[58:63],{10{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:31]<={reg_A[27:31],{11{1'b0}}};
								result[32:47]<={reg_A[43:47],{11{1'b0}}};
								result[48:63]<={reg_A[59:63],{11{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:31]<={reg_A[28:31],{12{1'b0}}};
								result[32:47]<={reg_A[44:47],{12{1'b0}}};
								result[48:63]<={reg_A[60:63],{12{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:31]<={reg_A[29:31],{13{1'b0}}};
								result[32:47]<={reg_A[45:47],{13{1'b0}}};
								result[48:63]<={reg_A[61:63],{13{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:31]<={reg_A[30:31],{14{1'b0}}};
								result[32:47]<={reg_A[46:47],{14{1'b0}}};
								result[48:63]<={reg_A[62:63],{14{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:31]<={reg_A[31],{15{1'b0}}};
								result[32:47]<={reg_A[47],{15{1'b0}}};
								result[48:63]<={reg_A[63],{15{1'b0}}};
								result[64:127]<=64'd0;
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:63]<=reg_A[0:63];
								result[64:127]<=64'd0;
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:63]<={reg_A[33:63],{1'b0}};
								result[64:127]<=64'd0;
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:63]<={reg_A[34:63],{2{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:63]<={reg_A[35:63],{3{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:63]<={reg_A[36:63],{4{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:63]<={reg_A[37:63],{5{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:63]<={reg_A[38:63],{6{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:63]<={reg_A[39:63],{7{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:63]<={reg_A[40:63],{8{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:63]<={reg_A[41:63],{9{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:63]<={reg_A[42:63],{10{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:63]<={reg_A[43:63],{11{1'b0}}};
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:63]<={reg_A[44:63],{12{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:63]<={reg_A[45:63],{13{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:63]<={reg_A[46:63],{14{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:63]<={reg_A[47:63],{15{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:63]<={reg_A[48:63],{16{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:63]<={reg_A[49:63],{17{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:63]<={reg_A[50:63],{18{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:63]<={reg_A[51:63],{19{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:63]<={reg_A[52:63],{20{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:63]<={reg_A[53:63],{21{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:63]<={reg_A[54:63],{22{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:63]<={reg_A[55:63],{23{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:63]<={reg_A[56:63],{24{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:63]<={reg_A[57:63],{25{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:63]<={reg_A[58:63],{26{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:63]<={reg_A[59:63],{27{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:63]<={reg_A[60:63],{28{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:63]<={reg_A[61:63],{29{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:63]<={reg_A[62:63],{30{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:63]<={reg_A[63],{31{1'b0}}};
								result[64:127]<=64'd0;
								end
						endcase
						end
					endcase
					end

					`dd:	// aluwslli SLLI `dd
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:63]<=64'd0;
								result[64:127]<=reg_A[64:127];
								end
							3'd1:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[65:71],{1'b0}};
								result[72:79]<={reg_A[73:79],{1'b0}};
								result[80:87]<={reg_A[81:87],{1'b0}};
								result[88:95]<={reg_A[89:95],{1'b0}};
								result[96:103]<={reg_A[97:103],{1'b0}};
								result[104:111]<={reg_A[105:111],{1'b0}};
								result[112:119]<={reg_A[113:119],{1'b0}};
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[66:71],{2{1'b0}}};
								result[72:79]<={reg_A[74:79],{2{1'b0}}};
								result[80:87]<={reg_A[82:87],{2{1'b0}}};
								result[88:95]<={reg_A[90:95],{2{1'b0}}};
								result[96:103]<={reg_A[98:103],{2{1'b0}}};
								result[104:111]<={reg_A[106:111],{2{1'b0}}};
								result[112:119]<={reg_A[114:119],{2{1'b0}}};
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[67:71],{3{1'b0}}};
								result[72:79]<={reg_A[75:79],{3{1'b0}}};
								result[80:87]<={reg_A[83:87],{3{1'b0}}};
								result[88:95]<={reg_A[91:95],{3{1'b0}}};
								result[96:103]<={reg_A[99:103],{3{1'b0}}};
								result[104:111]<={reg_A[107:111],{3{1'b0}}};
								result[112:119]<={reg_A[115:119],{3{1'b0}}};
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[68:71],{4{1'b0}}};
								result[72:79]<={reg_A[76:79],{4{1'b0}}};
								result[80:87]<={reg_A[84:87],{4{1'b0}}};
								result[88:95]<={reg_A[92:95],{4{1'b0}}};
								result[96:103]<={reg_A[100:103],{4{1'b0}}};
								result[104:111]<={reg_A[108:111],{4{1'b0}}};
								result[112:119]<={reg_A[116:119],{4{1'b0}}};
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[69:71],{5{1'b0}}};
								result[72:79]<={reg_A[77:79],{5{1'b0}}};
								result[80:87]<={reg_A[85:87],{5{1'b0}}};
								result[88:95]<={reg_A[93:95],{5{1'b0}}};
								result[96:103]<={reg_A[101:103],{5{1'b0}}};
								result[104:111]<={reg_A[109:111],{5{1'b0}}};
								result[112:119]<={reg_A[117:119],{5{1'b0}}};
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[70:71],{6{1'b0}}};
								result[72:79]<={reg_A[78:79],{6{1'b0}}};
								result[80:87]<={reg_A[86:87],{6{1'b0}}};
								result[88:95]<={reg_A[94:95],{6{1'b0}}};
								result[96:103]<={reg_A[102:103],{6{1'b0}}};
								result[104:111]<={reg_A[110:111],{6{1'b0}}};
								result[112:119]<={reg_A[118:119],{6{1'b0}}};
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[71],{7{1'b0}}};
								result[72:79]<={reg_A[79],{7{1'b0}}};
								result[80:87]<={reg_A[87],{7{1'b0}}};
								result[88:95]<={reg_A[95],{7{1'b0}}};
								result[96:103]<={reg_A[103],{7{1'b0}}};
								result[104:111]<={reg_A[111],{7{1'b0}}};
								result[112:119]<={reg_A[119],{7{1'b0}}};
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:63]<=64'd0;
								result[64:127]<=reg_A[64:127];
								end
							4'd1:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[65:79],{1'b0}};
								result[80:95]<={reg_A[81:95],{1'b0}};
								result[96:111]<={reg_A[97:111],{1'b0}};
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[66:79],{2{1'b0}}};
								result[80:95]<={reg_A[82:95],{2{1'b0}}};
								result[96:111]<={reg_A[98:111],{2{1'b0}}};
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[67:79],{3{1'b0}}};
								result[80:95]<={reg_A[83:95],{3{1'b0}}};
								result[96:111]<={reg_A[99:111],{3{1'b0}}};
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[68:79],{4{1'b0}}};
								result[80:95]<={reg_A[84:95],{4{1'b0}}};
								result[96:111]<={reg_A[100:111],{4{1'b0}}};
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[69:79],{5{1'b0}}};
								result[80:95]<={reg_A[85:95],{5{1'b0}}};
								result[96:111]<={reg_A[101:111],{5{1'b0}}};
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[70:79],{6{1'b0}}};
								result[80:95]<={reg_A[86:95],{6{1'b0}}};
								result[96:111]<={reg_A[102:111],{6{1'b0}}};
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[71:79],{7{1'b0}}};
								result[80:95]<={reg_A[87:95],{7{1'b0}}};
								result[96:111]<={reg_A[103:111],{7{1'b0}}};
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[72:79],{8{1'b0}}};
								result[80:95]<={reg_A[88:95],{8{1'b0}}};
								result[96:111]<={reg_A[104:111],{8{1'b0}}};
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[73:79],{9{1'b0}}};
								result[80:95]<={reg_A[89:95],{9{1'b0}}};
								result[96:111]<={reg_A[105:111],{9{1'b0}}};
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[74:79],{10{1'b0}}};
								result[80:95]<={reg_A[90:95],{10{1'b0}}};
								result[96:111]<={reg_A[106:111],{10{1'b0}}};
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[75:79],{11{1'b0}}};
								result[80:95]<={reg_A[91:95],{11{1'b0}}};
								result[96:111]<={reg_A[107:111],{11{1'b0}}};
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[76:79],{12{1'b0}}};
								result[80:95]<={reg_A[92:95],{12{1'b0}}};
								result[96:111]<={reg_A[108:111],{12{1'b0}}};
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[77:79],{13{1'b0}}};
								result[80:95]<={reg_A[93:95],{13{1'b0}}};
								result[96:111]<={reg_A[109:111],{13{1'b0}}};
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[78:79],{14{1'b0}}};
								result[80:95]<={reg_A[94:95],{14{1'b0}}};
								result[96:111]<={reg_A[110:111],{14{1'b0}}};
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[79],{15{1'b0}}};
								result[80:95]<={reg_A[95],{15{1'b0}}};
								result[96:111]<={reg_A[111],{15{1'b0}}};
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:63]<=64'd0;
								result[64:127]<=reg_A[64:127];
								end
							5'd1:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[65:95],{1'b0}};
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[66:95],{2{1'b0}}};
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[67:95],{3{1'b0}}};
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[68:95],{4{1'b0}}};
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[69:95],{5{1'b0}}};
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[70:95],{6{1'b0}}};
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[71:95],{7{1'b0}}};
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[72:95],{8{1'b0}}};
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[73:95],{9{1'b0}}};
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[74:95],{10{1'b0}}};
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[76:95],{12{1'b0}}};
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[77:95],{13{1'b0}}};
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[78:95],{14{1'b0}}};
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[79:95],{15{1'b0}}};
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[80:95],{16{1'b0}}};
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[81:95],{17{1'b0}}};
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[82:95],{18{1'b0}}};
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[83:95],{19{1'b0}}};
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[84:95],{20{1'b0}}};
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[85:95],{21{1'b0}}};
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[86:95],{22{1'b0}}};
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[87:95],{23{1'b0}}};
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[88:95],{24{1'b0}}};
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[89:95],{25{1'b0}}};
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[90:95],{26{1'b0}}};
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[91:95],{27{1'b0}}};
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[92:95],{28{1'b0}}};
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[93:95],{29{1'b0}}};
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[94:95],{30{1'b0}}};
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[95],{31{1'b0}}};
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end

					`ee:	// aluwslli SLLI `ee
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:7]<=reg_A[0:7];
								result[8:15]<=8'b0;
								result[16:23]<=reg_A[16:23];
								result[24:31]<=8'b0;
								result[32:39]<=reg_A[33:39];
								result[40:47]<=8'b0;
								result[48:55]<=reg_A[48:55];
								result[56:63]<=8'b0;
								result[64:71]<=reg_A[64:71];
								result[72:79]<=8'b0;
								result[80:87]<=reg_A[80:87];
								result[88:95]<=8'b0;
								result[96:103]<=reg_A[96:103];
								result[104:111]<=8'b0;
								result[112:119]<=reg_A[112:119];
								result[120:127]<=8'b0;
								
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[17:23],{1'b0}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[33:39],{1'b0}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[49:55],{1'b0}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[65:71],{1'b0}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[81:87],{1'b0}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[97:103],{1'b0}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[113:119],{1'b0}};
								result[120:127]<=8'b0;
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[18:23],{2{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[34:39],{2{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[50:55],{2{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[66:71],{2{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[82:87],{2{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[98:103],{2{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[114:119],{2{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[19:23],{3{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[35:39],{3{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[51:55],{3{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[67:71],{3{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[83:87],{3{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[99:103],{3{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[115:119],{3{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[20:23],{4{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[36:39],{4{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[52:55],{4{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[68:71],{4{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[84:87],{4{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[100:103],{4{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[116:119],{4{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[21:23],{5{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[37:39],{5{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[53:55],{5{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[69:71],{5{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[85:87],{5{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[101:103],{5{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[117:119],{5{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[22:23],{6{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[38:39],{6{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[54:55],{6{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[70:71],{6{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[86:87],{6{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[102:103],{6{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[118:119],{6{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[23],{7{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[39],{7{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[55],{7{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[71],{7{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[87],{7{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[103],{7{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[119],{7{1'b0}}};
								result[120:127]<=8'b0;
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[33:47],{1'b0}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[65:79],{1'b0}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[97:111],{1'b0}};
								result[112:127]<=16'b0;
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[34:47],{2{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[66:79],{2{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[98:111],{2{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[35:47],{3{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[67:79],{3{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[99:111],{3{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[36:47],{4{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[68:79],{4{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[100:111],{4{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[37:47],{5{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[69:79],{5{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[101:111],{5{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[38:47],{6{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[70:79],{6{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[102:111],{6{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[39:47],{7{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[71:79],{7{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[103:111],{7{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[40:47],{8{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[72:79],{8{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[104:111],{8{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[41:47],{9{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[73:79],{9{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[105:111],{9{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[42:47],{10{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[74:79],{10{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[106:111],{10{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[43:47],{11{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[75:79],{11{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[107:111],{11{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[44:47],{12{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[76:79],{12{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[108:111],{12{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[45:47],{13{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[77:79],{13{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[109:111],{13{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[46:47],{14{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[78:79],{14{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[110:111],{14{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[47],{15{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[79],{15{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[111],{15{1'b0}}};
								result[112:127]<=16'b0;
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[65:95],{1'b0}};
								result[96:127]<=32'b0;
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[66:95],{2{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[67:95],{3{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[68:95],{4{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[69:95],{5{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[70:95],{6{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[71:95],{7{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[72:95],{8{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[73:95],{9{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[74:95],{10{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[76:95],{12{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[77:95],{13{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[78:95],{14{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[79:95],{15{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[80:95],{16{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[81:95],{17{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[82:95],{18{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[83:95],{19{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[84:95],{20{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[85:95],{21{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[86:95],{22{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[87:95],{23{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[88:95],{24{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[89:95],{25{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[90:95],{26{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[91:95],{27{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[92:95],{28{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[93:95],{29{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[94:95],{30{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[95],{31{1'b0}}};
								result[96:127]<=32'b0;
								end
						endcase
						end
					endcase
					end

					`oo:	// aluwslli SLLI `oo
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							3'd1:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[9:15],{1'b0}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[25:31],{1'b0}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[41:47],{1'b0}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[57:63],{1'b0}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[73:79],{1'b0}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[89:95],{1'b0}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[105:111],{1'b0}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[10:15],{2{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[26:31],{2{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[42:47],{2{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[58:63],{2{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[74:79],{2{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[90:95],{2{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[106:111],{2{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[11:15],{3{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[27:31],{3{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[43:47],{3{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[59:63],{3{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[75:79],{3{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[91:95],{3{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[107:111],{3{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[12:15],{4{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[28:31],{4{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[44:47],{4{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[60:63],{4{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[76:79],{4{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[92:95],{4{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[108:111],{4{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[13:15],{5{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[29:31],{5{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[45:47],{5{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[61:63],{5{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[77:79],{5{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[93:95],{5{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[109:111],{5{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[14:15],{6{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[30:31],{6{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[46:47],{6{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[62:63],{6{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[78:79],{6{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[94:95],{6{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[110:111],{6{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[15],{7{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[31],{7{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[47],{7{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[63],{7{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[79],{7{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[95],{7{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[111],{7{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							4'd1:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[17:31],{1'b0}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[49:63],{1'b0}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[81:95],{1'b0}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[18:31],{2{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[50:63],{2{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[82:95],{2{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[19:31],{3{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[51:63],{3{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[83:95],{3{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[20:31],{4{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[52:63],{4{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[84:95],{4{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[21:31],{5{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[52:63],{5{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[85:95],{5{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[22:31],{6{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[53:63],{6{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[86:95],{6{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[23:31],{7{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[54:63],{7{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[87:95],{7{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[24:31],{8{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[55:63],{8{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[88:95],{8{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[25:31],{9{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[56:63],{9{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[89:95],{9{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[26:31],{10{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[58:63],{10{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[90:95],{10{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[27:31],{11{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[59:63],{11{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[91:95],{11{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[28:31],{12{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[60:63],{12{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[92:95],{12{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[29:31],{13{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[61:63],{13{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[93:95],{13{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[30:31],{14{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[62:63],{14{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[94:95],{14{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[31],{15{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[63],{15{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[95],{15{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							5'd1:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[33:63],{1'b0}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[34:63],{2{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[35:63],{3{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[36:63],{4{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[37:63],{5{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[38:63],{6{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[39:63],{7{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[40:63],{8{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[41:63],{9{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[42:63],{10{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[43:63],{11{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[44:63],{12{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[45:63],{13{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[46:63],{14{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[47:63],{15{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[48:63],{16{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[49:63],{17{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[50:63],{18{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[51:63],{19{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[52:63],{20{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[53:63],{21{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[54:63],{22{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[55:63],{23{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[56:63],{24{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[57:63],{25{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[58:63],{26{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[59:63],{27{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[60:63],{28{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[61:63],{29{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[62:63],{30{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[63],{31{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end

					`mm:	// aluwslli SLLI `mm
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:7]<=reg_A[0:7];
								result[8:127]<=119'b0;
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:127]<=119'b0;
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:127]<=119'b0;
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:15]<=reg_A[0:15];
								result[16:127]<=112'b0;
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:127]<=112'b0;
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:127]<=112'b0;
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:31]<=reg_A[0:31];
								result[32:127]<=96'b0;
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:127]<=96'b0;
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:127]<=96'b0;
								end
						endcase
						end
					endcase
					end

					`ll:	// aluwslli SLLI `ll
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:119]<=120'b0;
								result[120:127]<=reg_A[120:127];
								end
							3'd1:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:111]<=112'b0;
								result[112:127]<=reg_A[112:127];
								end
							4'd1:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:95]<=96'b0;
								result[96:127]<=reg_A[96:127];
								end
							5'd1:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end
				endcase
			end

			// ================================================
			
			// PRM instruction
			
			`aluwprm:
			begin
				case(ctrl_ppp)
					`aa:	// aluwprm PRM `aa
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase

						case(reg_B[12:15]) //byte1
						4'd0:
							result[8:15]<=reg_A[0:7];
						4'd1:
							result[8:15]<=reg_A[8:15];
						4'd2:
							result[8:15]<=reg_A[16:23];
						4'd3:
							result[8:15]<=reg_A[24:31];
						4'd4:
							result[8:15]<=reg_A[32:39];
						4'd5:
							result[8:15]<=reg_A[40:47];
						4'd6:
							result[8:15]<=reg_A[48:55];
						4'd7:
							result[8:15]<=reg_A[56:63];
						4'd8:
							result[8:15]<=reg_A[64:71];
						4'd9:
							result[8:15]<=reg_A[72:79];
						4'd10:
							result[8:15]<=reg_A[80:87];
						4'd11:
							result[8:15]<=reg_A[88:95];
						4'd12:
							result[8:15]<=reg_A[96:103];
						4'd13:
							result[8:15]<=reg_A[104:111];
						4'd14:
							result[8:15]<=reg_A[112:119];
						4'd15:
							result[8:15]<=reg_A[120:127];
						endcase

						case(reg_B[20:23]) //byte2
						4'd0:
							result[16:23]<=reg_A[0:7];
						4'd1:
							result[16:23]<=reg_A[8:15];
						4'd2:
							result[16:23]<=reg_A[16:23];
						4'd3:
							result[16:23]<=reg_A[24:31];
						4'd4:
							result[16:23]<=reg_A[32:39];
						4'd5:
							result[16:23]<=reg_A[40:47];
						4'd6:
							result[16:23]<=reg_A[48:55];
						4'd7:
							result[16:23]<=reg_A[56:63];
						4'd8:
							result[16:23]<=reg_A[64:71];
						4'd9:
							result[16:23]<=reg_A[72:79];
						4'd10:
							result[16:23]<=reg_A[80:87];
						4'd11:
							result[16:23]<=reg_A[88:95];
						4'd12:
							result[16:23]<=reg_A[96:103];
						4'd13:
							result[16:23]<=reg_A[104:111];
						4'd14:
							result[16:23]<=reg_A[112:119];
						4'd15:
							result[16:23]<=reg_A[120:127];
						endcase

						case(reg_B[28:31]) //byte3
						4'd0:
							result[24:31]<=reg_A[0:7];
						4'd1:
							result[24:31]<=reg_A[8:15];
						4'd2:
							result[24:31]<=reg_A[16:23];
						4'd3:
							result[24:31]<=reg_A[24:31];
						4'd4:
							result[24:31]<=reg_A[32:39];
						4'd5:
							result[24:31]<=reg_A[40:47];
						4'd6:
							result[24:31]<=reg_A[48:55];
						4'd7:
							result[24:31]<=reg_A[56:63];
						4'd8:
							result[24:31]<=reg_A[64:71];
						4'd9:
							result[24:31]<=reg_A[72:79];
						4'd10:
							result[24:31]<=reg_A[80:87];
						4'd11:
							result[24:31]<=reg_A[88:95];
						4'd12:
							result[24:31]<=reg_A[96:103];
						4'd13:
							result[24:31]<=reg_A[104:111];
						4'd14:
							result[24:31]<=reg_A[112:119];
						4'd15:
							result[24:31]<=reg_A[120:127];
						endcase

						case(reg_B[36:39]) //byte4
						4'd0:
							result[32:39]<=reg_A[0:7];
						4'd1:
							result[32:39]<=reg_A[8:15];
						4'd2:
							result[32:39]<=reg_A[16:23];
						4'd3:
							result[32:39]<=reg_A[24:31];
						4'd4:
							result[32:39]<=reg_A[32:39];
						4'd5:
							result[32:39]<=reg_A[40:47];
						4'd6:
							result[32:39]<=reg_A[48:55];
						4'd7:
							result[32:39]<=reg_A[56:63];
						4'd8:
							result[32:39]<=reg_A[64:71];
						4'd9:
							result[32:39]<=reg_A[72:79];
						4'd10:
							result[32:39]<=reg_A[80:87];
						4'd11:
							result[32:39]<=reg_A[88:95];
						4'd12:
							result[32:39]<=reg_A[96:103];
						4'd13:
							result[32:39]<=reg_A[104:111];
						4'd14:
							result[32:39]<=reg_A[112:119];
						4'd15:
							result[32:39]<=reg_A[120:127];
						endcase

						case(reg_B[44:47]) //byte5
						4'd0:
							result[40:47]<=reg_A[0:7];
						4'd1:
							result[40:47]<=reg_A[8:15];
						4'd2:
							result[40:47]<=reg_A[16:23];
						4'd3:
							result[40:47]<=reg_A[24:31];
						4'd4:
							result[40:47]<=reg_A[32:39];
						4'd5:
							result[40:47]<=reg_A[40:47];
						4'd6:
							result[40:47]<=reg_A[48:55];
						4'd7:
							result[40:47]<=reg_A[56:63];
						4'd8:
							result[40:47]<=reg_A[64:71];
						4'd9:
							result[40:47]<=reg_A[72:79];
						4'd10:
							result[40:47]<=reg_A[80:87];
						4'd11:
							result[40:47]<=reg_A[88:95];
						4'd12:
							result[40:47]<=reg_A[96:103];
						4'd13:
							result[40:47]<=reg_A[104:111];
						4'd14:
							result[40:47]<=reg_A[112:119];
						4'd15:
							result[40:47]<=reg_A[120:127];
						endcase

						case(reg_B[52:55]) //byte6
						4'd0:
							result[48:55]<=reg_A[0:7];
						4'd1:
							result[48:55]<=reg_A[8:15];
						4'd2:
							result[48:55]<=reg_A[16:23];
						4'd3:
							result[48:55]<=reg_A[24:31];
						4'd4:
							result[48:55]<=reg_A[32:39];
						4'd5:
							result[48:55]<=reg_A[40:47];
						4'd6:
							result[48:55]<=reg_A[48:55];
						4'd7:
							result[48:55]<=reg_A[56:63];
						4'd8:
							result[48:55]<=reg_A[64:71];
						4'd9:
							result[48:55]<=reg_A[72:79];
						4'd10:
							result[48:55]<=reg_A[80:87];
						4'd11:
							result[48:55]<=reg_A[88:95];
						4'd12:
							result[48:55]<=reg_A[96:103];
						4'd13:
							result[48:55]<=reg_A[104:111];
						4'd14:
							result[48:55]<=reg_A[112:119];
						4'd15:
							result[48:55]<=reg_A[120:127];
						endcase

						case(reg_B[60:63]) //byte7
						4'd0:
							result[56:63]<=reg_A[0:7];
						4'd1:
							result[56:63]<=reg_A[8:15];
						4'd2:
							result[56:63]<=reg_A[16:23];
						4'd3:
							result[56:63]<=reg_A[24:31];
						4'd4:
							result[56:63]<=reg_A[32:39];
						4'd5:
							result[56:63]<=reg_A[40:47];
						4'd6:
							result[56:63]<=reg_A[48:55];
						4'd7:
							result[56:63]<=reg_A[56:63];
						4'd8:
							result[56:63]<=reg_A[64:71];
						4'd9:
							result[56:63]<=reg_A[72:79];
						4'd10:
							result[56:63]<=reg_A[80:87];
						4'd11:
							result[56:63]<=reg_A[88:95];
						4'd12:
							result[56:63]<=reg_A[96:103];
						4'd13:
							result[56:63]<=reg_A[104:111];
						4'd14:
							result[56:63]<=reg_A[112:119];
						4'd15:
							result[56:63]<=reg_A[120:127];
						endcase

						case(reg_B[68:71]) //byte8
						4'd0:
							result[64:71]<=reg_A[0:7];
						4'd1:
							result[64:71]<=reg_A[8:15];
						4'd2:
							result[64:71]<=reg_A[16:23];
						4'd3:
							result[64:71]<=reg_A[24:31];
						4'd4:
							result[64:71]<=reg_A[32:39];
						4'd5:
							result[64:71]<=reg_A[40:47];
						4'd6:
							result[64:71]<=reg_A[48:55];
						4'd7:
							result[64:71]<=reg_A[56:63];
						4'd8:
							result[64:71]<=reg_A[64:71];
						4'd9:
							result[64:71]<=reg_A[72:79];
						4'd10:
							result[64:71]<=reg_A[80:87];
						4'd11:
							result[64:71]<=reg_A[88:95];
						4'd12:
							result[64:71]<=reg_A[96:103];
						4'd13:
							result[64:71]<=reg_A[104:111];
						4'd14:
							result[64:71]<=reg_A[112:119];
						4'd15:
							result[64:71]<=reg_A[120:127];
						endcase

						case(reg_B[76:79]) //byte9
						4'd0:
							result[72:79]<=reg_A[0:7];
						4'd1:
							result[72:79]<=reg_A[8:15];
						4'd2:
							result[72:79]<=reg_A[16:23];
						4'd3:
							result[72:79]<=reg_A[24:31];
						4'd4:
							result[72:79]<=reg_A[32:39];
						4'd5:
							result[72:79]<=reg_A[40:47];
						4'd6:
							result[72:79]<=reg_A[48:55];
						4'd7:
							result[72:79]<=reg_A[56:63];
						4'd8:
							result[72:79]<=reg_A[64:71];
						4'd9:
							result[72:79]<=reg_A[72:79];
						4'd10:
							result[72:79]<=reg_A[80:87];
						4'd11:
							result[72:79]<=reg_A[88:95];
						4'd12:
							result[72:79]<=reg_A[96:103];
						4'd13:
							result[72:79]<=reg_A[104:111];
						4'd14:
							result[72:79]<=reg_A[112:119];
						4'd15:
							result[72:79]<=reg_A[120:127];
						endcase

						case(reg_B[84:87]) //byte10
						4'd0:
							result[80:87]<=reg_A[0:7];
						4'd1:
							result[80:87]<=reg_A[8:15];
						4'd2:
							result[80:87]<=reg_A[16:23];
						4'd3:
							result[80:87]<=reg_A[24:31];
						4'd4:
							result[80:87]<=reg_A[32:39];
						4'd5:
							result[80:87]<=reg_A[40:47];
						4'd6:
							result[80:87]<=reg_A[48:55];
						4'd7:
							result[80:87]<=reg_A[56:63];
						4'd8:
							result[80:87]<=reg_A[64:71];
						4'd9:
							result[80:87]<=reg_A[72:79];
						4'd10:
							result[80:87]<=reg_A[80:87];
						4'd11:
							result[80:87]<=reg_A[88:95];
						4'd12:
							result[80:87]<=reg_A[96:103];
						4'd13:
							result[80:87]<=reg_A[104:111];
						4'd14:
							result[80:87]<=reg_A[112:119];
						4'd15:
							result[80:87]<=reg_A[120:127];
						endcase

						case(reg_B[92:95]) //byte11
						4'd0:
							result[88:95]<=reg_A[0:7];
						4'd1:
							result[88:95]<=reg_A[8:15];
						4'd2:
							result[88:95]<=reg_A[16:23];
						4'd3:
							result[88:95]<=reg_A[24:31];
						4'd4:
							result[88:95]<=reg_A[32:39];
						4'd5:
							result[88:95]<=reg_A[40:47];
						4'd6:
							result[88:95]<=reg_A[48:55];
						4'd7:
							result[88:95]<=reg_A[56:63];
						4'd8:
							result[88:95]<=reg_A[64:71];
						4'd9:
							result[88:95]<=reg_A[72:79];
						4'd10:
							result[88:95]<=reg_A[80:87];
						4'd11:
							result[88:95]<=reg_A[88:95];
						4'd12:
							result[88:95]<=reg_A[96:103];
						4'd13:
							result[88:95]<=reg_A[104:111];
						4'd14:
							result[88:95]<=reg_A[112:119];
						4'd15:
							result[88:95]<=reg_A[120:127];
						endcase

						case(reg_B[100:103]) //byte12
						4'd0:
							result[96:103]<=reg_A[0:7];
						4'd1:
							result[96:103]<=reg_A[8:15];
						4'd2:
							result[96:103]<=reg_A[16:23];
						4'd3:
							result[96:103]<=reg_A[24:31];
						4'd4:
							result[96:103]<=reg_A[32:39];
						4'd5:
							result[96:103]<=reg_A[40:47];
						4'd6:
							result[96:103]<=reg_A[48:55];
						4'd7:
							result[96:103]<=reg_A[56:63];
						4'd8:
							result[96:103]<=reg_A[64:71];
						4'd9:
							result[96:103]<=reg_A[72:79];
						4'd10:
							result[96:103]<=reg_A[80:87];
						4'd11:
							result[96:103]<=reg_A[88:95];
						4'd12:
							result[96:103]<=reg_A[96:103];
						4'd13:
							result[96:103]<=reg_A[104:111];
						4'd14:
							result[96:103]<=reg_A[112:119];
						4'd15:
							result[96:103]<=reg_A[120:127];
						endcase

						case(reg_B[108:111]) //byte13
						4'd0:
							result[104:111]<=reg_A[0:7];
						4'd1:
							result[104:111]<=reg_A[8:15];
						4'd2:
							result[104:111]<=reg_A[16:23];
						4'd3:
							result[104:111]<=reg_A[24:31];
						4'd4:
							result[104:111]<=reg_A[32:39];
						4'd5:
							result[104:111]<=reg_A[40:47];
						4'd6:
							result[104:111]<=reg_A[48:55];
						4'd7:
							result[104:111]<=reg_A[56:63];
						4'd8:
							result[104:111]<=reg_A[64:71];
						4'd9:
							result[104:111]<=reg_A[72:79];
						4'd10:
							result[104:111]<=reg_A[80:87];
						4'd11:
							result[104:111]<=reg_A[88:95];
						4'd12:
							result[104:111]<=reg_A[96:103];
						4'd13:
							result[104:111]<=reg_A[104:111];
						4'd14:
							result[104:111]<=reg_A[112:119];
						4'd15:
							result[104:111]<=reg_A[120:127];
						endcase

						case(reg_B[116:119]) //byte14
						4'd0:
							result[112:119]<=reg_A[112:119];
						4'd1:
							result[112:119]<=reg_A[8:15];
						4'd2:
							result[112:119]<=reg_A[16:23];
						4'd3:
							result[112:119]<=reg_A[24:31];
						4'd4:
							result[112:119]<=reg_A[32:39];
						4'd5:
							result[112:119]<=reg_A[40:47];
						4'd6:
							result[112:119]<=reg_A[48:55];
						4'd7:
							result[112:119]<=reg_A[56:63];
						4'd8:
							result[112:119]<=reg_A[64:71];
						4'd9:
							result[112:119]<=reg_A[72:79];
						4'd10:
							result[112:119]<=reg_A[80:87];
						4'd11:
							result[112:119]<=reg_A[88:95];
						4'd12:
							result[112:119]<=reg_A[96:103];
						4'd13:
							result[112:119]<=reg_A[104:111];
						4'd14:
							result[112:119]<=reg_A[112:119];
						4'd15:
							result[112:119]<=reg_A[120:127];
						endcase

						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					`uu:	// aluwprm PRM `uu
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase

						case(reg_B[12:15]) //byte1
						4'd0:
							result[8:15]<=reg_A[0:7];
						4'd1:
							result[8:15]<=reg_A[8:15];
						4'd2:
							result[8:15]<=reg_A[16:23];
						4'd3:
							result[8:15]<=reg_A[24:31];
						4'd4:
							result[8:15]<=reg_A[32:39];
						4'd5:
							result[8:15]<=reg_A[40:47];
						4'd6:
							result[8:15]<=reg_A[48:55];
						4'd7:
							result[8:15]<=reg_A[56:63];
						4'd8:
							result[8:15]<=reg_A[64:71];
						4'd9:
							result[8:15]<=reg_A[72:79];
						4'd10:
							result[8:15]<=reg_A[80:87];
						4'd11:
							result[8:15]<=reg_A[88:95];
						4'd12:
							result[8:15]<=reg_A[96:103];
						4'd13:
							result[8:15]<=reg_A[104:111];
						4'd14:
							result[8:15]<=reg_A[112:119];
						4'd15:
							result[8:15]<=reg_A[120:127];
						endcase

						case(reg_B[20:23]) //byte2
						4'd0:
							result[16:23]<=reg_A[0:7];
						4'd1:
							result[16:23]<=reg_A[8:15];
						4'd2:
							result[16:23]<=reg_A[16:23];
						4'd3:
							result[16:23]<=reg_A[24:31];
						4'd4:
							result[16:23]<=reg_A[32:39];
						4'd5:
							result[16:23]<=reg_A[40:47];
						4'd6:
							result[16:23]<=reg_A[48:55];
						4'd7:
							result[16:23]<=reg_A[56:63];
						4'd8:
							result[16:23]<=reg_A[64:71];
						4'd9:
							result[16:23]<=reg_A[72:79];
						4'd10:
							result[16:23]<=reg_A[80:87];
						4'd11:
							result[16:23]<=reg_A[88:95];
						4'd12:
							result[16:23]<=reg_A[96:103];
						4'd13:
							result[16:23]<=reg_A[104:111];
						4'd14:
							result[16:23]<=reg_A[112:119];
						4'd15:
							result[16:23]<=reg_A[120:127];
						endcase

						case(reg_B[28:31]) //byte3
						4'd0:
							result[24:31]<=reg_A[0:7];
						4'd1:
							result[24:31]<=reg_A[8:15];
						4'd2:
							result[24:31]<=reg_A[16:23];
						4'd3:
							result[24:31]<=reg_A[24:31];
						4'd4:
							result[24:31]<=reg_A[32:39];
						4'd5:
							result[24:31]<=reg_A[40:47];
						4'd6:
							result[24:31]<=reg_A[48:55];
						4'd7:
							result[24:31]<=reg_A[56:63];
						4'd8:
							result[24:31]<=reg_A[64:71];
						4'd9:
							result[24:31]<=reg_A[72:79];
						4'd10:
							result[24:31]<=reg_A[80:87];
						4'd11:
							result[24:31]<=reg_A[88:95];
						4'd12:
							result[24:31]<=reg_A[96:103];
						4'd13:
							result[24:31]<=reg_A[104:111];
						4'd14:
							result[24:31]<=reg_A[112:119];
						4'd15:
							result[24:31]<=reg_A[120:127];
						endcase

						case(reg_B[36:39]) //byte4
						4'd0:
							result[32:39]<=reg_A[0:7];
						4'd1:
							result[32:39]<=reg_A[8:15];
						4'd2:
							result[32:39]<=reg_A[16:23];
						4'd3:
							result[32:39]<=reg_A[24:31];
						4'd4:
							result[32:39]<=reg_A[32:39];
						4'd5:
							result[32:39]<=reg_A[40:47];
						4'd6:
							result[32:39]<=reg_A[48:55];
						4'd7:
							result[32:39]<=reg_A[56:63];
						4'd8:
							result[32:39]<=reg_A[64:71];
						4'd9:
							result[32:39]<=reg_A[72:79];
						4'd10:
							result[32:39]<=reg_A[80:87];
						4'd11:
							result[32:39]<=reg_A[88:95];
						4'd12:
							result[32:39]<=reg_A[96:103];
						4'd13:
							result[32:39]<=reg_A[104:111];
						4'd14:
							result[32:39]<=reg_A[112:119];
						4'd15:
							result[32:39]<=reg_A[120:127];
						endcase

						case(reg_B[44:47]) //byte5
						4'd0:
							result[40:47]<=reg_A[0:7];
						4'd1:
							result[40:47]<=reg_A[8:15];
						4'd2:
							result[40:47]<=reg_A[16:23];
						4'd3:
							result[40:47]<=reg_A[24:31];
						4'd4:
							result[40:47]<=reg_A[32:39];
						4'd5:
							result[40:47]<=reg_A[40:47];
						4'd6:
							result[40:47]<=reg_A[48:55];
						4'd7:
							result[40:47]<=reg_A[56:63];
						4'd8:
							result[40:47]<=reg_A[64:71];
						4'd9:
							result[40:47]<=reg_A[72:79];
						4'd10:
							result[40:47]<=reg_A[80:87];
						4'd11:
							result[40:47]<=reg_A[88:95];
						4'd12:
							result[40:47]<=reg_A[96:103];
						4'd13:
							result[40:47]<=reg_A[104:111];
						4'd14:
							result[40:47]<=reg_A[112:119];
						4'd15:
							result[40:47]<=reg_A[120:127];
						endcase

						case(reg_B[52:55]) //byte6
						4'd0:
							result[48:55]<=reg_A[0:7];
						4'd1:
							result[48:55]<=reg_A[8:15];
						4'd2:
							result[48:55]<=reg_A[16:23];
						4'd3:
							result[48:55]<=reg_A[24:31];
						4'd4:
							result[48:55]<=reg_A[32:39];
						4'd5:
							result[48:55]<=reg_A[40:47];
						4'd6:
							result[48:55]<=reg_A[48:55];
						4'd7:
							result[48:55]<=reg_A[56:63];
						4'd8:
							result[48:55]<=reg_A[64:71];
						4'd9:
							result[48:55]<=reg_A[72:79];
						4'd10:
							result[48:55]<=reg_A[80:87];
						4'd11:
							result[48:55]<=reg_A[88:95];
						4'd12:
							result[48:55]<=reg_A[96:103];
						4'd13:
							result[48:55]<=reg_A[104:111];
						4'd14:
							result[48:55]<=reg_A[112:119];
						4'd15:
							result[48:55]<=reg_A[120:127];
						endcase

						case(reg_B[60:63]) //byte7
						4'd0:
							result[56:63]<=reg_A[0:7];
						4'd1:
							result[56:63]<=reg_A[8:15];
						4'd2:
							result[56:63]<=reg_A[16:23];
						4'd3:
							result[56:63]<=reg_A[24:31];
						4'd4:
							result[56:63]<=reg_A[32:39];
						4'd5:
							result[56:63]<=reg_A[40:47];
						4'd6:
							result[56:63]<=reg_A[48:55];
						4'd7:
							result[56:63]<=reg_A[56:63];
						4'd8:
							result[56:63]<=reg_A[64:71];
						4'd9:
							result[56:63]<=reg_A[72:79];
						4'd10:
							result[56:63]<=reg_A[80:87];
						4'd11:
							result[56:63]<=reg_A[88:95];
						4'd12:
							result[56:63]<=reg_A[96:103];
						4'd13:
							result[56:63]<=reg_A[104:111];
						4'd14:
							result[56:63]<=reg_A[112:119];
						4'd15:
							result[56:63]<=reg_A[120:127];
						endcase

						//bytes8-15
						result[64:127]<=64'd0;
					end
					`dd:	// aluwprm PRM `dd
					begin
						//bytes0-7
						result[0:63]<=64'd0;

						case(reg_B[68:71]) //byte8
						4'd0:
							result[64:71]<=reg_A[0:7];
						4'd1:
							result[64:71]<=reg_A[8:15];
						4'd2:
							result[64:71]<=reg_A[16:23];
						4'd3:
							result[64:71]<=reg_A[24:31];
						4'd4:
							result[64:71]<=reg_A[32:39];
						4'd5:
							result[64:71]<=reg_A[40:47];
						4'd6:
							result[64:71]<=reg_A[48:55];
						4'd7:
							result[64:71]<=reg_A[56:63];
						4'd8:
							result[64:71]<=reg_A[64:71];
						4'd9:
							result[64:71]<=reg_A[72:79];
						4'd10:
							result[64:71]<=reg_A[80:87];
						4'd11:
							result[64:71]<=reg_A[88:95];
						4'd12:
							result[64:71]<=reg_A[96:103];
						4'd13:
							result[64:71]<=reg_A[104:111];
						4'd14:
							result[64:71]<=reg_A[112:119];
						4'd15:
							result[64:71]<=reg_A[120:127];
						endcase

						case(reg_B[76:79]) //byte9
						4'd0:
							result[72:79]<=reg_A[0:7];
						4'd1:
							result[72:79]<=reg_A[8:15];
						4'd2:
							result[72:79]<=reg_A[16:23];
						4'd3:
							result[72:79]<=reg_A[24:31];
						4'd4:
							result[72:79]<=reg_A[32:39];
						4'd5:
							result[72:79]<=reg_A[40:47];
						4'd6:
							result[72:79]<=reg_A[48:55];
						4'd7:
							result[72:79]<=reg_A[56:63];
						4'd8:
							result[72:79]<=reg_A[64:71];
						4'd9:
							result[72:79]<=reg_A[72:79];
						4'd10:
							result[72:79]<=reg_A[80:87];
						4'd11:
							result[72:79]<=reg_A[88:95];
						4'd12:
							result[72:79]<=reg_A[96:103];
						4'd13:
							result[72:79]<=reg_A[104:111];
						4'd14:
							result[72:79]<=reg_A[112:119];
						4'd15:
							result[72:79]<=reg_A[120:127];
						endcase

						case(reg_B[84:87]) //byte10
						4'd0:
							result[80:87]<=reg_A[0:7];
						4'd1:
							result[80:87]<=reg_A[8:15];
						4'd2:
							result[80:87]<=reg_A[16:23];
						4'd3:
							result[80:87]<=reg_A[24:31];
						4'd4:
							result[80:87]<=reg_A[32:39];
						4'd5:
							result[80:87]<=reg_A[40:47];
						4'd6:
							result[80:87]<=reg_A[48:55];
						4'd7:
							result[80:87]<=reg_A[56:63];
						4'd8:
							result[80:87]<=reg_A[64:71];
						4'd9:
							result[80:87]<=reg_A[72:79];
						4'd10:
							result[80:87]<=reg_A[80:87];
						4'd11:
							result[80:87]<=reg_A[88:95];
						4'd12:
							result[80:87]<=reg_A[96:103];
						4'd13:
							result[80:87]<=reg_A[104:111];
						4'd14:
							result[80:87]<=reg_A[112:119];
						4'd15:
							result[80:87]<=reg_A[120:127];
						endcase

						case(reg_B[92:95]) //byte11
						4'd0:
							result[88:95]<=reg_A[0:7];
						4'd1:
							result[88:95]<=reg_A[8:15];
						4'd2:
							result[88:95]<=reg_A[16:23];
						4'd3:
							result[88:95]<=reg_A[24:31];
						4'd4:
							result[88:95]<=reg_A[32:39];
						4'd5:
							result[88:95]<=reg_A[40:47];
						4'd6:
							result[88:95]<=reg_A[48:55];
						4'd7:
							result[88:95]<=reg_A[56:63];
						4'd8:
							result[88:95]<=reg_A[64:71];
						4'd9:
							result[88:95]<=reg_A[72:79];
						4'd10:
							result[88:95]<=reg_A[80:87];
						4'd11:
							result[88:95]<=reg_A[88:95];
						4'd12:
							result[88:95]<=reg_A[96:103];
						4'd13:
							result[88:95]<=reg_A[104:111];
						4'd14:
							result[88:95]<=reg_A[112:119];
						4'd15:
							result[88:95]<=reg_A[120:127];
						endcase

						case(reg_B[100:103]) //byte12
						4'd0:
							result[96:103]<=reg_A[0:7];
						4'd1:
							result[96:103]<=reg_A[8:15];
						4'd2:
							result[96:103]<=reg_A[16:23];
						4'd3:
							result[96:103]<=reg_A[24:31];
						4'd4:
							result[96:103]<=reg_A[32:39];
						4'd5:
							result[96:103]<=reg_A[40:47];
						4'd6:
							result[96:103]<=reg_A[48:55];
						4'd7:
							result[96:103]<=reg_A[56:63];
						4'd8:
							result[96:103]<=reg_A[64:71];
						4'd9:
							result[96:103]<=reg_A[72:79];
						4'd10:
							result[96:103]<=reg_A[80:87];
						4'd11:
							result[96:103]<=reg_A[88:95];
						4'd12:
							result[96:103]<=reg_A[96:103];
						4'd13:
							result[96:103]<=reg_A[104:111];
						4'd14:
							result[96:103]<=reg_A[112:119];
						4'd15:
							result[96:103]<=reg_A[120:127];
						endcase

						case(reg_B[108:111]) //byte13
						4'd0:
							result[104:111]<=reg_A[0:7];
						4'd1:
							result[104:111]<=reg_A[8:15];
						4'd2:
							result[104:111]<=reg_A[16:23];
						4'd3:
							result[104:111]<=reg_A[24:31];
						4'd4:
							result[104:111]<=reg_A[32:39];
						4'd5:
							result[104:111]<=reg_A[40:47];
						4'd6:
							result[104:111]<=reg_A[48:55];
						4'd7:
							result[104:111]<=reg_A[56:63];
						4'd8:
							result[104:111]<=reg_A[64:71];
						4'd9:
							result[104:111]<=reg_A[72:79];
						4'd10:
							result[104:111]<=reg_A[80:87];
						4'd11:
							result[104:111]<=reg_A[88:95];
						4'd12:
							result[104:111]<=reg_A[96:103];
						4'd13:
							result[104:111]<=reg_A[104:111];
						4'd14:
							result[104:111]<=reg_A[112:119];
						4'd15:
							result[104:111]<=reg_A[120:127];
						endcase

						case(reg_B[116:119]) //byte14
						4'd0:
							result[112:119]<=reg_A[0:7];
						4'd1:
							result[112:119]<=reg_A[8:15];
						4'd2:
							result[112:119]<=reg_A[16:23];
						4'd3:
							result[112:119]<=reg_A[24:31];
						4'd4:
							result[112:119]<=reg_A[32:39];
						4'd5:
							result[112:119]<=reg_A[40:47];
						4'd6:
							result[112:119]<=reg_A[48:55];
						4'd7:
							result[112:119]<=reg_A[56:63];
						4'd8:
							result[112:119]<=reg_A[64:71];
						4'd9:
							result[112:119]<=reg_A[72:79];
						4'd10:
							result[112:119]<=reg_A[80:87];
						4'd11:
							result[112:119]<=reg_A[88:95];
						4'd12:
							result[112:119]<=reg_A[96:103];
						4'd13:
							result[112:119]<=reg_A[104:111];
						4'd14:
							result[112:119]<=reg_A[112:119];
						4'd15:
							result[112:119]<=reg_A[120:127];
						endcase

						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					`ee:	// aluwprm PRM `ee
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase

						//byte1
						result[8:15]<=8'd0;

						case(reg_B[20:23]) //byte2
						4'd0:
							result[16:23]<=reg_A[0:7];
						4'd1:
							result[16:23]<=reg_A[8:15];
						4'd2:
							result[16:23]<=reg_A[16:23];
						4'd3:
							result[16:23]<=reg_A[24:31];
						4'd4:
							result[16:23]<=reg_A[32:39];
						4'd5:
							result[16:23]<=reg_A[40:47];
						4'd6:
							result[16:23]<=reg_A[48:55];
						4'd7:
							result[16:23]<=reg_A[56:63];
						4'd8:
							result[16:23]<=reg_A[64:71];
						4'd9:
							result[16:23]<=reg_A[72:79];
						4'd10:
							result[16:23]<=reg_A[80:87];
						4'd11:
							result[16:23]<=reg_A[88:95];
						4'd12:
							result[16:23]<=reg_A[96:103];
						4'd13:
							result[16:23]<=reg_A[104:111];
						4'd14:
							result[16:23]<=reg_A[112:119];
						4'd15:
							result[16:23]<=reg_A[120:127];
						endcase

						//byte3
						result[24:31]<=8'd0;

						case(reg_B[36:39]) //byte4
						4'd0:
							result[32:39]<=reg_A[0:7];
						4'd1:
							result[32:39]<=reg_A[8:15];
						4'd2:
							result[32:39]<=reg_A[16:23];
						4'd3:
							result[32:39]<=reg_A[24:31];
						4'd4:
							result[32:39]<=reg_A[32:39];
						4'd5:
							result[32:39]<=reg_A[40:47];
						4'd6:
							result[32:39]<=reg_A[48:55];
						4'd7:
							result[32:39]<=reg_A[56:63];
						4'd8:
							result[32:39]<=reg_A[64:71];
						4'd9:
							result[32:39]<=reg_A[72:79];
						4'd10:
							result[32:39]<=reg_A[80:87];
						4'd11:
							result[32:39]<=reg_A[88:95];
						4'd12:
							result[32:39]<=reg_A[96:103];
						4'd13:
							result[32:39]<=reg_A[104:111];
						4'd14:
							result[32:39]<=reg_A[112:119];
						4'd15:
							result[32:39]<=reg_A[120:127];
						endcase

						//byte5
						result[40:47]<=8'd0;

						case(reg_B[52:55]) //byte6
						4'd0:
							result[48:55]<=reg_A[0:7];
						4'd1:
							result[48:55]<=reg_A[8:15];
						4'd2:
							result[48:55]<=reg_A[16:23];
						4'd3:
							result[48:55]<=reg_A[24:31];
						4'd4:
							result[48:55]<=reg_A[32:39];
						4'd5:
							result[48:55]<=reg_A[40:47];
						4'd6:
							result[48:55]<=reg_A[48:55];
						4'd7:
							result[48:55]<=reg_A[56:63];
						4'd8:
							result[48:55]<=reg_A[64:71];
						4'd9:
							result[48:55]<=reg_A[72:79];
						4'd10:
							result[48:55]<=reg_A[80:87];
						4'd11:
							result[48:55]<=reg_A[88:95];
						4'd12:
							result[48:55]<=reg_A[96:103];
						4'd13:
							result[48:55]<=reg_A[104:111];
						4'd14:
							result[48:55]<=reg_A[112:119];
						4'd15:
							result[48:55]<=reg_A[120:127];
						endcase

						//byte7
						result[56:63]<=8'd0;

						case(reg_B[68:71]) //byte8
						4'd0:
							result[64:71]<=reg_A[0:7];
						4'd1:
							result[64:71]<=reg_A[8:15];
						4'd2:
							result[64:71]<=reg_A[16:23];
						4'd3:
							result[64:71]<=reg_A[24:31];
						4'd4:
							result[64:71]<=reg_A[32:39];
						4'd5:
							result[64:71]<=reg_A[40:47];
						4'd6:
							result[64:71]<=reg_A[48:55];
						4'd7:
							result[64:71]<=reg_A[56:63];
						4'd8:
							result[64:71]<=reg_A[64:71];
						4'd9:
							result[64:71]<=reg_A[72:79];
						4'd10:
							result[64:71]<=reg_A[80:87];
						4'd11:
							result[64:71]<=reg_A[88:95];
						4'd12:
							result[64:71]<=reg_A[96:103];
						4'd13:
							result[64:71]<=reg_A[104:111];
						4'd14:
							result[64:71]<=reg_A[112:119];
						4'd15:
							result[64:71]<=reg_A[120:127];
						endcase

						//byte9
						result[72:79]<=8'd0;

						case(reg_B[84:87]) //byte10
						4'd0:
							result[80:87]<=reg_A[0:7];
						4'd1:
							result[80:87]<=reg_A[8:15];
						4'd2:
							result[80:87]<=reg_A[16:23];
						4'd3:
							result[80:87]<=reg_A[24:31];
						4'd4:
							result[80:87]<=reg_A[32:39];
						4'd5:
							result[80:87]<=reg_A[40:47];
						4'd6:
							result[80:87]<=reg_A[48:55];
						4'd7:
							result[80:87]<=reg_A[56:63];
						4'd8:
							result[80:87]<=reg_A[64:71];
						4'd9:
							result[80:87]<=reg_A[72:79];
						4'd10:
							result[80:87]<=reg_A[80:87];
						4'd11:
							result[80:87]<=reg_A[88:95];
						4'd12:
							result[80:87]<=reg_A[96:103];
						4'd13:
							result[80:87]<=reg_A[104:111];
						4'd14:
							result[80:87]<=reg_A[112:119];
						4'd15:
							result[80:87]<=reg_A[120:127];
						endcase

						//byte11
						result[88:95]<=8'd0;

						case(reg_B[100:103]) //byte12
						4'd0:
							result[96:103]<=reg_A[0:7];
						4'd1:
							result[96:103]<=reg_A[8:15];
						4'd2:
							result[96:103]<=reg_A[16:23];
						4'd3:
							result[96:103]<=reg_A[24:31];
						4'd4:
							result[96:103]<=reg_A[32:39];
						4'd5:
							result[96:103]<=reg_A[40:47];
						4'd6:
							result[96:103]<=reg_A[48:55];
						4'd7:
							result[96:103]<=reg_A[56:63];
						4'd8:
							result[96:103]<=reg_A[64:71];
						4'd9:
							result[96:103]<=reg_A[72:79];
						4'd10:
							result[96:103]<=reg_A[80:87];
						4'd11:
							result[96:103]<=reg_A[88:95];
						4'd12:
							result[96:103]<=reg_A[96:103];
						4'd13:
							result[96:103]<=reg_A[104:111];
						4'd14:
							result[96:103]<=reg_A[112:119];
						4'd15:
							result[96:103]<=reg_A[120:127];
						endcase

						//byte13
						result[104:111]<=8'd0;

						case(reg_B[116:119]) //byte14
						4'd0:
							result[112:119]<=reg_A[112:119];
						4'd1:
							result[112:119]<=reg_A[8:15];
						4'd2:
							result[112:119]<=reg_A[16:23];
						4'd3:
							result[112:119]<=reg_A[24:31];
						4'd4:
							result[112:119]<=reg_A[32:39];
						4'd5:
							result[112:119]<=reg_A[40:47];
						4'd6:
							result[112:119]<=reg_A[48:55];
						4'd7:
							result[112:119]<=reg_A[56:63];
						4'd8:
							result[112:119]<=reg_A[64:71];
						4'd9:
							result[112:119]<=reg_A[72:79];
						4'd10:
							result[112:119]<=reg_A[80:87];
						4'd11:
							result[112:119]<=reg_A[88:95];
						4'd12:
							result[112:119]<=reg_A[96:103];
						4'd13:
							result[112:119]<=reg_A[104:111];
						4'd14:
							result[112:119]<=reg_A[112:119];
						4'd15:
							result[112:119]<=reg_A[120:127];
						endcase

						//byte15
						result[120:127]<=8'd0;

					end
					`oo:	// aluwprm PRM `oo
					begin
						//byte0
						result[0:7]<=8'd0;

						case(reg_B[12:15]) //byte1
						4'd0:
							result[8:15]<=reg_A[0:7];
						4'd1:
							result[8:15]<=reg_A[8:15];
						4'd2:
							result[8:15]<=reg_A[16:23];
						4'd3:
							result[8:15]<=reg_A[24:31];
						4'd4:
							result[8:15]<=reg_A[32:39];
						4'd5:
							result[8:15]<=reg_A[40:47];
						4'd6:
							result[8:15]<=reg_A[48:55];
						4'd7:
							result[8:15]<=reg_A[56:63];
						4'd8:
							result[8:15]<=reg_A[64:71];
						4'd9:
							result[8:15]<=reg_A[72:79];
						4'd10:
							result[8:15]<=reg_A[80:87];
						4'd11:
							result[8:15]<=reg_A[88:95];
						4'd12:
							result[8:15]<=reg_A[96:103];
						4'd13:
							result[8:15]<=reg_A[104:111];
						4'd14:
							result[8:15]<=reg_A[112:119];
						4'd15:
							result[8:15]<=reg_A[120:127];
						endcase

						//byte2
						result[16:23]<=8'd0;

						case(reg_B[28:31]) //byte3
						4'd0:
							result[24:31]<=reg_A[0:7];
						4'd1:
							result[24:31]<=reg_A[8:15];
						4'd2:
							result[24:31]<=reg_A[16:23];
						4'd3:
							result[24:31]<=reg_A[24:31];
						4'd4:
							result[24:31]<=reg_A[32:39];
						4'd5:
							result[24:31]<=reg_A[40:47];
						4'd6:
							result[24:31]<=reg_A[48:55];
						4'd7:
							result[24:31]<=reg_A[56:63];
						4'd8:
							result[24:31]<=reg_A[64:71];
						4'd9:
							result[24:31]<=reg_A[72:79];
						4'd10:
							result[24:31]<=reg_A[80:87];
						4'd11:
							result[24:31]<=reg_A[88:95];
						4'd12:
							result[24:31]<=reg_A[96:103];
						4'd13:
							result[24:31]<=reg_A[104:111];
						4'd14:
							result[24:31]<=reg_A[112:119];
						4'd15:
							result[24:31]<=reg_A[120:127];
						endcase

						//byte4
						result[32:39]<=8'd0;

						case(reg_B[44:47]) //byte5
						4'd0:
							result[40:47]<=reg_A[0:7];
						4'd1:
							result[40:47]<=reg_A[8:15];
						4'd2:
							result[40:47]<=reg_A[16:23];
						4'd3:
							result[40:47]<=reg_A[24:31];
						4'd4:
							result[40:47]<=reg_A[32:39];
						4'd5:
							result[40:47]<=reg_A[40:47];
						4'd6:
							result[40:47]<=reg_A[48:55];
						4'd7:
							result[40:47]<=reg_A[56:63];
						4'd8:
							result[40:47]<=reg_A[64:71];
						4'd9:
							result[40:47]<=reg_A[72:79];
						4'd10:
							result[40:47]<=reg_A[80:87];
						4'd11:
							result[40:47]<=reg_A[88:95];
						4'd12:
							result[40:47]<=reg_A[96:103];
						4'd13:
							result[40:47]<=reg_A[104:111];
						4'd14:
							result[40:47]<=reg_A[112:119];
						4'd15:
							result[40:47]<=reg_A[120:127];
						endcase

						//byte6
						result[48:55]<=8'd0;

						case(reg_B[60:63]) //byte7
						4'd0:
							result[56:63]<=reg_A[0:7];
						4'd1:
							result[56:63]<=reg_A[8:15];
						4'd2:
							result[56:63]<=reg_A[16:23];
						4'd3:
							result[56:63]<=reg_A[24:31];
						4'd4:
							result[56:63]<=reg_A[32:39];
						4'd5:
							result[56:63]<=reg_A[40:47];
						4'd6:
							result[56:63]<=reg_A[48:55];
						4'd7:
							result[56:63]<=reg_A[56:63];
						4'd8:
							result[56:63]<=reg_A[64:71];
						4'd9:
							result[56:63]<=reg_A[72:79];
						4'd10:
							result[56:63]<=reg_A[80:87];
						4'd11:
							result[56:63]<=reg_A[88:95];
						4'd12:
							result[56:63]<=reg_A[96:103];
						4'd13:
							result[56:63]<=reg_A[104:111];
						4'd14:
							result[56:63]<=reg_A[112:119];
						4'd15:
							result[56:63]<=reg_A[120:127];
						endcase

						//byte8
						result[64:71]<=8'd0;

						case(reg_B[76:79]) //byte9
						4'd0:
							result[72:79]<=reg_A[0:7];
						4'd1:
							result[72:79]<=reg_A[8:15];
						4'd2:
							result[72:79]<=reg_A[16:23];
						4'd3:
							result[72:79]<=reg_A[24:31];
						4'd4:
							result[72:79]<=reg_A[32:39];
						4'd5:
							result[72:79]<=reg_A[40:47];
						4'd6:
							result[72:79]<=reg_A[48:55];
						4'd7:
							result[72:79]<=reg_A[56:63];
						4'd8:
							result[72:79]<=reg_A[64:71];
						4'd9:
							result[72:79]<=reg_A[72:79];
						4'd10:
							result[72:79]<=reg_A[80:87];
						4'd11:
							result[72:79]<=reg_A[88:95];
						4'd12:
							result[72:79]<=reg_A[96:103];
						4'd13:
							result[72:79]<=reg_A[104:111];
						4'd14:
							result[72:79]<=reg_A[112:119];
						4'd15:
							result[72:79]<=reg_A[120:127];
						endcase

						//byte10
						result[80:87]<=8'd0;
						
						case(reg_B[92:95]) //byte11
						4'd0:
							result[88:95]<=reg_A[0:7];
						4'd1:
							result[88:95]<=reg_A[8:15];
						4'd2:
							result[88:95]<=reg_A[16:23];
						4'd3:
							result[88:95]<=reg_A[24:31];
						4'd4:
							result[88:95]<=reg_A[32:39];
						4'd5:
							result[88:95]<=reg_A[40:47];
						4'd6:
							result[88:95]<=reg_A[48:55];
						4'd7:
							result[88:95]<=reg_A[56:63];
						4'd8:
							result[88:95]<=reg_A[64:71];
						4'd9:
							result[88:95]<=reg_A[72:79];
						4'd10:
							result[88:95]<=reg_A[80:87];
						4'd11:
							result[88:95]<=reg_A[88:95];
						4'd12:
							result[88:95]<=reg_A[96:103];
						4'd13:
							result[88:95]<=reg_A[104:111];
						4'd14:
							result[88:95]<=reg_A[112:119];
						4'd15:
							result[88:95]<=reg_A[120:127];
						endcase

						//byte12
						result[96:103]<=8'd0;
						
						case(reg_B[108:111]) //byte13
						4'd0:
							result[104:111]<=reg_A[0:7];
						4'd1:
							result[104:111]<=reg_A[8:15];
						4'd2:
							result[104:111]<=reg_A[16:23];
						4'd3:
							result[104:111]<=reg_A[24:31];
						4'd4:
							result[104:111]<=reg_A[32:39];
						4'd5:
							result[104:111]<=reg_A[40:47];
						4'd6:
							result[104:111]<=reg_A[48:55];
						4'd7:
							result[104:111]<=reg_A[56:63];
						4'd8:
							result[104:111]<=reg_A[64:71];
						4'd9:
							result[104:111]<=reg_A[72:79];
						4'd10:
							result[104:111]<=reg_A[80:87];
						4'd11:
							result[104:111]<=reg_A[88:95];
						4'd12:
							result[104:111]<=reg_A[96:103];
						4'd13:
							result[104:111]<=reg_A[104:111];
						4'd14:
							result[104:111]<=reg_A[112:119];
						4'd15:
							result[104:111]<=reg_A[120:127];
						endcase
						
						//byte14
						result[112:119]<=8'd0;
						
						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					`mm:	// aluwprm PRM `mm
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase
						
						//bytes1-14
						result[8:127]<=120'd0;
						
					end
					`ll:	// aluwprm PRM `ll
					begin
						//bytes0-14
						result[0:119]<=120'd0;
						
						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					default:	// aluwprm PRM Default
					begin
						result<=128'd0;
					end
				endcase
			end


//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================

/*

			// ================================================
			
			// ADD instruction
			
			`aluwadd:
			begin
				case(ctrl_ppp)
					`aa:	// aluwadd AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
								result[8:15]<=reg_A[8:15]+reg_B[8:15];
								result[16:23]<=reg_A[16:23]+reg_B[16:23];
								result[24:31]<=reg_A[24:31]+reg_B[24:31];
								result[32:39]<=reg_A[32:39]+reg_B[32:39];
								result[40:47]<=reg_A[40:47]+reg_B[40:47];
								result[48:55]<=reg_A[48:55]+reg_B[48:55];
								result[56:63]<=reg_A[56:63]+reg_B[56:63];
								result[64:71]<=reg_A[64:71]+reg_B[64:71];
								result[72:79]<=reg_A[72:79]+reg_B[72:79];
								result[80:87]<=reg_A[80:87]+reg_B[80:87];
								result[88:95]<=reg_A[88:95]+reg_B[88:95];
								result[96:103]<=reg_A[96:103]+reg_B[96:103];
								result[104:111]<=reg_A[104:111]+reg_B[104:111];
								result[112:119]<=reg_A[112:119]+reg_B[112:119];
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
								result[16:31]<=reg_A[16:31]+reg_B[16:31];
								result[32:47]<=reg_A[32:47]+reg_B[32:47];
								result[48:63]<=reg_A[48:63]+reg_B[48:63];
								result[64:79]<=reg_A[64:79]+reg_B[64:79];
								result[80:95]<=reg_A[80:95]+reg_B[80:95];
								result[96:111]<=reg_A[96:111]+reg_B[96:111];
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
								result[32:63]<=reg_A[32:63]+reg_B[32:63];
								result[64:95]<=reg_A[64:95]+reg_B[64:95];
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:	// aluwadd AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwadd AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
								result[8:15]<=reg_A[8:15]+reg_B[8:15];
								result[16:23]<=reg_A[16:23]+reg_B[16:23];
								result[24:31]<=reg_A[24:31]+reg_B[24:31];
								result[32:39]<=reg_A[32:39]+reg_B[32:39];
								result[40:47]<=reg_A[40:47]+reg_B[40:47];
								result[48:55]<=reg_A[48:55]+reg_B[48:55];
								result[56:63]<=reg_A[56:63]+reg_B[56:63];
							end
							`w16:	// aluwadd AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
								result[16:31]<=reg_A[16:31]+reg_B[16:31];
								result[32:47]<=reg_A[32:47]+reg_B[32:47];
								result[48:63]<=reg_A[48:63]+reg_B[48:63];
							end
							`w32:	// aluwadd AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
								result[32:63]<=reg_A[32:63]+reg_B[32:63];
							end
							
							default:
							begin
								// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwadd AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]+reg_B[64:71];
								result[72:79]<=reg_A[72:79]+reg_B[72:79];
								result[80:87]<=reg_A[80:87]+reg_B[80:87];
								result[88:95]<=reg_A[88:95]+reg_B[88:95];
								result[96:103]<=reg_A[96:103]+reg_B[96:103];
								result[104:111]<=reg_A[104:111]+reg_B[104:111];
								result[112:119]<=reg_A[112:119]+reg_B[112:119];
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]+reg_B[64:79];
								result[80:95]<=reg_A[80:95]+reg_B[80:95];
								result[96:111]<=reg_A[96:111]+reg_B[96:111];
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]+reg_B[64:95];
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:
							begin
									// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwadd AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
								result[16:23]<=reg_A[16:23]+reg_B[16:23];
								result[32:39]<=reg_A[32:39]+reg_B[32:39];
								result[48:55]<=reg_A[48:55]+reg_B[48:55];
								result[64:71]<=reg_A[64:71]+reg_B[64:71];
								result[80:87]<=reg_A[80:87]+reg_B[80:87];
								result[96:103]<=reg_A[96:103]+reg_B[96:103];
								result[112:119]<=reg_A[112:119]+reg_B[112:119];
							end
							`w16:	// aluwadd AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
								result[32:47]<=reg_A[32:47]+reg_B[32:47];
								result[64:79]<=reg_A[64:79]+reg_B[64:79];
								result[96:111]<=reg_A[96:111]+reg_B[96:111];
							end
							`w32:	// aluwadd AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
								result[64:95]<=reg_A[64:95]+reg_B[64:95];
							end
							
							default:
							begin
								// aluwadd AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwadd AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]+reg_B[8:15];
								result[24:31]<=reg_A[24:31]+reg_B[24:31];
								result[40:47]<=reg_A[40:47]+reg_B[40:47];
								result[56:63]<=reg_A[56:63]+reg_B[56:63];
								result[72:79]<=reg_A[72:79]+reg_B[72:79];
								result[88:95]<=reg_A[88:95]+reg_B[88:95];
								result[104:111]<=reg_A[104:111]+reg_B[104:111];
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]+reg_B[16:31];
								result[48:63]<=reg_A[48:63]+reg_B[48:63];
								result[80:95]<=reg_A[80:95]+reg_B[80:95];
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]+reg_B[32:63];
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwadd AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
							end
							`w16:	// aluwadd AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
							end
							`w32:	// aluwadd AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
							end
							
							default:
							begin
								// aluwadd AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwadd AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwadd AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			// ================================================
			
			// AND instruction
			`aluwand:
			begin
				case(ctrl_ppp)
					`aa:	// aluwadd AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
								result[8:15]<=reg_A[8:15]&reg_B[8:15];
								result[16:23]<=reg_A[16:23]&reg_B[16:23];
								result[24:31]<=reg_A[24:31]&reg_B[24:31];
								result[32:39]<=reg_A[32:39]&reg_B[32:39];
								result[40:47]<=reg_A[40:47]&reg_B[40:47];
								result[48:55]<=reg_A[48:55]&reg_B[48:55];
								result[56:63]<=reg_A[56:63]&reg_B[56:63];
								result[64:71]<=reg_A[64:71]&reg_B[64:71];
								result[72:79]<=reg_A[72:79]&reg_B[72:79];
								result[80:87]<=reg_A[80:87]&reg_B[80:87];
								result[88:95]<=reg_A[88:95]&reg_B[88:95];
								result[96:103]<=reg_A[96:103]&reg_B[96:103];
								result[104:111]<=reg_A[104:111]&reg_B[104:111];
								result[112:119]<=reg_A[112:119]&reg_B[112:119];
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwadd AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
								result[16:31]<=reg_A[16:31]&reg_B[16:31];
								result[32:47]<=reg_A[32:47]&reg_B[32:47];
								result[48:63]<=reg_A[48:63]&reg_B[48:63];
								result[64:79]<=reg_A[64:79]&reg_B[64:79];
								result[80:95]<=reg_A[80:95]&reg_B[80:95];
								result[96:111]<=reg_A[96:111]&reg_B[96:111];
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwadd AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
								result[32:63]<=reg_A[32:63]&reg_B[32:63];
								result[64:95]<=reg_A[64:95]&reg_B[64:95];
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:	// aluwadd AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwadd AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
								result[8:15]<=reg_A[8:15]&reg_B[8:15];
								result[16:23]<=reg_A[16:23]&reg_B[16:23];
								result[24:31]<=reg_A[24:31]&reg_B[24:31];
								result[32:39]<=reg_A[32:39]&reg_B[32:39];
								result[40:47]<=reg_A[40:47]&reg_B[40:47];
								result[48:55]<=reg_A[48:55]&reg_B[48:55];
								result[56:63]<=reg_A[56:63]&reg_B[56:63];
							end
							`w16:	// aluwadd AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
								result[16:31]<=reg_A[16:31]&reg_B[16:31];
								result[32:47]<=reg_A[32:47]&reg_B[32:47];
								result[48:63]<=reg_A[48:63]&reg_B[48:63];
							end
							`w32:	// aluwadd AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
								result[32:63]<=reg_A[32:63]&reg_B[32:63];
							end
							
							default:
							begin
								// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwadd AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]&reg_B[64:71];
								result[72:79]<=reg_A[72:79]&reg_B[72:79];
								result[80:87]<=reg_A[80:87]&reg_B[80:87];
								result[88:95]<=reg_A[88:95]&reg_B[88:95];
								result[96:103]<=reg_A[96:103]&reg_B[96:103];
								result[104:111]<=reg_A[104:111]&reg_B[104:111];
								result[112:119]<=reg_A[112:119]&reg_B[112:119];
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwadd AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]&reg_B[64:79];
								result[80:95]<=reg_A[80:95]&reg_B[80:95];
								result[96:111]<=reg_A[96:111]&reg_B[96:111];
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwadd AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]&reg_B[64:95];
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:
							begin
									// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwadd AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
								result[16:23]<=reg_A[16:23]&reg_B[16:23];
								result[32:39]<=reg_A[32:39]&reg_B[32:39];
								result[48:55]<=reg_A[48:55]&reg_B[48:55];
								result[64:71]<=reg_A[64:71]&reg_B[64:71];
								result[80:87]<=reg_A[80:87]&reg_B[80:87];
								result[96:103]<=reg_A[96:103]&reg_B[96:103];
								result[112:119]<=reg_A[112:119]&reg_B[112:119];
							end
							`w16:	// aluwadd AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
								result[32:47]<=reg_A[32:47]&reg_B[32:47];
								result[64:79]<=reg_A[64:79]&reg_B[64:79];
								result[96:111]<=reg_A[96:111]&reg_B[96:111];
							end
							`w32:	// aluwadd AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
								result[64:95]<=reg_A[64:95]&reg_B[64:95];
							end
							
							default:
							begin
								// aluwadd AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwadd AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]&reg_B[8:15];
								result[24:31]<=reg_A[24:31]&reg_B[24:31];
								result[40:47]<=reg_A[40:47]&reg_B[40:47];
								result[56:63]<=reg_A[56:63]&reg_B[56:63];
								result[72:79]<=reg_A[72:79]&reg_B[72:79];
								result[88:95]<=reg_A[88:95]&reg_B[88:95];
								result[104:111]<=reg_A[104:111]&reg_B[104:111];
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwadd AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]&reg_B[16:31];
								result[48:63]<=reg_A[48:63]&reg_B[48:63];
								result[80:95]<=reg_A[80:95]&reg_B[80:95];
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwadd AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]&reg_B[32:63];
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwadd AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
							end
							`w16:	// aluwadd AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
							end
							`w32:	// aluwadd AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
							end
							
							default:
							begin
								// aluwadd AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwadd AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwadd AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwadd AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwadd AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			// ==============================================
			
			
			// ================================================
			
			// NOT instruction
			`aluwnot:
			begin
				case(ctrl_ppp)
					`aa:	// aluwadd AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `aa AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
								result[8:15]<=~reg_A[8:15];
								result[16:23]<=~reg_A[16:23];
								result[24:31]<=~reg_A[24:31];
								result[32:39]<=~reg_A[32:39];
								result[40:47]<=~reg_A[40:47];
								result[48:55]<=~reg_A[48:55];
								result[56:63]<=~reg_A[56:63];
								result[64:71]<=~reg_A[64:71];
								result[72:79]<=~reg_A[72:79];
								result[80:87]<=~reg_A[80:87];
								result[88:95]<=~reg_A[88:95];
								result[96:103]<=~reg_A[96:103];
								result[104:111]<=~reg_A[104:111];
								result[112:119]<=~reg_A[112:119];
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwadd AND `aa AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
								result[16:31]<=~reg_A[16:31];
								result[32:47]<=~reg_A[32:47];
								result[48:63]<=~reg_A[48:63];
								result[64:79]<=~reg_A[64:79];
								result[80:95]<=~reg_A[80:95];
								result[96:111]<=~reg_A[96:111];
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwadd AND `aa AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
								result[32:63]<=~reg_A[32:63];
								result[64:95]<=~reg_A[64:95];
								result[96:127]<=~reg_A[96:127];
							end
							
							default:	// aluwadd AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwadd AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `uu AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
								result[8:15]<=~reg_A[8:15];
								result[16:23]<=~reg_A[16:23];
								result[24:31]<=~reg_A[24:31];
								result[32:39]<=~reg_A[32:39];
								result[40:47]<=~reg_A[40:47];
								result[48:55]<=~reg_A[48:55];
								result[56:63]<=~reg_A[56:63];
							end
							`w16:	// aluwadd AND `uu AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
								result[16:31]<=~reg_A[16:31];
								result[32:47]<=~reg_A[32:47];
								result[48:63]<=~reg_A[48:63];
							end
							`w32:	// aluwadd AND `uu AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
								result[32:63]<=~reg_A[32:63];
							end
							
							default:
							begin
								// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwadd AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `dd AND `w8
							begin
								result[64:71]<=~reg_A[64:71];
								result[72:79]<=~reg_A[72:79];
								result[80:87]<=~reg_A[80:87];
								result[88:95]<=~reg_A[88:95];
								result[96:103]<=~reg_A[96:103];
								result[104:111]<=~reg_A[104:111];
								result[112:119]<=~reg_A[112:119];
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwadd AND `dd AND `w16
							begin
								result[64:79]<=~reg_A[64:79];
								result[80:95]<=~reg_A[80:95];
								result[96:111]<=~reg_A[96:111];
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwadd AND `dd AND `w32
							begin
								result[64:95]<=~reg_A[64:95];
								result[96:127]<=~reg_A[96:127];
							end
							
							default:
							begin
									// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwadd AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ee AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
								result[16:23]<=~reg_A[16:23];
								result[32:39]<=~reg_A[32:39];
								result[48:55]<=~reg_A[48:55];
								result[64:71]<=~reg_A[64:71];
								result[80:87]<=~reg_A[80:87];
								result[96:103]<=~reg_A[96:103];
								result[112:119]<=~reg_A[112:119];
							end
							`w16:	// aluwadd AND `ee AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
								result[32:47]<=~reg_A[32:47];
								result[64:79]<=~reg_A[64:79];
								result[96:111]<=~reg_A[96:111];
							end
							`w32:	// aluwadd AND `ee AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
								result[64:95]<=~reg_A[64:95];
							end
							
							default:
							begin
								// aluwadd AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwadd AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `oo AND `w8
							begin
								result[8:15]<=~reg_A[8:15];
								result[24:31]<=~reg_A[24:31];
								result[40:47]<=~reg_A[40:47];
								result[56:63]<=~reg_A[56:63];
								result[72:79]<=~reg_A[72:79];
								result[88:95]<=~reg_A[88:95];
								result[104:111]<=~reg_A[104:111];
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwadd AND `oo AND `w16
							begin
								result[16:31]<=~reg_A[16:31];
								result[48:63]<=~reg_A[48:63];
								result[80:95]<=~reg_A[80:95];
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwadd AND `oo AND `w32
							begin
								result[32:63]<=~reg_A[32:63];
								result[96:127]<=~reg_A[96:127];
							end
							
							default:
							begin
								// aluwadd AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwadd AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `mm AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
							end
							`w16:	// aluwadd AND `mm AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
							end
							`w32:	// aluwadd AND `mm AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
							end
							
							default:
							begin
								// aluwadd AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwadd AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ll AND `w8
							begin
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwadd AND `ll AND `w16
							begin
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwadd AND `ll AND `w32
							begin
								result[96:127]<=~reg_A[96:127];
							end
							
							default:
							begin
								// aluwadd AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwadd AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			
			
			// ================================================
			
						// OR instruction
			`aluwor:
			begin
				case(ctrl_ppp)
					`aa:	// aluwadd AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
								result[8:15]<=reg_A[8:15]|reg_B[8:15];
								result[16:23]<=reg_A[16:23]|reg_B[16:23];
								result[24:31]<=reg_A[24:31]|reg_B[24:31];
								result[32:39]<=reg_A[32:39]|reg_B[32:39];
								result[40:47]<=reg_A[40:47]|reg_B[40:47];
								result[48:55]<=reg_A[48:55]|reg_B[48:55];
								result[56:63]<=reg_A[56:63]|reg_B[56:63];
								result[64:71]<=reg_A[64:71]|reg_B[64:71];
								result[72:79]<=reg_A[72:79]|reg_B[72:79];
								result[80:87]<=reg_A[80:87]|reg_B[80:87];
								result[88:95]<=reg_A[88:95]|reg_B[88:95];
								result[96:103]<=reg_A[96:103]|reg_B[96:103];
								result[104:111]<=reg_A[104:111]|reg_B[104:111];
								result[112:119]<=reg_A[112:119]|reg_B[112:119];
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwadd AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
								result[16:31]<=reg_A[16:31]|reg_B[16:31];
								result[32:47]<=reg_A[32:47]|reg_B[32:47];
								result[48:63]<=reg_A[48:63]|reg_B[48:63];
								result[64:79]<=reg_A[64:79]|reg_B[64:79];
								result[80:95]<=reg_A[80:95]|reg_B[80:95];
								result[96:111]<=reg_A[96:111]|reg_B[96:111];
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwadd AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
								result[32:63]<=reg_A[32:63]|reg_B[32:63];
								result[64:95]<=reg_A[64:95]|reg_B[64:95];
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:	// aluwadd AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwadd AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
								result[8:15]<=reg_A[8:15]|reg_B[8:15];
								result[16:23]<=reg_A[16:23]|reg_B[16:23];
								result[24:31]<=reg_A[24:31]|reg_B[24:31];
								result[32:39]<=reg_A[32:39]|reg_B[32:39];
								result[40:47]<=reg_A[40:47]|reg_B[40:47];
								result[48:55]<=reg_A[48:55]|reg_B[48:55];
								result[56:63]<=reg_A[56:63]|reg_B[56:63];
							end
							`w16:	// aluwadd AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
								result[16:31]<=reg_A[16:31]|reg_B[16:31];
								result[32:47]<=reg_A[32:47]|reg_B[32:47];
								result[48:63]<=reg_A[48:63]|reg_B[48:63];
							end
							`w32:	// aluwadd AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
								result[32:63]<=reg_A[32:63]|reg_B[32:63];
							end
							
							default:
							begin
								// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwadd AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]|reg_B[64:71];
								result[72:79]<=reg_A[72:79]|reg_B[72:79];
								result[80:87]<=reg_A[80:87]|reg_B[80:87];
								result[88:95]<=reg_A[88:95]|reg_B[88:95];
								result[96:103]<=reg_A[96:103]|reg_B[96:103];
								result[104:111]<=reg_A[104:111]|reg_B[104:111];
								result[112:119]<=reg_A[112:119]|reg_B[112:119];
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwadd AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]|reg_B[64:79];
								result[80:95]<=reg_A[80:95]|reg_B[80:95];
								result[96:111]<=reg_A[96:111]|reg_B[96:111];
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwadd AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]|reg_B[64:95];
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:
							begin
									// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwadd AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
								result[16:23]<=reg_A[16:23]|reg_B[16:23];
								result[32:39]<=reg_A[32:39]|reg_B[32:39];
								result[48:55]<=reg_A[48:55]|reg_B[48:55];
								result[64:71]<=reg_A[64:71]|reg_B[64:71];
								result[80:87]<=reg_A[80:87]|reg_B[80:87];
								result[96:103]<=reg_A[96:103]|reg_B[96:103];
								result[112:119]<=reg_A[112:119]|reg_B[112:119];
							end
							`w16:	// aluwadd AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
								result[32:47]<=reg_A[32:47]|reg_B[32:47];
								result[64:79]<=reg_A[64:79]|reg_B[64:79];
								result[96:111]<=reg_A[96:111]|reg_B[96:111];
							end
							`w32:	// aluwadd AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
								result[64:95]<=reg_A[64:95]|reg_B[64:95];
							end
							
							default:
							begin
								// aluwadd AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwadd AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]|reg_B[8:15];
								result[24:31]<=reg_A[24:31]|reg_B[24:31];
								result[40:47]<=reg_A[40:47]|reg_B[40:47];
								result[56:63]<=reg_A[56:63]|reg_B[56:63];
								result[72:79]<=reg_A[72:79]|reg_B[72:79];
								result[88:95]<=reg_A[88:95]|reg_B[88:95];
								result[104:111]<=reg_A[104:111]|reg_B[104:111];
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwadd AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]|reg_B[16:31];
								result[48:63]<=reg_A[48:63]|reg_B[48:63];
								result[80:95]<=reg_A[80:95]|reg_B[80:95];
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwadd AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]|reg_B[32:63];
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwadd AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
							end
							`w16:	// aluwadd AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
							end
							`w32:	// aluwadd AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
							end
							
							default:
							begin
								// aluwadd AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwadd AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwadd AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwadd AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwadd AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			
			
*/			
			
			
			
			
			
			
			
			
			
			
			default:
			begin
				// Default arithmetic/logic operation
				result<=128'd0;
			end
		endcase
	end
	
	
	
	
endmodule
