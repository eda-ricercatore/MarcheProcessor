
module alu_DW_mult_uns_1 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176;

  NOR2X1 U17 ( .A(n1), .B(n9), .Y(product[0]) );
  NOR2X1 U18 ( .A(n1), .B(n10), .Y(n17) );
  NOR2X1 U19 ( .A(n1), .B(n11), .Y(n18) );
  NOR2X1 U20 ( .A(n1), .B(n12), .Y(n19) );
  NOR2X1 U21 ( .A(n1), .B(n13), .Y(n20) );
  NOR2X1 U22 ( .A(n1), .B(n14), .Y(n21) );
  NOR2X1 U23 ( .A(n1), .B(n15), .Y(n22) );
  NOR2X1 U24 ( .A(n1), .B(n16), .Y(n23) );
  NOR2X1 U25 ( .A(n2), .B(n9), .Y(n24) );
  NOR2X1 U26 ( .A(n2), .B(n10), .Y(n25) );
  NOR2X1 U27 ( .A(n2), .B(n11), .Y(n26) );
  NOR2X1 U28 ( .A(n2), .B(n12), .Y(n27) );
  NOR2X1 U29 ( .A(n2), .B(n13), .Y(n28) );
  NOR2X1 U30 ( .A(n2), .B(n14), .Y(n29) );
  NOR2X1 U31 ( .A(n2), .B(n15), .Y(n30) );
  NOR2X1 U32 ( .A(n2), .B(n16), .Y(n31) );
  NOR2X1 U33 ( .A(n3), .B(n9), .Y(n32) );
  NOR2X1 U34 ( .A(n3), .B(n10), .Y(n33) );
  NOR2X1 U35 ( .A(n3), .B(n11), .Y(n34) );
  NOR2X1 U36 ( .A(n3), .B(n12), .Y(n35) );
  NOR2X1 U37 ( .A(n3), .B(n13), .Y(n36) );
  NOR2X1 U38 ( .A(n3), .B(n14), .Y(n37) );
  NOR2X1 U39 ( .A(n3), .B(n15), .Y(n38) );
  NOR2X1 U40 ( .A(n3), .B(n16), .Y(n39) );
  NOR2X1 U41 ( .A(n4), .B(n9), .Y(n40) );
  NOR2X1 U42 ( .A(n4), .B(n10), .Y(n41) );
  NOR2X1 U43 ( .A(n4), .B(n11), .Y(n42) );
  NOR2X1 U44 ( .A(n4), .B(n12), .Y(n43) );
  NOR2X1 U45 ( .A(n4), .B(n13), .Y(n44) );
  NOR2X1 U46 ( .A(n4), .B(n14), .Y(n45) );
  NOR2X1 U47 ( .A(n4), .B(n15), .Y(n46) );
  NOR2X1 U48 ( .A(n4), .B(n16), .Y(n47) );
  NOR2X1 U49 ( .A(n5), .B(n9), .Y(n48) );
  NOR2X1 U50 ( .A(n5), .B(n10), .Y(n49) );
  NOR2X1 U51 ( .A(n5), .B(n11), .Y(n50) );
  NOR2X1 U52 ( .A(n5), .B(n12), .Y(n51) );
  NOR2X1 U53 ( .A(n5), .B(n13), .Y(n52) );
  NOR2X1 U54 ( .A(n5), .B(n14), .Y(n53) );
  NOR2X1 U55 ( .A(n5), .B(n15), .Y(n54) );
  NOR2X1 U56 ( .A(n5), .B(n16), .Y(n55) );
  NOR2X1 U57 ( .A(n6), .B(n9), .Y(n56) );
  NOR2X1 U58 ( .A(n6), .B(n10), .Y(n57) );
  NOR2X1 U59 ( .A(n6), .B(n11), .Y(n58) );
  NOR2X1 U60 ( .A(n6), .B(n12), .Y(n59) );
  NOR2X1 U61 ( .A(n6), .B(n13), .Y(n60) );
  NOR2X1 U62 ( .A(n6), .B(n14), .Y(n61) );
  NOR2X1 U63 ( .A(n6), .B(n15), .Y(n62) );
  NOR2X1 U64 ( .A(n6), .B(n16), .Y(n63) );
  NOR2X1 U65 ( .A(n7), .B(n9), .Y(n64) );
  NOR2X1 U66 ( .A(n7), .B(n10), .Y(n65) );
  NOR2X1 U67 ( .A(n7), .B(n11), .Y(n66) );
  NOR2X1 U68 ( .A(n7), .B(n12), .Y(n67) );
  NOR2X1 U69 ( .A(n7), .B(n13), .Y(n68) );
  NOR2X1 U70 ( .A(n7), .B(n14), .Y(n69) );
  NOR2X1 U71 ( .A(n7), .B(n15), .Y(n70) );
  NOR2X1 U72 ( .A(n7), .B(n16), .Y(n71) );
  NOR2X1 U73 ( .A(n8), .B(n9), .Y(n72) );
  NOR2X1 U74 ( .A(n8), .B(n10), .Y(n73) );
  NOR2X1 U75 ( .A(n8), .B(n11), .Y(n74) );
  NOR2X1 U76 ( .A(n8), .B(n12), .Y(n75) );
  NOR2X1 U77 ( .A(n8), .B(n13), .Y(n76) );
  NOR2X1 U78 ( .A(n8), .B(n14), .Y(n77) );
  NOR2X1 U79 ( .A(n8), .B(n15), .Y(n78) );
  NOR2X1 U80 ( .A(n8), .B(n16), .Y(n79) );
  HAX1 U81 ( .A(n18), .B(n25), .YC(n81), .YS(n80) );
  HAX1 U82 ( .A(n33), .B(n40), .YC(n83), .YS(n82) );
  FAX1 U83 ( .A(n19), .B(n26), .C(n81), .YC(n85), .YS(n84) );
  HAX1 U84 ( .A(n41), .B(n48), .YC(n87), .YS(n86) );
  FAX1 U85 ( .A(n20), .B(n34), .C(n27), .YC(n89), .YS(n88) );
  FAX1 U86 ( .A(n83), .B(n86), .C(n88), .YC(n91), .YS(n90) );
  HAX1 U87 ( .A(n49), .B(n56), .YC(n93), .YS(n92) );
  FAX1 U88 ( .A(n21), .B(n42), .C(n35), .YC(n95), .YS(n94) );
  FAX1 U89 ( .A(n28), .B(n87), .C(n92), .YC(n97), .YS(n96) );
  FAX1 U90 ( .A(n89), .B(n94), .C(n96), .YC(n99), .YS(n98) );
  HAX1 U91 ( .A(n57), .B(n64), .YC(n101), .YS(n100) );
  FAX1 U92 ( .A(n22), .B(n50), .C(n29), .YC(n103), .YS(n102) );
  FAX1 U93 ( .A(n36), .B(n43), .C(n93), .YC(n105), .YS(n104) );
  FAX1 U94 ( .A(n100), .B(n95), .C(n102), .YC(n107), .YS(n106) );
  FAX1 U95 ( .A(n97), .B(n104), .C(n106), .YC(n109), .YS(n108) );
  HAX1 U96 ( .A(n65), .B(n72), .YC(n111), .YS(n110) );
  FAX1 U97 ( .A(n23), .B(n58), .C(n30), .YC(n113), .YS(n112) );
  FAX1 U98 ( .A(n37), .B(n51), .C(n44), .YC(n115), .YS(n114) );
  FAX1 U99 ( .A(n101), .B(n110), .C(n103), .YC(n117), .YS(n116) );
  FAX1 U100 ( .A(n114), .B(n112), .C(n105), .YC(n119), .YS(n118) );
  FAX1 U101 ( .A(n107), .B(n116), .C(n118), .YC(n121), .YS(n120) );
  HAX1 U102 ( .A(n66), .B(n73), .YC(n123), .YS(n122) );
  FAX1 U103 ( .A(n52), .B(n59), .C(n31), .YC(n125), .YS(n124) );
  FAX1 U104 ( .A(n38), .B(n45), .C(n111), .YC(n127), .YS(n126) );
  FAX1 U105 ( .A(n122), .B(n113), .C(n115), .YC(n129), .YS(n128) );
  FAX1 U106 ( .A(n124), .B(n126), .C(n117), .YC(n131), .YS(n130) );
  FAX1 U107 ( .A(n128), .B(n119), .C(n130), .YC(n133), .YS(n132) );
  FAX1 U108 ( .A(n39), .B(n74), .C(n67), .YC(n135), .YS(n134) );
  FAX1 U109 ( .A(n60), .B(n53), .C(n46), .YC(n137), .YS(n136) );
  FAX1 U110 ( .A(n123), .B(n125), .C(n136), .YC(n139), .YS(n138) );
  FAX1 U111 ( .A(n134), .B(n127), .C(n129), .YC(n141), .YS(n140) );
  FAX1 U112 ( .A(n138), .B(n131), .C(n140), .YC(n143), .YS(n142) );
  FAX1 U113 ( .A(n47), .B(n75), .C(n68), .YC(n145), .YS(n144) );
  FAX1 U114 ( .A(n54), .B(n61), .C(n135), .YC(n147), .YS(n146) );
  FAX1 U115 ( .A(n137), .B(n144), .C(n139), .YC(n149), .YS(n148) );
  FAX1 U116 ( .A(n146), .B(n141), .C(n148), .YC(n151), .YS(n150) );
  FAX1 U117 ( .A(n55), .B(n76), .C(n69), .YC(n153), .YS(n152) );
  FAX1 U118 ( .A(n62), .B(n145), .C(n152), .YC(n155), .YS(n154) );
  FAX1 U119 ( .A(n147), .B(n154), .C(n149), .YC(n157), .YS(n156) );
  FAX1 U120 ( .A(n63), .B(n77), .C(n70), .YC(n159), .YS(n158) );
  FAX1 U121 ( .A(n153), .B(n158), .C(n155), .YC(n161), .YS(n160) );
  FAX1 U122 ( .A(n71), .B(n78), .C(n159), .YC(n163), .YS(n162) );
  HAX1 U123 ( .A(n24), .B(n17), .YC(n164), .YS(product[1]) );
  FAX1 U124 ( .A(n32), .B(n164), .C(n80), .YC(n165), .YS(product[2]) );
  FAX1 U125 ( .A(n82), .B(n165), .C(n84), .YC(n166), .YS(product[3]) );
  FAX1 U126 ( .A(n85), .B(n90), .C(n166), .YC(n167), .YS(product[4]) );
  FAX1 U127 ( .A(n91), .B(n98), .C(n167), .YC(n168), .YS(product[5]) );
  FAX1 U128 ( .A(n99), .B(n108), .C(n168), .YC(n169), .YS(product[6]) );
  FAX1 U129 ( .A(n109), .B(n120), .C(n169), .YC(n170), .YS(product[7]) );
  FAX1 U130 ( .A(n121), .B(n132), .C(n170), .YC(n171), .YS(product[8]) );
  FAX1 U131 ( .A(n133), .B(n142), .C(n171), .YC(n172), .YS(product[9]) );
  FAX1 U132 ( .A(n143), .B(n150), .C(n172), .YC(n173), .YS(product[10]) );
  FAX1 U133 ( .A(n151), .B(n156), .C(n173), .YC(n174), .YS(product[11]) );
  FAX1 U134 ( .A(n160), .B(n157), .C(n174), .YC(n175), .YS(product[12]) );
  FAX1 U135 ( .A(n162), .B(n161), .C(n175), .YC(n176), .YS(product[13]) );
  FAX1 U136 ( .A(n79), .B(n163), .C(n176), .YC(product[15]), .YS(product[14])
         );
  INVX2 U140 ( .A(b[0]), .Y(n9) );
  INVX2 U141 ( .A(b[1]), .Y(n10) );
  INVX2 U142 ( .A(b[2]), .Y(n11) );
  INVX2 U143 ( .A(b[3]), .Y(n12) );
  INVX2 U144 ( .A(b[4]), .Y(n13) );
  INVX2 U145 ( .A(b[5]), .Y(n14) );
  INVX2 U146 ( .A(b[6]), .Y(n15) );
  INVX2 U147 ( .A(b[7]), .Y(n16) );
  INVX2 U148 ( .A(a[0]), .Y(n1) );
  INVX2 U149 ( .A(a[1]), .Y(n2) );
  INVX2 U150 ( .A(a[2]), .Y(n3) );
  INVX2 U151 ( .A(a[3]), .Y(n4) );
  INVX2 U152 ( .A(a[4]), .Y(n5) );
  INVX2 U153 ( .A(a[5]), .Y(n6) );
  INVX2 U154 ( .A(a[6]), .Y(n7) );
  INVX2 U155 ( .A(a[7]), .Y(n8) );
endmodule


module alu_DW_mult_uns_2 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176;

  NOR2X1 U17 ( .A(n1), .B(n9), .Y(product[0]) );
  NOR2X1 U18 ( .A(n1), .B(n10), .Y(n17) );
  NOR2X1 U19 ( .A(n1), .B(n11), .Y(n18) );
  NOR2X1 U20 ( .A(n1), .B(n12), .Y(n19) );
  NOR2X1 U21 ( .A(n1), .B(n13), .Y(n20) );
  NOR2X1 U22 ( .A(n1), .B(n14), .Y(n21) );
  NOR2X1 U23 ( .A(n1), .B(n15), .Y(n22) );
  NOR2X1 U24 ( .A(n1), .B(n16), .Y(n23) );
  NOR2X1 U25 ( .A(n2), .B(n9), .Y(n24) );
  NOR2X1 U26 ( .A(n2), .B(n10), .Y(n25) );
  NOR2X1 U27 ( .A(n2), .B(n11), .Y(n26) );
  NOR2X1 U28 ( .A(n2), .B(n12), .Y(n27) );
  NOR2X1 U29 ( .A(n2), .B(n13), .Y(n28) );
  NOR2X1 U30 ( .A(n2), .B(n14), .Y(n29) );
  NOR2X1 U31 ( .A(n2), .B(n15), .Y(n30) );
  NOR2X1 U32 ( .A(n2), .B(n16), .Y(n31) );
  NOR2X1 U33 ( .A(n3), .B(n9), .Y(n32) );
  NOR2X1 U34 ( .A(n3), .B(n10), .Y(n33) );
  NOR2X1 U35 ( .A(n3), .B(n11), .Y(n34) );
  NOR2X1 U36 ( .A(n3), .B(n12), .Y(n35) );
  NOR2X1 U37 ( .A(n3), .B(n13), .Y(n36) );
  NOR2X1 U38 ( .A(n3), .B(n14), .Y(n37) );
  NOR2X1 U39 ( .A(n3), .B(n15), .Y(n38) );
  NOR2X1 U40 ( .A(n3), .B(n16), .Y(n39) );
  NOR2X1 U41 ( .A(n4), .B(n9), .Y(n40) );
  NOR2X1 U42 ( .A(n4), .B(n10), .Y(n41) );
  NOR2X1 U43 ( .A(n4), .B(n11), .Y(n42) );
  NOR2X1 U44 ( .A(n4), .B(n12), .Y(n43) );
  NOR2X1 U45 ( .A(n4), .B(n13), .Y(n44) );
  NOR2X1 U46 ( .A(n4), .B(n14), .Y(n45) );
  NOR2X1 U47 ( .A(n4), .B(n15), .Y(n46) );
  NOR2X1 U48 ( .A(n4), .B(n16), .Y(n47) );
  NOR2X1 U49 ( .A(n5), .B(n9), .Y(n48) );
  NOR2X1 U50 ( .A(n5), .B(n10), .Y(n49) );
  NOR2X1 U51 ( .A(n5), .B(n11), .Y(n50) );
  NOR2X1 U52 ( .A(n5), .B(n12), .Y(n51) );
  NOR2X1 U53 ( .A(n5), .B(n13), .Y(n52) );
  NOR2X1 U54 ( .A(n5), .B(n14), .Y(n53) );
  NOR2X1 U55 ( .A(n5), .B(n15), .Y(n54) );
  NOR2X1 U56 ( .A(n5), .B(n16), .Y(n55) );
  NOR2X1 U57 ( .A(n6), .B(n9), .Y(n56) );
  NOR2X1 U58 ( .A(n6), .B(n10), .Y(n57) );
  NOR2X1 U59 ( .A(n6), .B(n11), .Y(n58) );
  NOR2X1 U60 ( .A(n6), .B(n12), .Y(n59) );
  NOR2X1 U61 ( .A(n6), .B(n13), .Y(n60) );
  NOR2X1 U62 ( .A(n6), .B(n14), .Y(n61) );
  NOR2X1 U63 ( .A(n6), .B(n15), .Y(n62) );
  NOR2X1 U64 ( .A(n6), .B(n16), .Y(n63) );
  NOR2X1 U65 ( .A(n7), .B(n9), .Y(n64) );
  NOR2X1 U66 ( .A(n7), .B(n10), .Y(n65) );
  NOR2X1 U67 ( .A(n7), .B(n11), .Y(n66) );
  NOR2X1 U68 ( .A(n7), .B(n12), .Y(n67) );
  NOR2X1 U69 ( .A(n7), .B(n13), .Y(n68) );
  NOR2X1 U70 ( .A(n7), .B(n14), .Y(n69) );
  NOR2X1 U71 ( .A(n7), .B(n15), .Y(n70) );
  NOR2X1 U72 ( .A(n7), .B(n16), .Y(n71) );
  NOR2X1 U73 ( .A(n8), .B(n9), .Y(n72) );
  NOR2X1 U74 ( .A(n8), .B(n10), .Y(n73) );
  NOR2X1 U75 ( .A(n8), .B(n11), .Y(n74) );
  NOR2X1 U76 ( .A(n8), .B(n12), .Y(n75) );
  NOR2X1 U77 ( .A(n8), .B(n13), .Y(n76) );
  NOR2X1 U78 ( .A(n8), .B(n14), .Y(n77) );
  NOR2X1 U79 ( .A(n8), .B(n15), .Y(n78) );
  NOR2X1 U80 ( .A(n8), .B(n16), .Y(n79) );
  HAX1 U81 ( .A(n18), .B(n25), .YC(n81), .YS(n80) );
  HAX1 U82 ( .A(n33), .B(n40), .YC(n83), .YS(n82) );
  FAX1 U83 ( .A(n19), .B(n26), .C(n81), .YC(n85), .YS(n84) );
  HAX1 U84 ( .A(n41), .B(n48), .YC(n87), .YS(n86) );
  FAX1 U85 ( .A(n20), .B(n34), .C(n27), .YC(n89), .YS(n88) );
  FAX1 U86 ( .A(n83), .B(n86), .C(n88), .YC(n91), .YS(n90) );
  HAX1 U87 ( .A(n49), .B(n56), .YC(n93), .YS(n92) );
  FAX1 U88 ( .A(n21), .B(n42), .C(n35), .YC(n95), .YS(n94) );
  FAX1 U89 ( .A(n28), .B(n87), .C(n92), .YC(n97), .YS(n96) );
  FAX1 U90 ( .A(n89), .B(n94), .C(n96), .YC(n99), .YS(n98) );
  HAX1 U91 ( .A(n57), .B(n64), .YC(n101), .YS(n100) );
  FAX1 U92 ( .A(n22), .B(n50), .C(n29), .YC(n103), .YS(n102) );
  FAX1 U93 ( .A(n36), .B(n43), .C(n93), .YC(n105), .YS(n104) );
  FAX1 U94 ( .A(n100), .B(n95), .C(n102), .YC(n107), .YS(n106) );
  FAX1 U95 ( .A(n97), .B(n104), .C(n106), .YC(n109), .YS(n108) );
  HAX1 U96 ( .A(n65), .B(n72), .YC(n111), .YS(n110) );
  FAX1 U97 ( .A(n23), .B(n58), .C(n30), .YC(n113), .YS(n112) );
  FAX1 U98 ( .A(n37), .B(n51), .C(n44), .YC(n115), .YS(n114) );
  FAX1 U99 ( .A(n101), .B(n110), .C(n103), .YC(n117), .YS(n116) );
  FAX1 U100 ( .A(n114), .B(n112), .C(n105), .YC(n119), .YS(n118) );
  FAX1 U101 ( .A(n107), .B(n116), .C(n118), .YC(n121), .YS(n120) );
  HAX1 U102 ( .A(n66), .B(n73), .YC(n123), .YS(n122) );
  FAX1 U103 ( .A(n52), .B(n59), .C(n31), .YC(n125), .YS(n124) );
  FAX1 U104 ( .A(n38), .B(n45), .C(n111), .YC(n127), .YS(n126) );
  FAX1 U105 ( .A(n122), .B(n113), .C(n115), .YC(n129), .YS(n128) );
  FAX1 U106 ( .A(n124), .B(n126), .C(n117), .YC(n131), .YS(n130) );
  FAX1 U107 ( .A(n128), .B(n119), .C(n130), .YC(n133), .YS(n132) );
  FAX1 U108 ( .A(n39), .B(n74), .C(n67), .YC(n135), .YS(n134) );
  FAX1 U109 ( .A(n60), .B(n53), .C(n46), .YC(n137), .YS(n136) );
  FAX1 U110 ( .A(n123), .B(n125), .C(n136), .YC(n139), .YS(n138) );
  FAX1 U111 ( .A(n134), .B(n127), .C(n129), .YC(n141), .YS(n140) );
  FAX1 U112 ( .A(n138), .B(n131), .C(n140), .YC(n143), .YS(n142) );
  FAX1 U113 ( .A(n47), .B(n75), .C(n68), .YC(n145), .YS(n144) );
  FAX1 U114 ( .A(n54), .B(n61), .C(n135), .YC(n147), .YS(n146) );
  FAX1 U115 ( .A(n137), .B(n144), .C(n139), .YC(n149), .YS(n148) );
  FAX1 U116 ( .A(n146), .B(n141), .C(n148), .YC(n151), .YS(n150) );
  FAX1 U117 ( .A(n55), .B(n76), .C(n69), .YC(n153), .YS(n152) );
  FAX1 U118 ( .A(n62), .B(n145), .C(n152), .YC(n155), .YS(n154) );
  FAX1 U119 ( .A(n147), .B(n154), .C(n149), .YC(n157), .YS(n156) );
  FAX1 U120 ( .A(n63), .B(n77), .C(n70), .YC(n159), .YS(n158) );
  FAX1 U121 ( .A(n153), .B(n158), .C(n155), .YC(n161), .YS(n160) );
  FAX1 U122 ( .A(n71), .B(n78), .C(n159), .YC(n163), .YS(n162) );
  HAX1 U123 ( .A(n24), .B(n17), .YC(n164), .YS(product[1]) );
  FAX1 U124 ( .A(n32), .B(n164), .C(n80), .YC(n165), .YS(product[2]) );
  FAX1 U125 ( .A(n82), .B(n165), .C(n84), .YC(n166), .YS(product[3]) );
  FAX1 U126 ( .A(n85), .B(n90), .C(n166), .YC(n167), .YS(product[4]) );
  FAX1 U127 ( .A(n91), .B(n98), .C(n167), .YC(n168), .YS(product[5]) );
  FAX1 U128 ( .A(n99), .B(n108), .C(n168), .YC(n169), .YS(product[6]) );
  FAX1 U129 ( .A(n109), .B(n120), .C(n169), .YC(n170), .YS(product[7]) );
  FAX1 U130 ( .A(n121), .B(n132), .C(n170), .YC(n171), .YS(product[8]) );
  FAX1 U131 ( .A(n133), .B(n142), .C(n171), .YC(n172), .YS(product[9]) );
  FAX1 U132 ( .A(n143), .B(n150), .C(n172), .YC(n173), .YS(product[10]) );
  FAX1 U133 ( .A(n151), .B(n156), .C(n173), .YC(n174), .YS(product[11]) );
  FAX1 U134 ( .A(n160), .B(n157), .C(n174), .YC(n175), .YS(product[12]) );
  FAX1 U135 ( .A(n162), .B(n161), .C(n175), .YC(n176), .YS(product[13]) );
  FAX1 U136 ( .A(n79), .B(n163), .C(n176), .YC(product[15]), .YS(product[14])
         );
  INVX2 U140 ( .A(b[0]), .Y(n9) );
  INVX2 U141 ( .A(b[1]), .Y(n10) );
  INVX2 U142 ( .A(b[2]), .Y(n11) );
  INVX2 U143 ( .A(b[3]), .Y(n12) );
  INVX2 U144 ( .A(b[4]), .Y(n13) );
  INVX2 U145 ( .A(b[5]), .Y(n14) );
  INVX2 U146 ( .A(b[6]), .Y(n15) );
  INVX2 U147 ( .A(b[7]), .Y(n16) );
  INVX2 U148 ( .A(a[0]), .Y(n1) );
  INVX2 U149 ( .A(a[1]), .Y(n2) );
  INVX2 U150 ( .A(a[2]), .Y(n3) );
  INVX2 U151 ( .A(a[3]), .Y(n4) );
  INVX2 U152 ( .A(a[4]), .Y(n5) );
  INVX2 U153 ( .A(a[5]), .Y(n6) );
  INVX2 U154 ( .A(a[6]), .Y(n7) );
  INVX2 U155 ( .A(a[7]), .Y(n8) );
endmodule


module alu_DW_mult_uns_3 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176;

  NOR2X1 U17 ( .A(n1), .B(n9), .Y(product[0]) );
  NOR2X1 U18 ( .A(n1), .B(n10), .Y(n17) );
  NOR2X1 U19 ( .A(n1), .B(n11), .Y(n18) );
  NOR2X1 U20 ( .A(n1), .B(n12), .Y(n19) );
  NOR2X1 U21 ( .A(n1), .B(n13), .Y(n20) );
  NOR2X1 U22 ( .A(n1), .B(n14), .Y(n21) );
  NOR2X1 U23 ( .A(n1), .B(n15), .Y(n22) );
  NOR2X1 U24 ( .A(n1), .B(n16), .Y(n23) );
  NOR2X1 U25 ( .A(n2), .B(n9), .Y(n24) );
  NOR2X1 U26 ( .A(n2), .B(n10), .Y(n25) );
  NOR2X1 U27 ( .A(n2), .B(n11), .Y(n26) );
  NOR2X1 U28 ( .A(n2), .B(n12), .Y(n27) );
  NOR2X1 U29 ( .A(n2), .B(n13), .Y(n28) );
  NOR2X1 U30 ( .A(n2), .B(n14), .Y(n29) );
  NOR2X1 U31 ( .A(n2), .B(n15), .Y(n30) );
  NOR2X1 U32 ( .A(n2), .B(n16), .Y(n31) );
  NOR2X1 U33 ( .A(n3), .B(n9), .Y(n32) );
  NOR2X1 U34 ( .A(n3), .B(n10), .Y(n33) );
  NOR2X1 U35 ( .A(n3), .B(n11), .Y(n34) );
  NOR2X1 U36 ( .A(n3), .B(n12), .Y(n35) );
  NOR2X1 U37 ( .A(n3), .B(n13), .Y(n36) );
  NOR2X1 U38 ( .A(n3), .B(n14), .Y(n37) );
  NOR2X1 U39 ( .A(n3), .B(n15), .Y(n38) );
  NOR2X1 U40 ( .A(n3), .B(n16), .Y(n39) );
  NOR2X1 U41 ( .A(n4), .B(n9), .Y(n40) );
  NOR2X1 U42 ( .A(n4), .B(n10), .Y(n41) );
  NOR2X1 U43 ( .A(n4), .B(n11), .Y(n42) );
  NOR2X1 U44 ( .A(n4), .B(n12), .Y(n43) );
  NOR2X1 U45 ( .A(n4), .B(n13), .Y(n44) );
  NOR2X1 U46 ( .A(n4), .B(n14), .Y(n45) );
  NOR2X1 U47 ( .A(n4), .B(n15), .Y(n46) );
  NOR2X1 U48 ( .A(n4), .B(n16), .Y(n47) );
  NOR2X1 U49 ( .A(n5), .B(n9), .Y(n48) );
  NOR2X1 U50 ( .A(n5), .B(n10), .Y(n49) );
  NOR2X1 U51 ( .A(n5), .B(n11), .Y(n50) );
  NOR2X1 U52 ( .A(n5), .B(n12), .Y(n51) );
  NOR2X1 U53 ( .A(n5), .B(n13), .Y(n52) );
  NOR2X1 U54 ( .A(n5), .B(n14), .Y(n53) );
  NOR2X1 U55 ( .A(n5), .B(n15), .Y(n54) );
  NOR2X1 U56 ( .A(n5), .B(n16), .Y(n55) );
  NOR2X1 U57 ( .A(n6), .B(n9), .Y(n56) );
  NOR2X1 U58 ( .A(n6), .B(n10), .Y(n57) );
  NOR2X1 U59 ( .A(n6), .B(n11), .Y(n58) );
  NOR2X1 U60 ( .A(n6), .B(n12), .Y(n59) );
  NOR2X1 U61 ( .A(n6), .B(n13), .Y(n60) );
  NOR2X1 U62 ( .A(n6), .B(n14), .Y(n61) );
  NOR2X1 U63 ( .A(n6), .B(n15), .Y(n62) );
  NOR2X1 U64 ( .A(n6), .B(n16), .Y(n63) );
  NOR2X1 U65 ( .A(n7), .B(n9), .Y(n64) );
  NOR2X1 U66 ( .A(n7), .B(n10), .Y(n65) );
  NOR2X1 U67 ( .A(n7), .B(n11), .Y(n66) );
  NOR2X1 U68 ( .A(n7), .B(n12), .Y(n67) );
  NOR2X1 U69 ( .A(n7), .B(n13), .Y(n68) );
  NOR2X1 U70 ( .A(n7), .B(n14), .Y(n69) );
  NOR2X1 U71 ( .A(n7), .B(n15), .Y(n70) );
  NOR2X1 U72 ( .A(n7), .B(n16), .Y(n71) );
  NOR2X1 U73 ( .A(n8), .B(n9), .Y(n72) );
  NOR2X1 U74 ( .A(n8), .B(n10), .Y(n73) );
  NOR2X1 U75 ( .A(n8), .B(n11), .Y(n74) );
  NOR2X1 U76 ( .A(n8), .B(n12), .Y(n75) );
  NOR2X1 U77 ( .A(n8), .B(n13), .Y(n76) );
  NOR2X1 U78 ( .A(n8), .B(n14), .Y(n77) );
  NOR2X1 U79 ( .A(n8), .B(n15), .Y(n78) );
  NOR2X1 U80 ( .A(n8), .B(n16), .Y(n79) );
  HAX1 U81 ( .A(n18), .B(n25), .YC(n81), .YS(n80) );
  HAX1 U82 ( .A(n33), .B(n40), .YC(n83), .YS(n82) );
  FAX1 U83 ( .A(n19), .B(n26), .C(n81), .YC(n85), .YS(n84) );
  HAX1 U84 ( .A(n41), .B(n48), .YC(n87), .YS(n86) );
  FAX1 U85 ( .A(n20), .B(n34), .C(n27), .YC(n89), .YS(n88) );
  FAX1 U86 ( .A(n83), .B(n86), .C(n88), .YC(n91), .YS(n90) );
  HAX1 U87 ( .A(n49), .B(n56), .YC(n93), .YS(n92) );
  FAX1 U88 ( .A(n21), .B(n42), .C(n35), .YC(n95), .YS(n94) );
  FAX1 U89 ( .A(n28), .B(n87), .C(n92), .YC(n97), .YS(n96) );
  FAX1 U90 ( .A(n89), .B(n94), .C(n96), .YC(n99), .YS(n98) );
  HAX1 U91 ( .A(n57), .B(n64), .YC(n101), .YS(n100) );
  FAX1 U92 ( .A(n22), .B(n50), .C(n29), .YC(n103), .YS(n102) );
  FAX1 U93 ( .A(n36), .B(n43), .C(n93), .YC(n105), .YS(n104) );
  FAX1 U94 ( .A(n100), .B(n95), .C(n102), .YC(n107), .YS(n106) );
  FAX1 U95 ( .A(n97), .B(n104), .C(n106), .YC(n109), .YS(n108) );
  HAX1 U96 ( .A(n65), .B(n72), .YC(n111), .YS(n110) );
  FAX1 U97 ( .A(n23), .B(n58), .C(n30), .YC(n113), .YS(n112) );
  FAX1 U98 ( .A(n37), .B(n51), .C(n44), .YC(n115), .YS(n114) );
  FAX1 U99 ( .A(n101), .B(n110), .C(n103), .YC(n117), .YS(n116) );
  FAX1 U100 ( .A(n114), .B(n112), .C(n105), .YC(n119), .YS(n118) );
  FAX1 U101 ( .A(n107), .B(n116), .C(n118), .YC(n121), .YS(n120) );
  HAX1 U102 ( .A(n66), .B(n73), .YC(n123), .YS(n122) );
  FAX1 U103 ( .A(n52), .B(n59), .C(n31), .YC(n125), .YS(n124) );
  FAX1 U104 ( .A(n38), .B(n45), .C(n111), .YC(n127), .YS(n126) );
  FAX1 U105 ( .A(n122), .B(n113), .C(n115), .YC(n129), .YS(n128) );
  FAX1 U106 ( .A(n124), .B(n126), .C(n117), .YC(n131), .YS(n130) );
  FAX1 U107 ( .A(n128), .B(n119), .C(n130), .YC(n133), .YS(n132) );
  FAX1 U108 ( .A(n39), .B(n74), .C(n67), .YC(n135), .YS(n134) );
  FAX1 U109 ( .A(n60), .B(n53), .C(n46), .YC(n137), .YS(n136) );
  FAX1 U110 ( .A(n123), .B(n125), .C(n136), .YC(n139), .YS(n138) );
  FAX1 U111 ( .A(n134), .B(n127), .C(n129), .YC(n141), .YS(n140) );
  FAX1 U112 ( .A(n138), .B(n131), .C(n140), .YC(n143), .YS(n142) );
  FAX1 U113 ( .A(n47), .B(n75), .C(n68), .YC(n145), .YS(n144) );
  FAX1 U114 ( .A(n54), .B(n61), .C(n135), .YC(n147), .YS(n146) );
  FAX1 U115 ( .A(n137), .B(n144), .C(n139), .YC(n149), .YS(n148) );
  FAX1 U116 ( .A(n146), .B(n141), .C(n148), .YC(n151), .YS(n150) );
  FAX1 U117 ( .A(n55), .B(n76), .C(n69), .YC(n153), .YS(n152) );
  FAX1 U118 ( .A(n62), .B(n145), .C(n152), .YC(n155), .YS(n154) );
  FAX1 U119 ( .A(n147), .B(n154), .C(n149), .YC(n157), .YS(n156) );
  FAX1 U120 ( .A(n63), .B(n77), .C(n70), .YC(n159), .YS(n158) );
  FAX1 U121 ( .A(n153), .B(n158), .C(n155), .YC(n161), .YS(n160) );
  FAX1 U122 ( .A(n71), .B(n78), .C(n159), .YC(n163), .YS(n162) );
  HAX1 U123 ( .A(n24), .B(n17), .YC(n164), .YS(product[1]) );
  FAX1 U124 ( .A(n32), .B(n164), .C(n80), .YC(n165), .YS(product[2]) );
  FAX1 U125 ( .A(n82), .B(n165), .C(n84), .YC(n166), .YS(product[3]) );
  FAX1 U126 ( .A(n85), .B(n90), .C(n166), .YC(n167), .YS(product[4]) );
  FAX1 U127 ( .A(n91), .B(n98), .C(n167), .YC(n168), .YS(product[5]) );
  FAX1 U128 ( .A(n99), .B(n108), .C(n168), .YC(n169), .YS(product[6]) );
  FAX1 U129 ( .A(n109), .B(n120), .C(n169), .YC(n170), .YS(product[7]) );
  FAX1 U130 ( .A(n121), .B(n132), .C(n170), .YC(n171), .YS(product[8]) );
  FAX1 U131 ( .A(n133), .B(n142), .C(n171), .YC(n172), .YS(product[9]) );
  FAX1 U132 ( .A(n143), .B(n150), .C(n172), .YC(n173), .YS(product[10]) );
  FAX1 U133 ( .A(n151), .B(n156), .C(n173), .YC(n174), .YS(product[11]) );
  FAX1 U134 ( .A(n160), .B(n157), .C(n174), .YC(n175), .YS(product[12]) );
  FAX1 U135 ( .A(n162), .B(n161), .C(n175), .YC(n176), .YS(product[13]) );
  FAX1 U136 ( .A(n79), .B(n163), .C(n176), .YC(product[15]), .YS(product[14])
         );
  INVX2 U140 ( .A(b[0]), .Y(n9) );
  INVX2 U141 ( .A(b[1]), .Y(n10) );
  INVX2 U142 ( .A(b[2]), .Y(n11) );
  INVX2 U143 ( .A(b[3]), .Y(n12) );
  INVX2 U144 ( .A(b[4]), .Y(n13) );
  INVX2 U145 ( .A(b[5]), .Y(n14) );
  INVX2 U146 ( .A(b[6]), .Y(n15) );
  INVX2 U147 ( .A(b[7]), .Y(n16) );
  INVX2 U148 ( .A(a[0]), .Y(n1) );
  INVX2 U149 ( .A(a[1]), .Y(n2) );
  INVX2 U150 ( .A(a[2]), .Y(n3) );
  INVX2 U151 ( .A(a[3]), .Y(n4) );
  INVX2 U152 ( .A(a[4]), .Y(n5) );
  INVX2 U153 ( .A(a[5]), .Y(n6) );
  INVX2 U154 ( .A(a[6]), .Y(n7) );
  INVX2 U155 ( .A(a[7]), .Y(n8) );
endmodule


module alu_DW_mult_uns_4 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n15, n25, n26, n50, n60, n80, n85, n86, n101, n102, n117, n118, n133,
         n134, n149, n150, n160, n165, n176, n178, n187, n188, n189, n190,
         n191, n192, n193, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n221, n222, n223, n224, n225,
         n226, n227, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n940,
         n941, n942, n943, n944, n945, n946, n947;

  NAND2X1 OR_NOTi ( .A(n176), .B(n878), .Y(n236) );
  INVX1 U1 ( .A(n831), .Y(n176) );
  OAI21X1 AO21i ( .A(n165), .B(a[0]), .C(a[1]), .Y(n403) );
  INVX1 U12 ( .A(n846), .Y(n165) );
  NAND2X1 OR_NOTi1 ( .A(n160), .B(n876), .Y(n253) );
  INVX1 U13 ( .A(n831), .Y(n160) );
  OAI21X1 AO21i1 ( .A(n149), .B(n150), .C(a[3]), .Y(n421) );
  INVX1 U23 ( .A(n860), .Y(n150) );
  INVX1 U15 ( .A(n844), .Y(n149) );
  NAND2X1 OR_NOTi2 ( .A(n160), .B(n874), .Y(n270) );
  OAI21X1 AO21i2 ( .A(n133), .B(n134), .C(a[5]), .Y(n439) );
  INVX1 U25 ( .A(n858), .Y(n134) );
  INVX1 U18 ( .A(n842), .Y(n133) );
  NAND2X1 OR_NOTi3 ( .A(n160), .B(n872), .Y(n287) );
  OAI21X1 AO21i3 ( .A(n117), .B(n118), .C(a[7]), .Y(n457) );
  INVX1 U27 ( .A(n856), .Y(n118) );
  INVX1 U111 ( .A(n840), .Y(n117) );
  NAND2X1 OR_NOTi4 ( .A(n80), .B(n870), .Y(n304) );
  OAI21X1 AO21i4 ( .A(n101), .B(n102), .C(a[9]), .Y(n475) );
  INVX1 U29 ( .A(n854), .Y(n102) );
  INVX1 U114 ( .A(n838), .Y(n101) );
  NAND2X1 OR_NOTi5 ( .A(n80), .B(n868), .Y(n321) );
  OAI21X1 AO21i5 ( .A(n85), .B(n86), .C(a[11]), .Y(n493) );
  INVX1 U211 ( .A(n852), .Y(n86) );
  INVX1 U117 ( .A(n836), .Y(n85) );
  NAND2X1 OR_NOTi6 ( .A(n80), .B(n866), .Y(n338) );
  INVX1 U118 ( .A(n830), .Y(n80) );
  OAI21X1 AO21i6 ( .A(n50), .B(n60), .C(a[13]), .Y(n511) );
  INVX1 U213 ( .A(n850), .Y(n60) );
  INVX1 U120 ( .A(n834), .Y(n50) );
  NAND2X1 OR_NOTi7 ( .A(n176), .B(n864), .Y(n355) );
  OAI21X1 AO21i7 ( .A(n25), .B(n26), .C(a[15]), .Y(n529) );
  INVX1 U215 ( .A(n848), .Y(n26) );
  INVX1 U123 ( .A(n832), .Y(n25) );
  XOR2X1 U217 ( .A(n538), .B(n795), .Y(n15) );
  XOR2X1 U125 ( .A(n529), .B(n15), .Y(n798) );
  INVX2 U4 ( .A(a[0]), .Y(n195) );
  XOR2X1 U5 ( .A(a[0]), .B(a[1]), .Y(n212) );
  NAND2X1 U6 ( .A(n195), .B(n212), .Y(n204) );
  XNOR2X1 U7 ( .A(a[2]), .B(a[1]), .Y(n196) );
  XOR2X1 U8 ( .A(a[2]), .B(a[3]), .Y(n213) );
  NAND2X1 U9 ( .A(n213), .B(n196), .Y(n205) );
  XNOR2X1 U10 ( .A(a[4]), .B(a[3]), .Y(n197) );
  XOR2X1 U20 ( .A(a[4]), .B(a[5]), .Y(n214) );
  NAND2X1 U30 ( .A(n214), .B(n197), .Y(n206) );
  XNOR2X1 U38 ( .A(a[6]), .B(a[5]), .Y(n198) );
  XOR2X1 U39 ( .A(a[6]), .B(a[7]), .Y(n215) );
  NAND2X1 U40 ( .A(n215), .B(n198), .Y(n207) );
  XNOR2X1 U41 ( .A(a[8]), .B(a[7]), .Y(n199) );
  XOR2X1 U42 ( .A(a[8]), .B(a[9]), .Y(n216) );
  NAND2X1 U43 ( .A(n216), .B(n199), .Y(n208) );
  XNOR2X1 U44 ( .A(a[10]), .B(a[9]), .Y(n200) );
  XOR2X1 U45 ( .A(a[10]), .B(a[11]), .Y(n217) );
  NAND2X1 U46 ( .A(n217), .B(n200), .Y(n209) );
  XNOR2X1 U47 ( .A(a[12]), .B(a[11]), .Y(n201) );
  XOR2X1 U48 ( .A(a[12]), .B(a[13]), .Y(n218) );
  NAND2X1 U49 ( .A(n218), .B(n201), .Y(n210) );
  XNOR2X1 U50 ( .A(a[14]), .B(a[13]), .Y(n202) );
  XOR2X1 U51 ( .A(a[14]), .B(a[15]), .Y(n219) );
  NAND2X1 U52 ( .A(n219), .B(n202), .Y(n211) );
  INVX2 U53 ( .A(a[15]), .Y(n178) );
  INVX2 U54 ( .A(n879), .Y(n187) );
  INVX2 U55 ( .A(n877), .Y(n188) );
  INVX2 U56 ( .A(n875), .Y(n189) );
  INVX2 U57 ( .A(n873), .Y(n190) );
  INVX2 U58 ( .A(n871), .Y(n191) );
  INVX2 U59 ( .A(n869), .Y(n192) );
  INVX2 U60 ( .A(n867), .Y(n193) );
  XNOR2X1 U78 ( .A(n879), .B(n831), .Y(n237) );
  XNOR2X1 U79 ( .A(n879), .B(n221), .Y(n238) );
  XNOR2X1 U80 ( .A(n879), .B(n222), .Y(n239) );
  XNOR2X1 U81 ( .A(n879), .B(n223), .Y(n240) );
  XNOR2X1 U82 ( .A(n879), .B(n224), .Y(n241) );
  XNOR2X1 U83 ( .A(n879), .B(n225), .Y(n242) );
  XNOR2X1 U84 ( .A(n879), .B(n226), .Y(n243) );
  XNOR2X1 U85 ( .A(n879), .B(n227), .Y(n244) );
  XNOR2X1 U86 ( .A(n878), .B(b[8]), .Y(n245) );
  XNOR2X1 U87 ( .A(n878), .B(b[9]), .Y(n246) );
  XNOR2X1 U88 ( .A(n878), .B(b[10]), .Y(n247) );
  XNOR2X1 U89 ( .A(n878), .B(b[11]), .Y(n248) );
  XNOR2X1 U90 ( .A(n878), .B(b[12]), .Y(n249) );
  XNOR2X1 U91 ( .A(n878), .B(b[13]), .Y(n250) );
  XNOR2X1 U92 ( .A(n878), .B(b[14]), .Y(n251) );
  XNOR2X1 U93 ( .A(n878), .B(b[15]), .Y(n252) );
  OAI22X1 U94 ( .A(n863), .B(n238), .C(n237), .D(n847), .Y(n387) );
  OAI22X1 U95 ( .A(n863), .B(n239), .C(n238), .D(n847), .Y(n388) );
  OAI22X1 U96 ( .A(n863), .B(n240), .C(n239), .D(n847), .Y(n389) );
  OAI22X1 U97 ( .A(n863), .B(n241), .C(n240), .D(n847), .Y(n390) );
  OAI22X1 U98 ( .A(n863), .B(n242), .C(n241), .D(n847), .Y(n391) );
  OAI22X1 U99 ( .A(n863), .B(n243), .C(n242), .D(n847), .Y(n392) );
  OAI22X1 U100 ( .A(n863), .B(n244), .C(n243), .D(n847), .Y(n393) );
  OAI22X1 U101 ( .A(n863), .B(n245), .C(n244), .D(n847), .Y(n394) );
  OAI22X1 U102 ( .A(n863), .B(n246), .C(n245), .D(n847), .Y(n395) );
  OAI22X1 U103 ( .A(n862), .B(n247), .C(n246), .D(n846), .Y(n396) );
  OAI22X1 U104 ( .A(n862), .B(n248), .C(n247), .D(n846), .Y(n397) );
  OAI22X1 U105 ( .A(n862), .B(n249), .C(n248), .D(n846), .Y(n398) );
  OAI22X1 U106 ( .A(n862), .B(n250), .C(n249), .D(n846), .Y(n399) );
  OAI22X1 U107 ( .A(n862), .B(n251), .C(n250), .D(n846), .Y(n400) );
  OAI22X1 U108 ( .A(n862), .B(n252), .C(n251), .D(n846), .Y(n401) );
  OAI22X1 U109 ( .A(n862), .B(n187), .C(n252), .D(n846), .Y(n402) );
  OAI22X1 U127 ( .A(n862), .B(n236), .C(n187), .D(n846), .Y(n539) );
  XNOR2X1 U128 ( .A(n877), .B(n831), .Y(n254) );
  XNOR2X1 U129 ( .A(n877), .B(n221), .Y(n255) );
  XNOR2X1 U130 ( .A(n877), .B(n222), .Y(n256) );
  XNOR2X1 U131 ( .A(n877), .B(n223), .Y(n257) );
  XNOR2X1 U132 ( .A(n877), .B(n224), .Y(n258) );
  XNOR2X1 U133 ( .A(n877), .B(n225), .Y(n259) );
  XNOR2X1 U134 ( .A(n877), .B(n226), .Y(n260) );
  XNOR2X1 U135 ( .A(n877), .B(n227), .Y(n261) );
  XNOR2X1 U136 ( .A(n876), .B(b[8]), .Y(n262) );
  XNOR2X1 U137 ( .A(n876), .B(b[9]), .Y(n263) );
  XNOR2X1 U138 ( .A(n876), .B(b[10]), .Y(n264) );
  XNOR2X1 U139 ( .A(n876), .B(b[11]), .Y(n265) );
  XNOR2X1 U140 ( .A(n876), .B(b[12]), .Y(n266) );
  XNOR2X1 U141 ( .A(n876), .B(b[13]), .Y(n267) );
  XNOR2X1 U142 ( .A(n876), .B(b[14]), .Y(n268) );
  XNOR2X1 U143 ( .A(n876), .B(b[15]), .Y(n269) );
  OAI22X1 U144 ( .A(n255), .B(n861), .C(n254), .D(n845), .Y(n405) );
  OAI22X1 U145 ( .A(n256), .B(n861), .C(n255), .D(n845), .Y(n406) );
  OAI22X1 U146 ( .A(n257), .B(n861), .C(n256), .D(n845), .Y(n407) );
  OAI22X1 U147 ( .A(n258), .B(n861), .C(n257), .D(n845), .Y(n408) );
  OAI22X1 U148 ( .A(n259), .B(n861), .C(n258), .D(n845), .Y(n409) );
  OAI22X1 U149 ( .A(n260), .B(n861), .C(n259), .D(n845), .Y(n410) );
  OAI22X1 U150 ( .A(n261), .B(n861), .C(n260), .D(n845), .Y(n411) );
  OAI22X1 U151 ( .A(n262), .B(n861), .C(n261), .D(n845), .Y(n412) );
  OAI22X1 U152 ( .A(n263), .B(n861), .C(n262), .D(n845), .Y(n413) );
  OAI22X1 U153 ( .A(n264), .B(n860), .C(n263), .D(n844), .Y(n414) );
  OAI22X1 U154 ( .A(n265), .B(n860), .C(n264), .D(n844), .Y(n415) );
  OAI22X1 U155 ( .A(n266), .B(n860), .C(n265), .D(n844), .Y(n416) );
  OAI22X1 U156 ( .A(n267), .B(n860), .C(n266), .D(n844), .Y(n417) );
  OAI22X1 U157 ( .A(n268), .B(n860), .C(n267), .D(n844), .Y(n418) );
  OAI22X1 U158 ( .A(n269), .B(n860), .C(n268), .D(n844), .Y(n419) );
  OAI22X1 U159 ( .A(n188), .B(n860), .C(n269), .D(n844), .Y(n420) );
  OAI22X1 U160 ( .A(n860), .B(n253), .C(n188), .D(n844), .Y(n540) );
  XNOR2X1 U161 ( .A(n875), .B(n831), .Y(n271) );
  XNOR2X1 U162 ( .A(n875), .B(n221), .Y(n272) );
  XNOR2X1 U163 ( .A(n875), .B(n222), .Y(n273) );
  XNOR2X1 U164 ( .A(n875), .B(n223), .Y(n274) );
  XNOR2X1 U165 ( .A(n875), .B(n224), .Y(n275) );
  XNOR2X1 U166 ( .A(n875), .B(n225), .Y(n276) );
  XNOR2X1 U167 ( .A(n875), .B(n226), .Y(n277) );
  XNOR2X1 U168 ( .A(n875), .B(n227), .Y(n278) );
  XNOR2X1 U169 ( .A(n874), .B(b[8]), .Y(n279) );
  XNOR2X1 U170 ( .A(n874), .B(b[9]), .Y(n280) );
  XNOR2X1 U171 ( .A(n874), .B(b[10]), .Y(n281) );
  XNOR2X1 U172 ( .A(n874), .B(b[11]), .Y(n282) );
  XNOR2X1 U173 ( .A(n874), .B(b[12]), .Y(n283) );
  XNOR2X1 U174 ( .A(n874), .B(b[13]), .Y(n284) );
  XNOR2X1 U175 ( .A(n874), .B(b[14]), .Y(n285) );
  XNOR2X1 U176 ( .A(n874), .B(b[15]), .Y(n286) );
  OAI22X1 U177 ( .A(n272), .B(n859), .C(n271), .D(n843), .Y(n423) );
  OAI22X1 U178 ( .A(n273), .B(n859), .C(n272), .D(n843), .Y(n424) );
  OAI22X1 U179 ( .A(n274), .B(n859), .C(n273), .D(n843), .Y(n425) );
  OAI22X1 U180 ( .A(n275), .B(n859), .C(n274), .D(n843), .Y(n426) );
  OAI22X1 U181 ( .A(n276), .B(n859), .C(n275), .D(n843), .Y(n427) );
  OAI22X1 U182 ( .A(n277), .B(n859), .C(n276), .D(n843), .Y(n428) );
  OAI22X1 U183 ( .A(n278), .B(n859), .C(n277), .D(n843), .Y(n429) );
  OAI22X1 U184 ( .A(n279), .B(n859), .C(n278), .D(n843), .Y(n430) );
  OAI22X1 U185 ( .A(n280), .B(n859), .C(n279), .D(n843), .Y(n431) );
  OAI22X1 U186 ( .A(n281), .B(n858), .C(n280), .D(n842), .Y(n432) );
  OAI22X1 U187 ( .A(n282), .B(n858), .C(n281), .D(n842), .Y(n433) );
  OAI22X1 U188 ( .A(n283), .B(n858), .C(n282), .D(n842), .Y(n434) );
  OAI22X1 U189 ( .A(n284), .B(n858), .C(n283), .D(n842), .Y(n435) );
  OAI22X1 U190 ( .A(n285), .B(n858), .C(n284), .D(n842), .Y(n436) );
  OAI22X1 U191 ( .A(n286), .B(n858), .C(n285), .D(n842), .Y(n437) );
  OAI22X1 U192 ( .A(n189), .B(n858), .C(n286), .D(n842), .Y(n438) );
  OAI22X1 U193 ( .A(n858), .B(n270), .C(n189), .D(n842), .Y(n541) );
  XNOR2X1 U194 ( .A(n873), .B(n831), .Y(n288) );
  XNOR2X1 U195 ( .A(n873), .B(n221), .Y(n289) );
  XNOR2X1 U196 ( .A(n873), .B(n222), .Y(n290) );
  XNOR2X1 U197 ( .A(n873), .B(n223), .Y(n291) );
  XNOR2X1 U198 ( .A(n873), .B(n224), .Y(n292) );
  XNOR2X1 U199 ( .A(n873), .B(n225), .Y(n293) );
  XNOR2X1 U200 ( .A(n873), .B(n226), .Y(n294) );
  XNOR2X1 U201 ( .A(n873), .B(n227), .Y(n295) );
  XNOR2X1 U202 ( .A(n872), .B(b[8]), .Y(n296) );
  XNOR2X1 U203 ( .A(n872), .B(b[9]), .Y(n297) );
  XNOR2X1 U204 ( .A(n872), .B(b[10]), .Y(n298) );
  XNOR2X1 U205 ( .A(n872), .B(b[11]), .Y(n299) );
  XNOR2X1 U206 ( .A(n872), .B(b[12]), .Y(n300) );
  XNOR2X1 U207 ( .A(n872), .B(b[13]), .Y(n301) );
  XNOR2X1 U208 ( .A(n872), .B(b[14]), .Y(n302) );
  XNOR2X1 U209 ( .A(n872), .B(b[15]), .Y(n303) );
  OAI22X1 U218 ( .A(n289), .B(n857), .C(n288), .D(n841), .Y(n441) );
  OAI22X1 U219 ( .A(n290), .B(n857), .C(n289), .D(n841), .Y(n442) );
  OAI22X1 U220 ( .A(n291), .B(n857), .C(n290), .D(n841), .Y(n443) );
  OAI22X1 U221 ( .A(n292), .B(n857), .C(n291), .D(n841), .Y(n444) );
  OAI22X1 U222 ( .A(n293), .B(n857), .C(n292), .D(n841), .Y(n445) );
  OAI22X1 U223 ( .A(n294), .B(n857), .C(n293), .D(n841), .Y(n446) );
  OAI22X1 U224 ( .A(n295), .B(n857), .C(n294), .D(n841), .Y(n447) );
  OAI22X1 U225 ( .A(n296), .B(n857), .C(n295), .D(n841), .Y(n448) );
  OAI22X1 U226 ( .A(n297), .B(n857), .C(n296), .D(n841), .Y(n449) );
  OAI22X1 U227 ( .A(n298), .B(n856), .C(n297), .D(n840), .Y(n450) );
  OAI22X1 U228 ( .A(n299), .B(n856), .C(n298), .D(n840), .Y(n451) );
  OAI22X1 U229 ( .A(n300), .B(n856), .C(n299), .D(n840), .Y(n452) );
  OAI22X1 U230 ( .A(n301), .B(n856), .C(n300), .D(n840), .Y(n453) );
  OAI22X1 U231 ( .A(n302), .B(n856), .C(n301), .D(n840), .Y(n454) );
  OAI22X1 U232 ( .A(n303), .B(n856), .C(n302), .D(n840), .Y(n455) );
  OAI22X1 U233 ( .A(n190), .B(n856), .C(n303), .D(n840), .Y(n456) );
  OAI22X1 U234 ( .A(n856), .B(n287), .C(n190), .D(n840), .Y(n542) );
  XNOR2X1 U235 ( .A(n871), .B(n831), .Y(n305) );
  XNOR2X1 U236 ( .A(n871), .B(n221), .Y(n306) );
  XNOR2X1 U237 ( .A(n871), .B(n222), .Y(n307) );
  XNOR2X1 U238 ( .A(n871), .B(n223), .Y(n308) );
  XNOR2X1 U239 ( .A(n871), .B(n224), .Y(n309) );
  XNOR2X1 U240 ( .A(n871), .B(n225), .Y(n310) );
  XNOR2X1 U241 ( .A(n871), .B(n226), .Y(n311) );
  XNOR2X1 U242 ( .A(n871), .B(n227), .Y(n312) );
  XNOR2X1 U243 ( .A(n870), .B(b[8]), .Y(n313) );
  XNOR2X1 U244 ( .A(n870), .B(b[9]), .Y(n314) );
  XNOR2X1 U245 ( .A(n870), .B(b[10]), .Y(n315) );
  XNOR2X1 U246 ( .A(n870), .B(b[11]), .Y(n316) );
  XNOR2X1 U247 ( .A(n870), .B(b[12]), .Y(n317) );
  XNOR2X1 U248 ( .A(n870), .B(b[13]), .Y(n318) );
  XNOR2X1 U249 ( .A(n870), .B(b[14]), .Y(n319) );
  XNOR2X1 U250 ( .A(n870), .B(b[15]), .Y(n320) );
  OAI22X1 U251 ( .A(n306), .B(n855), .C(n305), .D(n839), .Y(n459) );
  OAI22X1 U252 ( .A(n307), .B(n855), .C(n306), .D(n839), .Y(n460) );
  OAI22X1 U253 ( .A(n308), .B(n855), .C(n307), .D(n839), .Y(n461) );
  OAI22X1 U254 ( .A(n309), .B(n855), .C(n308), .D(n839), .Y(n462) );
  OAI22X1 U255 ( .A(n310), .B(n855), .C(n309), .D(n839), .Y(n463) );
  OAI22X1 U256 ( .A(n311), .B(n855), .C(n310), .D(n839), .Y(n464) );
  OAI22X1 U257 ( .A(n312), .B(n855), .C(n311), .D(n839), .Y(n465) );
  OAI22X1 U258 ( .A(n313), .B(n855), .C(n312), .D(n839), .Y(n466) );
  OAI22X1 U259 ( .A(n314), .B(n855), .C(n313), .D(n839), .Y(n467) );
  OAI22X1 U260 ( .A(n315), .B(n854), .C(n314), .D(n838), .Y(n468) );
  OAI22X1 U261 ( .A(n316), .B(n854), .C(n315), .D(n838), .Y(n469) );
  OAI22X1 U262 ( .A(n317), .B(n854), .C(n316), .D(n838), .Y(n470) );
  OAI22X1 U263 ( .A(n318), .B(n854), .C(n317), .D(n838), .Y(n471) );
  OAI22X1 U264 ( .A(n319), .B(n854), .C(n318), .D(n838), .Y(n472) );
  OAI22X1 U265 ( .A(n320), .B(n854), .C(n319), .D(n838), .Y(n473) );
  OAI22X1 U266 ( .A(n191), .B(n854), .C(n320), .D(n838), .Y(n474) );
  OAI22X1 U267 ( .A(n854), .B(n304), .C(n191), .D(n838), .Y(n543) );
  XNOR2X1 U268 ( .A(n869), .B(n831), .Y(n322) );
  XNOR2X1 U269 ( .A(n869), .B(n221), .Y(n323) );
  XNOR2X1 U270 ( .A(n869), .B(n222), .Y(n324) );
  XNOR2X1 U271 ( .A(n869), .B(n223), .Y(n325) );
  XNOR2X1 U272 ( .A(n869), .B(n224), .Y(n326) );
  XNOR2X1 U273 ( .A(n869), .B(n225), .Y(n327) );
  XNOR2X1 U274 ( .A(n869), .B(n226), .Y(n328) );
  XNOR2X1 U275 ( .A(n869), .B(n227), .Y(n329) );
  XNOR2X1 U276 ( .A(n868), .B(b[8]), .Y(n330) );
  XNOR2X1 U277 ( .A(n868), .B(b[9]), .Y(n331) );
  XNOR2X1 U278 ( .A(n868), .B(b[10]), .Y(n332) );
  XNOR2X1 U279 ( .A(n868), .B(b[11]), .Y(n333) );
  XNOR2X1 U280 ( .A(n868), .B(b[12]), .Y(n334) );
  XNOR2X1 U281 ( .A(n868), .B(b[13]), .Y(n335) );
  XNOR2X1 U282 ( .A(n868), .B(b[14]), .Y(n336) );
  XNOR2X1 U283 ( .A(n868), .B(b[15]), .Y(n337) );
  OAI22X1 U284 ( .A(n323), .B(n853), .C(n322), .D(n837), .Y(n477) );
  OAI22X1 U285 ( .A(n324), .B(n853), .C(n323), .D(n837), .Y(n478) );
  OAI22X1 U286 ( .A(n325), .B(n853), .C(n324), .D(n837), .Y(n479) );
  OAI22X1 U287 ( .A(n326), .B(n853), .C(n325), .D(n837), .Y(n480) );
  OAI22X1 U288 ( .A(n327), .B(n853), .C(n326), .D(n837), .Y(n481) );
  OAI22X1 U289 ( .A(n328), .B(n853), .C(n327), .D(n837), .Y(n482) );
  OAI22X1 U290 ( .A(n329), .B(n853), .C(n328), .D(n837), .Y(n483) );
  OAI22X1 U291 ( .A(n330), .B(n853), .C(n329), .D(n837), .Y(n484) );
  OAI22X1 U292 ( .A(n331), .B(n853), .C(n330), .D(n837), .Y(n485) );
  OAI22X1 U293 ( .A(n332), .B(n852), .C(n331), .D(n836), .Y(n486) );
  OAI22X1 U294 ( .A(n333), .B(n852), .C(n332), .D(n836), .Y(n487) );
  OAI22X1 U295 ( .A(n334), .B(n852), .C(n333), .D(n836), .Y(n488) );
  OAI22X1 U296 ( .A(n335), .B(n852), .C(n334), .D(n836), .Y(n489) );
  OAI22X1 U297 ( .A(n336), .B(n852), .C(n335), .D(n836), .Y(n490) );
  OAI22X1 U298 ( .A(n337), .B(n852), .C(n336), .D(n836), .Y(n491) );
  OAI22X1 U299 ( .A(n192), .B(n852), .C(n337), .D(n836), .Y(n492) );
  OAI22X1 U300 ( .A(n852), .B(n321), .C(n192), .D(n836), .Y(n544) );
  XNOR2X1 U301 ( .A(n867), .B(n831), .Y(n339) );
  XNOR2X1 U302 ( .A(n867), .B(n221), .Y(n340) );
  XNOR2X1 U303 ( .A(n867), .B(n222), .Y(n341) );
  XNOR2X1 U304 ( .A(n867), .B(n223), .Y(n342) );
  XNOR2X1 U305 ( .A(n867), .B(n224), .Y(n343) );
  XNOR2X1 U306 ( .A(n867), .B(n225), .Y(n344) );
  XNOR2X1 U307 ( .A(n867), .B(n226), .Y(n345) );
  XNOR2X1 U308 ( .A(n867), .B(n227), .Y(n346) );
  XNOR2X1 U309 ( .A(n866), .B(b[8]), .Y(n347) );
  XNOR2X1 U310 ( .A(n866), .B(b[9]), .Y(n348) );
  XNOR2X1 U311 ( .A(n866), .B(b[10]), .Y(n349) );
  XNOR2X1 U312 ( .A(n866), .B(b[11]), .Y(n350) );
  XNOR2X1 U313 ( .A(n866), .B(b[12]), .Y(n351) );
  XNOR2X1 U314 ( .A(n866), .B(b[13]), .Y(n352) );
  XNOR2X1 U315 ( .A(n866), .B(b[14]), .Y(n353) );
  XNOR2X1 U316 ( .A(n866), .B(b[15]), .Y(n354) );
  OAI22X1 U317 ( .A(n340), .B(n851), .C(n339), .D(n835), .Y(n495) );
  OAI22X1 U318 ( .A(n341), .B(n851), .C(n340), .D(n835), .Y(n496) );
  OAI22X1 U319 ( .A(n342), .B(n851), .C(n341), .D(n835), .Y(n497) );
  OAI22X1 U320 ( .A(n343), .B(n851), .C(n342), .D(n835), .Y(n498) );
  OAI22X1 U321 ( .A(n344), .B(n851), .C(n343), .D(n835), .Y(n499) );
  OAI22X1 U322 ( .A(n345), .B(n851), .C(n344), .D(n835), .Y(n500) );
  OAI22X1 U323 ( .A(n346), .B(n851), .C(n345), .D(n835), .Y(n501) );
  OAI22X1 U324 ( .A(n347), .B(n851), .C(n346), .D(n835), .Y(n502) );
  OAI22X1 U325 ( .A(n348), .B(n851), .C(n347), .D(n835), .Y(n503) );
  OAI22X1 U326 ( .A(n349), .B(n850), .C(n348), .D(n834), .Y(n504) );
  OAI22X1 U327 ( .A(n350), .B(n850), .C(n349), .D(n834), .Y(n505) );
  OAI22X1 U328 ( .A(n351), .B(n850), .C(n350), .D(n834), .Y(n506) );
  OAI22X1 U329 ( .A(n352), .B(n850), .C(n351), .D(n834), .Y(n507) );
  OAI22X1 U330 ( .A(n353), .B(n850), .C(n352), .D(n834), .Y(n508) );
  OAI22X1 U331 ( .A(n354), .B(n850), .C(n353), .D(n834), .Y(n509) );
  OAI22X1 U332 ( .A(n193), .B(n850), .C(n354), .D(n834), .Y(n510) );
  OAI22X1 U333 ( .A(n850), .B(n338), .C(n193), .D(n834), .Y(n545) );
  XNOR2X1 U334 ( .A(n865), .B(n831), .Y(n356) );
  XNOR2X1 U335 ( .A(n865), .B(n221), .Y(n357) );
  XNOR2X1 U336 ( .A(n865), .B(n222), .Y(n358) );
  XNOR2X1 U337 ( .A(n865), .B(n223), .Y(n359) );
  XNOR2X1 U338 ( .A(n865), .B(n224), .Y(n360) );
  XNOR2X1 U339 ( .A(n865), .B(n225), .Y(n361) );
  XNOR2X1 U340 ( .A(n865), .B(n226), .Y(n362) );
  XNOR2X1 U341 ( .A(n865), .B(n227), .Y(n363) );
  XNOR2X1 U342 ( .A(n864), .B(b[8]), .Y(n364) );
  XNOR2X1 U343 ( .A(n864), .B(b[9]), .Y(n365) );
  XNOR2X1 U344 ( .A(n864), .B(b[10]), .Y(n366) );
  XNOR2X1 U345 ( .A(n864), .B(b[11]), .Y(n367) );
  XNOR2X1 U346 ( .A(n864), .B(b[12]), .Y(n368) );
  XNOR2X1 U347 ( .A(n864), .B(b[13]), .Y(n369) );
  XNOR2X1 U348 ( .A(n864), .B(b[14]), .Y(n370) );
  XNOR2X1 U349 ( .A(n864), .B(b[15]), .Y(n371) );
  OAI22X1 U350 ( .A(n357), .B(n849), .C(n356), .D(n833), .Y(n513) );
  OAI22X1 U351 ( .A(n358), .B(n849), .C(n357), .D(n833), .Y(n514) );
  OAI22X1 U352 ( .A(n359), .B(n849), .C(n358), .D(n833), .Y(n515) );
  OAI22X1 U353 ( .A(n360), .B(n849), .C(n359), .D(n833), .Y(n516) );
  OAI22X1 U354 ( .A(n361), .B(n849), .C(n360), .D(n833), .Y(n517) );
  OAI22X1 U355 ( .A(n362), .B(n849), .C(n361), .D(n833), .Y(n518) );
  OAI22X1 U356 ( .A(n363), .B(n849), .C(n362), .D(n833), .Y(n519) );
  OAI22X1 U357 ( .A(n364), .B(n849), .C(n363), .D(n833), .Y(n520) );
  OAI22X1 U358 ( .A(n365), .B(n849), .C(n364), .D(n833), .Y(n521) );
  OAI22X1 U359 ( .A(n366), .B(n848), .C(n365), .D(n832), .Y(n522) );
  OAI22X1 U360 ( .A(n367), .B(n848), .C(n366), .D(n832), .Y(n523) );
  OAI22X1 U361 ( .A(n368), .B(n848), .C(n367), .D(n832), .Y(n524) );
  OAI22X1 U362 ( .A(n369), .B(n848), .C(n368), .D(n832), .Y(n525) );
  OAI22X1 U363 ( .A(n370), .B(n848), .C(n369), .D(n832), .Y(n526) );
  OAI22X1 U364 ( .A(n371), .B(n848), .C(n370), .D(n832), .Y(n527) );
  OAI22X1 U365 ( .A(n178), .B(n848), .C(n371), .D(n832), .Y(n528) );
  OAI22X1 U366 ( .A(n848), .B(n355), .C(n178), .D(n832), .Y(n546) );
  INVX2 U367 ( .A(n221), .Y(n372) );
  INVX2 U368 ( .A(n222), .Y(n373) );
  INVX2 U369 ( .A(n223), .Y(n374) );
  INVX2 U370 ( .A(n224), .Y(n375) );
  INVX2 U371 ( .A(n225), .Y(n376) );
  INVX2 U372 ( .A(n226), .Y(n377) );
  INVX2 U373 ( .A(n227), .Y(n378) );
  INVX2 U374 ( .A(b[8]), .Y(n379) );
  INVX2 U375 ( .A(b[9]), .Y(n380) );
  INVX2 U376 ( .A(b[10]), .Y(n381) );
  INVX2 U377 ( .A(b[11]), .Y(n382) );
  INVX2 U378 ( .A(b[12]), .Y(n383) );
  INVX2 U379 ( .A(b[13]), .Y(n384) );
  INVX2 U380 ( .A(b[14]), .Y(n385) );
  INVX2 U381 ( .A(b[15]), .Y(n386) );
  NOR2X1 U382 ( .A(n372), .B(n203), .Y(n675) );
  NOR2X1 U383 ( .A(n373), .B(n203), .Y(n531) );
  NOR2X1 U384 ( .A(n374), .B(n203), .Y(n532) );
  NOR2X1 U385 ( .A(n375), .B(n203), .Y(n705) );
  NOR2X1 U386 ( .A(n376), .B(n203), .Y(n533) );
  NOR2X1 U387 ( .A(n377), .B(n203), .Y(n731) );
  NOR2X1 U388 ( .A(n378), .B(n203), .Y(n534) );
  NOR2X1 U389 ( .A(n379), .B(n203), .Y(n753) );
  NOR2X1 U390 ( .A(n380), .B(n203), .Y(n535) );
  NOR2X1 U391 ( .A(n381), .B(n203), .Y(n771) );
  NOR2X1 U392 ( .A(n382), .B(n203), .Y(n536) );
  NOR2X1 U393 ( .A(n383), .B(n203), .Y(n785) );
  NOR2X1 U394 ( .A(n384), .B(n203), .Y(n537) );
  NOR2X1 U395 ( .A(n385), .B(n203), .Y(n795) );
  NOR2X1 U396 ( .A(n386), .B(n203), .Y(n538) );
  HAX1 U397 ( .A(n389), .B(n405), .YC(n548), .YS(n547) );
  FAX1 U398 ( .A(n390), .B(n406), .C(n548), .YC(n550), .YS(n549) );
  HAX1 U399 ( .A(n391), .B(n541), .YC(n552), .YS(n551) );
  FAX1 U400 ( .A(n407), .B(n423), .C(n551), .YC(n554), .YS(n553) );
  FAX1 U401 ( .A(n392), .B(n424), .C(n408), .YC(n556), .YS(n555) );
  FAX1 U402 ( .A(n552), .B(n943), .C(n555), .YC(n558), .YS(n557) );
  HAX1 U403 ( .A(n393), .B(n542), .YC(n560), .YS(n559) );
  FAX1 U404 ( .A(n409), .B(n441), .C(n425), .YC(n562), .YS(n561) );
  FAX1 U405 ( .A(n559), .B(n556), .C(n561), .YC(n564), .YS(n563) );
  FAX1 U406 ( .A(n394), .B(n426), .C(n442), .YC(n566), .YS(n565) );
  FAX1 U407 ( .A(n410), .B(n560), .C(n946), .YC(n568), .YS(n567) );
  FAX1 U408 ( .A(n562), .B(n565), .C(n567), .YC(n570), .YS(n569) );
  HAX1 U409 ( .A(n395), .B(n543), .YC(n572), .YS(n571) );
  FAX1 U410 ( .A(n443), .B(n459), .C(n427), .YC(n574), .YS(n573) );
  FAX1 U411 ( .A(n411), .B(n571), .C(n566), .YC(n576), .YS(n575) );
  FAX1 U412 ( .A(n573), .B(n568), .C(n575), .YC(n578), .YS(n577) );
  FAX1 U413 ( .A(n396), .B(n412), .C(n428), .YC(n580), .YS(n579) );
  FAX1 U414 ( .A(n444), .B(n460), .C(n572), .YC(n582), .YS(n581) );
  FAX1 U415 ( .A(n941), .B(n574), .C(n579), .YC(n584), .YS(n583) );
  FAX1 U416 ( .A(n581), .B(n576), .C(n583), .YC(n586), .YS(n585) );
  HAX1 U417 ( .A(n397), .B(n544), .YC(n588), .YS(n587) );
  FAX1 U418 ( .A(n445), .B(n477), .C(n413), .YC(n590), .YS(n589) );
  FAX1 U419 ( .A(n429), .B(n461), .C(n587), .YC(n592), .YS(n591) );
  FAX1 U420 ( .A(n580), .B(n589), .C(n582), .YC(n594), .YS(n593) );
  FAX1 U421 ( .A(n591), .B(n584), .C(n593), .YC(n596), .YS(n595) );
  FAX1 U422 ( .A(n398), .B(n414), .C(n478), .YC(n598), .YS(n597) );
  FAX1 U423 ( .A(n430), .B(n462), .C(n446), .YC(n600), .YS(n599) );
  FAX1 U424 ( .A(n588), .B(n942), .C(n590), .YC(n602), .YS(n601) );
  FAX1 U425 ( .A(n597), .B(n599), .C(n592), .YC(n604), .YS(n603) );
  FAX1 U426 ( .A(n601), .B(n594), .C(n603), .YC(n606), .YS(n605) );
  HAX1 U427 ( .A(n399), .B(n545), .YC(n608), .YS(n607) );
  FAX1 U428 ( .A(n463), .B(n415), .C(n431), .YC(n610), .YS(n609) );
  FAX1 U429 ( .A(n447), .B(n495), .C(n479), .YC(n612), .YS(n611) );
  FAX1 U430 ( .A(n607), .B(n598), .C(n600), .YC(n614), .YS(n613) );
  FAX1 U431 ( .A(n611), .B(n609), .C(n602), .YC(n616), .YS(n615) );
  FAX1 U432 ( .A(n613), .B(n604), .C(n615), .YC(n618), .YS(n617) );
  FAX1 U433 ( .A(n400), .B(n416), .C(n432), .YC(n620), .YS(n619) );
  FAX1 U434 ( .A(n448), .B(n496), .C(n480), .YC(n622), .YS(n621) );
  FAX1 U435 ( .A(n464), .B(n608), .C(n945), .YC(n624), .YS(n623) );
  FAX1 U436 ( .A(n610), .B(n612), .C(n619), .YC(n626), .YS(n625) );
  FAX1 U437 ( .A(n621), .B(n623), .C(n614), .YC(n628), .YS(n627) );
  FAX1 U438 ( .A(n625), .B(n616), .C(n627), .YC(n630), .YS(n629) );
  HAX1 U439 ( .A(n401), .B(n546), .YC(n632), .YS(n631) );
  FAX1 U440 ( .A(n465), .B(n513), .C(n497), .YC(n634), .YS(n633) );
  FAX1 U441 ( .A(n417), .B(n481), .C(n449), .YC(n636), .YS(n635) );
  FAX1 U442 ( .A(n433), .B(n631), .C(n620), .YC(n638), .YS(n637) );
  FAX1 U443 ( .A(n622), .B(n635), .C(n633), .YC(n640), .YS(n639) );
  FAX1 U444 ( .A(n624), .B(n626), .C(n637), .YC(n642), .YS(n641) );
  FAX1 U445 ( .A(n639), .B(n628), .C(n641), .YC(n644), .YS(n643) );
  FAX1 U446 ( .A(n402), .B(n418), .C(n947), .YC(n646), .YS(n645) );
  FAX1 U447 ( .A(n434), .B(n514), .C(n498), .YC(n648), .YS(n647) );
  FAX1 U448 ( .A(n450), .B(n482), .C(n466), .YC(n650), .YS(n649) );
  FAX1 U449 ( .A(n632), .B(n634), .C(n636), .YC(n652), .YS(n651) );
  FAX1 U450 ( .A(n645), .B(n649), .C(n647), .YC(n654), .YS(n653) );
  FAX1 U451 ( .A(n638), .B(n640), .C(n651), .YC(n656), .YS(n655) );
  FAX1 U452 ( .A(n653), .B(n642), .C(n655), .YC(n658), .YS(n657) );
  INVX2 U453 ( .A(n675), .Y(n659) );
  FAX1 U454 ( .A(n659), .B(n499), .C(n451), .YC(n661), .YS(n660) );
  FAX1 U455 ( .A(n467), .B(n483), .C(n515), .YC(n663), .YS(n662) );
  FAX1 U456 ( .A(n419), .B(n435), .C(n403), .YC(n665), .YS(n664) );
  FAX1 U457 ( .A(n646), .B(n648), .C(n650), .YC(n667), .YS(n666) );
  FAX1 U458 ( .A(n660), .B(n662), .C(n664), .YC(n669), .YS(n668) );
  FAX1 U459 ( .A(n652), .B(n654), .C(n666), .YC(n671), .YS(n670) );
  FAX1 U460 ( .A(n668), .B(n656), .C(n670), .YC(n673), .YS(n672) );
  FAX1 U462 ( .A(n531), .B(n659), .C(n420), .YC(n677), .YS(n676) );
  FAX1 U463 ( .A(n436), .B(n516), .C(n452), .YC(n679), .YS(n678) );
  FAX1 U464 ( .A(n468), .B(n500), .C(n484), .YC(n681), .YS(n680) );
  FAX1 U465 ( .A(n661), .B(n663), .C(n676), .YC(n683), .YS(n682) );
  FAX1 U466 ( .A(n680), .B(n678), .C(n665), .YC(n685), .YS(n684) );
  FAX1 U467 ( .A(n667), .B(n682), .C(n669), .YC(n687), .YS(n686) );
  FAX1 U468 ( .A(n684), .B(n671), .C(n686), .YC(n689), .YS(n688) );
  FAX1 U469 ( .A(n675), .B(n532), .C(n469), .YC(n691), .YS(n690) );
  FAX1 U470 ( .A(n485), .B(n501), .C(n517), .YC(n693), .YS(n692) );
  FAX1 U471 ( .A(n437), .B(n453), .C(n421), .YC(n695), .YS(n694) );
  FAX1 U472 ( .A(n677), .B(n679), .C(n681), .YC(n697), .YS(n696) );
  FAX1 U473 ( .A(n690), .B(n692), .C(n694), .YC(n699), .YS(n698) );
  FAX1 U474 ( .A(n683), .B(n696), .C(n685), .YC(n701), .YS(n700) );
  FAX1 U475 ( .A(n698), .B(n687), .C(n700), .YC(n703), .YS(n702) );
  INVX2 U476 ( .A(n705), .Y(n704) );
  FAX1 U477 ( .A(n704), .B(n438), .C(n454), .YC(n707), .YS(n706) );
  FAX1 U478 ( .A(n518), .B(n470), .C(n486), .YC(n709), .YS(n708) );
  FAX1 U479 ( .A(n502), .B(n691), .C(n693), .YC(n711), .YS(n710) );
  FAX1 U480 ( .A(n706), .B(n708), .C(n695), .YC(n713), .YS(n712) );
  FAX1 U481 ( .A(n697), .B(n710), .C(n699), .YC(n715), .YS(n714) );
  FAX1 U482 ( .A(n712), .B(n701), .C(n714), .YC(n717), .YS(n716) );
  FAX1 U483 ( .A(n705), .B(n533), .C(n471), .YC(n719), .YS(n718) );
  FAX1 U484 ( .A(n487), .B(n519), .C(n455), .YC(n721), .YS(n720) );
  FAX1 U485 ( .A(n503), .B(n439), .C(n707), .YC(n723), .YS(n722) );
  FAX1 U486 ( .A(n709), .B(n718), .C(n720), .YC(n725), .YS(n724) );
  FAX1 U487 ( .A(n711), .B(n722), .C(n713), .YC(n727), .YS(n726) );
  FAX1 U488 ( .A(n724), .B(n715), .C(n726), .YC(n729), .YS(n728) );
  INVX2 U489 ( .A(n731), .Y(n730) );
  FAX1 U490 ( .A(n730), .B(n456), .C(n472), .YC(n733), .YS(n732) );
  FAX1 U491 ( .A(n520), .B(n504), .C(n488), .YC(n735), .YS(n734) );
  FAX1 U492 ( .A(n719), .B(n721), .C(n732), .YC(n737), .YS(n736) );
  FAX1 U493 ( .A(n734), .B(n723), .C(n725), .YC(n739), .YS(n738) );
  FAX1 U494 ( .A(n736), .B(n727), .C(n738), .YC(n741), .YS(n740) );
  FAX1 U495 ( .A(n731), .B(n534), .C(n489), .YC(n743), .YS(n742) );
  FAX1 U496 ( .A(n505), .B(n521), .C(n473), .YC(n745), .YS(n744) );
  FAX1 U497 ( .A(n457), .B(n733), .C(n735), .YC(n747), .YS(n746) );
  FAX1 U498 ( .A(n742), .B(n744), .C(n737), .YC(n749), .YS(n748) );
  FAX1 U499 ( .A(n746), .B(n739), .C(n748), .YC(n751), .YS(n750) );
  INVX2 U500 ( .A(n753), .Y(n752) );
  FAX1 U501 ( .A(n752), .B(n474), .C(n490), .YC(n755), .YS(n754) );
  FAX1 U502 ( .A(n506), .B(n522), .C(n743), .YC(n757), .YS(n756) );
  FAX1 U503 ( .A(n745), .B(n754), .C(n756), .YC(n759), .YS(n758) );
  FAX1 U504 ( .A(n747), .B(n749), .C(n758), .YC(n761), .YS(n760) );
  FAX1 U505 ( .A(n753), .B(n535), .C(n491), .YC(n763), .YS(n762) );
  FAX1 U506 ( .A(n523), .B(n507), .C(n475), .YC(n765), .YS(n764) );
  FAX1 U507 ( .A(n755), .B(n762), .C(n764), .YC(n767), .YS(n766) );
  FAX1 U508 ( .A(n757), .B(n766), .C(n759), .YC(n769), .YS(n768) );
  INVX2 U509 ( .A(n771), .Y(n770) );
  FAX1 U510 ( .A(n770), .B(n492), .C(n508), .YC(n773), .YS(n772) );
  FAX1 U511 ( .A(n524), .B(n763), .C(n772), .YC(n775), .YS(n774) );
  FAX1 U512 ( .A(n765), .B(n774), .C(n767), .YC(n777), .YS(n776) );
  FAX1 U513 ( .A(n771), .B(n536), .C(n509), .YC(n779), .YS(n778) );
  FAX1 U514 ( .A(n525), .B(n493), .C(n773), .YC(n781), .YS(n780) );
  FAX1 U515 ( .A(n778), .B(n775), .C(n780), .YC(n783), .YS(n782) );
  INVX2 U516 ( .A(n785), .Y(n784) );
  FAX1 U517 ( .A(n784), .B(n510), .C(n526), .YC(n787), .YS(n786) );
  FAX1 U518 ( .A(n779), .B(n786), .C(n781), .YC(n789), .YS(n788) );
  FAX1 U519 ( .A(n785), .B(n537), .C(n527), .YC(n791), .YS(n790) );
  FAX1 U520 ( .A(n511), .B(n787), .C(n790), .YC(n793), .YS(n792) );
  INVX2 U521 ( .A(n795), .Y(n794) );
  FAX1 U522 ( .A(n794), .B(n528), .C(n791), .YC(n797), .YS(n796) );
  HAX1 U523 ( .A(n539), .B(n387), .YC(n799), .YS(product[1]) );
  FAX1 U524 ( .A(n388), .B(n799), .C(n944), .YC(n800), .YS(product[2]) );
  FAX1 U525 ( .A(n540), .B(n547), .C(n800), .YC(n801), .YS(product[3]) );
  FAX1 U526 ( .A(n940), .B(n549), .C(n801), .YC(n802), .YS(product[4]) );
  FAX1 U527 ( .A(n550), .B(n553), .C(n802), .YC(n803), .YS(product[5]) );
  FAX1 U528 ( .A(n554), .B(n557), .C(n803), .YC(n804), .YS(product[6]) );
  FAX1 U529 ( .A(n558), .B(n563), .C(n804), .YC(n805), .YS(product[7]) );
  FAX1 U530 ( .A(n564), .B(n569), .C(n805), .YC(n806), .YS(product[8]) );
  FAX1 U531 ( .A(n570), .B(n577), .C(n806), .YC(n807), .YS(product[9]) );
  FAX1 U532 ( .A(n578), .B(n585), .C(n807), .YC(n808), .YS(product[10]) );
  FAX1 U533 ( .A(n586), .B(n595), .C(n808), .YC(n809), .YS(product[11]) );
  FAX1 U534 ( .A(n596), .B(n605), .C(n809), .YC(n810), .YS(product[12]) );
  FAX1 U535 ( .A(n606), .B(n617), .C(n810), .YC(n811), .YS(product[13]) );
  FAX1 U536 ( .A(n618), .B(n629), .C(n811), .YC(n812), .YS(product[14]) );
  FAX1 U537 ( .A(n630), .B(n643), .C(n812), .YC(n813), .YS(product[15]) );
  FAX1 U538 ( .A(n644), .B(n657), .C(n813), .YC(n814), .YS(product[16]) );
  FAX1 U539 ( .A(n658), .B(n672), .C(n814), .YC(n815), .YS(product[17]) );
  FAX1 U540 ( .A(n673), .B(n688), .C(n815), .YC(n816), .YS(product[18]) );
  FAX1 U541 ( .A(n689), .B(n702), .C(n816), .YC(n817), .YS(product[19]) );
  FAX1 U542 ( .A(n703), .B(n716), .C(n817), .YC(n818), .YS(product[20]) );
  FAX1 U543 ( .A(n717), .B(n728), .C(n818), .YC(n819), .YS(product[21]) );
  FAX1 U544 ( .A(n729), .B(n740), .C(n819), .YC(n820), .YS(product[22]) );
  FAX1 U545 ( .A(n741), .B(n750), .C(n820), .YC(n821), .YS(product[23]) );
  FAX1 U546 ( .A(n751), .B(n760), .C(n821), .YC(n822), .YS(product[24]) );
  FAX1 U547 ( .A(n761), .B(n768), .C(n822), .YC(n823), .YS(product[25]) );
  FAX1 U548 ( .A(n776), .B(n769), .C(n823), .YC(n824), .YS(product[26]) );
  FAX1 U549 ( .A(n782), .B(n777), .C(n824), .YC(n825), .YS(product[27]) );
  FAX1 U550 ( .A(n788), .B(n783), .C(n825), .YC(n826), .YS(product[28]) );
  FAX1 U551 ( .A(n792), .B(n789), .C(n826), .YC(n827), .YS(product[29]) );
  FAX1 U552 ( .A(n796), .B(n793), .C(n827), .YC(n828), .YS(product[30]) );
  XOR2X1 U553 ( .A(n797), .B(n798), .Y(n829) );
  XOR2X1 U554 ( .A(n828), .B(n829), .Y(product[31]) );
  AND2X2 U607 ( .A(n831), .B(a[0]), .Y(product[0]) );
  AND2X2 U608 ( .A(n830), .B(n134), .Y(n940) );
  AND2X2 U609 ( .A(n830), .B(n86), .Y(n941) );
  AND2X2 U610 ( .A(n830), .B(n60), .Y(n942) );
  AND2X2 U611 ( .A(n830), .B(n118), .Y(n943) );
  AND2X2 U612 ( .A(n831), .B(n150), .Y(n944) );
  AND2X2 U613 ( .A(n830), .B(n26), .Y(n945) );
  AND2X2 U614 ( .A(n830), .B(n102), .Y(n946) );
  AND2X2 U615 ( .A(n830), .B(a[15]), .Y(n947) );
  BUFX2 U616 ( .A(n205), .Y(n845) );
  BUFX2 U617 ( .A(n206), .Y(n843) );
  BUFX2 U618 ( .A(n207), .Y(n841) );
  BUFX2 U619 ( .A(n208), .Y(n839) );
  BUFX2 U620 ( .A(n209), .Y(n837) );
  BUFX2 U621 ( .A(n210), .Y(n835) );
  BUFX2 U622 ( .A(n211), .Y(n833) );
  BUFX2 U623 ( .A(n204), .Y(n847) );
  BUFX2 U624 ( .A(n196), .Y(n861) );
  BUFX2 U625 ( .A(n197), .Y(n859) );
  BUFX2 U626 ( .A(n198), .Y(n857) );
  BUFX2 U627 ( .A(n199), .Y(n855) );
  BUFX2 U628 ( .A(n200), .Y(n853) );
  BUFX2 U629 ( .A(n201), .Y(n851) );
  BUFX2 U630 ( .A(n202), .Y(n849) );
  BUFX2 U631 ( .A(n196), .Y(n860) );
  BUFX2 U632 ( .A(n197), .Y(n858) );
  BUFX2 U633 ( .A(n198), .Y(n856) );
  BUFX2 U634 ( .A(n199), .Y(n854) );
  BUFX2 U635 ( .A(n200), .Y(n852) );
  BUFX2 U636 ( .A(n201), .Y(n850) );
  BUFX2 U637 ( .A(n202), .Y(n848) );
  BUFX2 U638 ( .A(n195), .Y(n862) );
  BUFX2 U639 ( .A(n205), .Y(n844) );
  BUFX2 U640 ( .A(n206), .Y(n842) );
  BUFX2 U641 ( .A(n207), .Y(n840) );
  BUFX2 U642 ( .A(n208), .Y(n838) );
  BUFX2 U643 ( .A(n209), .Y(n836) );
  BUFX2 U644 ( .A(n211), .Y(n832) );
  BUFX2 U645 ( .A(n210), .Y(n834) );
  BUFX2 U646 ( .A(n204), .Y(n846) );
  BUFX2 U647 ( .A(n195), .Y(n863) );
  BUFX2 U648 ( .A(b[0]), .Y(n831) );
  BUFX2 U649 ( .A(a[1]), .Y(n879) );
  BUFX2 U650 ( .A(a[5]), .Y(n875) );
  BUFX2 U651 ( .A(a[3]), .Y(n877) );
  BUFX2 U652 ( .A(a[7]), .Y(n873) );
  BUFX2 U653 ( .A(a[9]), .Y(n871) );
  BUFX2 U654 ( .A(a[11]), .Y(n869) );
  BUFX2 U655 ( .A(a[13]), .Y(n867) );
  BUFX2 U656 ( .A(a[15]), .Y(n865) );
  BUFX2 U657 ( .A(a[1]), .Y(n878) );
  BUFX2 U658 ( .A(a[3]), .Y(n876) );
  BUFX2 U659 ( .A(a[5]), .Y(n874) );
  BUFX2 U660 ( .A(a[7]), .Y(n872) );
  BUFX2 U661 ( .A(a[9]), .Y(n870) );
  BUFX2 U662 ( .A(a[11]), .Y(n868) );
  BUFX2 U663 ( .A(a[13]), .Y(n866) );
  BUFX2 U664 ( .A(a[15]), .Y(n864) );
  BUFX2 U665 ( .A(n178), .Y(n203) );
  BUFX2 U666 ( .A(b[0]), .Y(n830) );
  BUFX2 U667 ( .A(b[1]), .Y(n221) );
  BUFX2 U668 ( .A(b[2]), .Y(n222) );
  BUFX2 U669 ( .A(b[3]), .Y(n223) );
  BUFX2 U670 ( .A(b[4]), .Y(n224) );
  BUFX2 U671 ( .A(b[5]), .Y(n225) );
  BUFX2 U672 ( .A(b[6]), .Y(n226) );
  BUFX2 U673 ( .A(b[7]), .Y(n227) );
endmodule


module alu_DW_mult_uns_5 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n15, n25, n26, n50, n60, n80, n85, n86, n101, n102, n117, n118, n133,
         n134, n149, n150, n160, n165, n176, n178, n187, n188, n189, n190,
         n191, n192, n193, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n221, n222, n223, n224, n225,
         n226, n227, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n939,
         n940, n941, n942, n943, n944, n945, n947;

  NAND2X1 OR_NOTi ( .A(n176), .B(n878), .Y(n236) );
  INVX1 U1 ( .A(n831), .Y(n176) );
  OAI21X1 AO21i ( .A(n165), .B(a[0]), .C(a[1]), .Y(n403) );
  INVX1 U12 ( .A(n846), .Y(n165) );
  NAND2X1 OR_NOTi1 ( .A(n160), .B(n876), .Y(n253) );
  INVX1 U13 ( .A(n831), .Y(n160) );
  OAI21X1 AO21i1 ( .A(n149), .B(n150), .C(a[3]), .Y(n421) );
  INVX1 U23 ( .A(n860), .Y(n150) );
  INVX1 U15 ( .A(n844), .Y(n149) );
  NAND2X1 OR_NOTi2 ( .A(n160), .B(n874), .Y(n270) );
  OAI21X1 AO21i2 ( .A(n133), .B(n134), .C(a[5]), .Y(n439) );
  INVX1 U25 ( .A(n858), .Y(n134) );
  INVX1 U18 ( .A(n842), .Y(n133) );
  NAND2X1 OR_NOTi3 ( .A(n160), .B(n872), .Y(n287) );
  OAI21X1 AO21i3 ( .A(n117), .B(n118), .C(a[7]), .Y(n457) );
  INVX1 U27 ( .A(n856), .Y(n118) );
  INVX1 U111 ( .A(n840), .Y(n117) );
  NAND2X1 OR_NOTi4 ( .A(n80), .B(n870), .Y(n304) );
  OAI21X1 AO21i4 ( .A(n101), .B(n102), .C(a[9]), .Y(n475) );
  INVX1 U29 ( .A(n854), .Y(n102) );
  INVX1 U114 ( .A(n838), .Y(n101) );
  NAND2X1 OR_NOTi5 ( .A(n80), .B(n868), .Y(n321) );
  OAI21X1 AO21i5 ( .A(n85), .B(n86), .C(a[11]), .Y(n493) );
  INVX1 U211 ( .A(n852), .Y(n86) );
  INVX1 U117 ( .A(n836), .Y(n85) );
  NAND2X1 OR_NOTi6 ( .A(n80), .B(n866), .Y(n338) );
  INVX1 U118 ( .A(n830), .Y(n80) );
  OAI21X1 AO21i6 ( .A(n50), .B(n60), .C(a[13]), .Y(n511) );
  INVX1 U213 ( .A(n850), .Y(n60) );
  INVX1 U120 ( .A(n834), .Y(n50) );
  NAND2X1 OR_NOTi7 ( .A(n176), .B(n864), .Y(n355) );
  OAI21X1 AO21i7 ( .A(n25), .B(n26), .C(a[15]), .Y(n529) );
  INVX1 U215 ( .A(n848), .Y(n26) );
  INVX1 U123 ( .A(n832), .Y(n25) );
  XOR2X1 U217 ( .A(n538), .B(n795), .Y(n15) );
  XOR2X1 U125 ( .A(n529), .B(n15), .Y(n798) );
  INVX2 U4 ( .A(a[0]), .Y(n195) );
  XOR2X1 U5 ( .A(a[0]), .B(a[1]), .Y(n212) );
  NAND2X1 U6 ( .A(n195), .B(n212), .Y(n204) );
  XNOR2X1 U7 ( .A(a[2]), .B(a[1]), .Y(n196) );
  XOR2X1 U8 ( .A(a[2]), .B(a[3]), .Y(n213) );
  NAND2X1 U9 ( .A(n213), .B(n196), .Y(n205) );
  XNOR2X1 U10 ( .A(a[4]), .B(a[3]), .Y(n197) );
  XOR2X1 U20 ( .A(a[4]), .B(a[5]), .Y(n214) );
  NAND2X1 U30 ( .A(n214), .B(n197), .Y(n206) );
  XNOR2X1 U38 ( .A(a[6]), .B(a[5]), .Y(n198) );
  XOR2X1 U39 ( .A(a[6]), .B(a[7]), .Y(n215) );
  NAND2X1 U40 ( .A(n215), .B(n198), .Y(n207) );
  XNOR2X1 U41 ( .A(a[8]), .B(a[7]), .Y(n199) );
  XOR2X1 U42 ( .A(a[8]), .B(a[9]), .Y(n216) );
  NAND2X1 U43 ( .A(n216), .B(n199), .Y(n208) );
  XNOR2X1 U44 ( .A(a[10]), .B(a[9]), .Y(n200) );
  XOR2X1 U45 ( .A(a[10]), .B(a[11]), .Y(n217) );
  NAND2X1 U46 ( .A(n217), .B(n200), .Y(n209) );
  XNOR2X1 U47 ( .A(a[12]), .B(a[11]), .Y(n201) );
  XOR2X1 U48 ( .A(a[12]), .B(a[13]), .Y(n218) );
  NAND2X1 U49 ( .A(n218), .B(n201), .Y(n210) );
  XNOR2X1 U50 ( .A(a[14]), .B(a[13]), .Y(n202) );
  XOR2X1 U51 ( .A(a[14]), .B(a[15]), .Y(n219) );
  NAND2X1 U52 ( .A(n219), .B(n202), .Y(n211) );
  INVX2 U53 ( .A(a[15]), .Y(n178) );
  INVX2 U54 ( .A(n879), .Y(n187) );
  INVX2 U55 ( .A(n877), .Y(n188) );
  INVX2 U56 ( .A(n875), .Y(n189) );
  INVX2 U57 ( .A(n873), .Y(n190) );
  INVX2 U58 ( .A(n871), .Y(n191) );
  INVX2 U59 ( .A(n869), .Y(n192) );
  INVX2 U60 ( .A(n867), .Y(n193) );
  XNOR2X1 U78 ( .A(n879), .B(n831), .Y(n237) );
  XNOR2X1 U79 ( .A(n879), .B(n221), .Y(n238) );
  XNOR2X1 U80 ( .A(n879), .B(n222), .Y(n239) );
  XNOR2X1 U81 ( .A(n879), .B(n223), .Y(n240) );
  XNOR2X1 U82 ( .A(n879), .B(n224), .Y(n241) );
  XNOR2X1 U83 ( .A(n879), .B(n225), .Y(n242) );
  XNOR2X1 U84 ( .A(n879), .B(n226), .Y(n243) );
  XNOR2X1 U85 ( .A(n879), .B(n227), .Y(n244) );
  XNOR2X1 U86 ( .A(n878), .B(b[8]), .Y(n245) );
  XNOR2X1 U87 ( .A(n878), .B(b[9]), .Y(n246) );
  XNOR2X1 U88 ( .A(n878), .B(b[10]), .Y(n247) );
  XNOR2X1 U89 ( .A(n878), .B(b[11]), .Y(n248) );
  XNOR2X1 U90 ( .A(n878), .B(b[12]), .Y(n249) );
  XNOR2X1 U91 ( .A(n878), .B(b[13]), .Y(n250) );
  XNOR2X1 U92 ( .A(n878), .B(b[14]), .Y(n251) );
  XNOR2X1 U93 ( .A(n878), .B(b[15]), .Y(n252) );
  OAI22X1 U94 ( .A(n863), .B(n238), .C(n237), .D(n847), .Y(n387) );
  OAI22X1 U95 ( .A(n863), .B(n239), .C(n238), .D(n847), .Y(n388) );
  OAI22X1 U96 ( .A(n863), .B(n240), .C(n239), .D(n847), .Y(n389) );
  OAI22X1 U97 ( .A(n863), .B(n241), .C(n240), .D(n847), .Y(n390) );
  OAI22X1 U98 ( .A(n863), .B(n242), .C(n241), .D(n847), .Y(n391) );
  OAI22X1 U99 ( .A(n863), .B(n243), .C(n242), .D(n847), .Y(n392) );
  OAI22X1 U100 ( .A(n863), .B(n244), .C(n243), .D(n847), .Y(n393) );
  OAI22X1 U101 ( .A(n863), .B(n245), .C(n244), .D(n847), .Y(n394) );
  OAI22X1 U102 ( .A(n863), .B(n246), .C(n245), .D(n847), .Y(n395) );
  OAI22X1 U103 ( .A(n862), .B(n247), .C(n246), .D(n846), .Y(n396) );
  OAI22X1 U104 ( .A(n862), .B(n248), .C(n247), .D(n846), .Y(n397) );
  OAI22X1 U105 ( .A(n862), .B(n249), .C(n248), .D(n846), .Y(n398) );
  OAI22X1 U106 ( .A(n862), .B(n250), .C(n249), .D(n846), .Y(n399) );
  OAI22X1 U107 ( .A(n862), .B(n251), .C(n250), .D(n846), .Y(n400) );
  OAI22X1 U108 ( .A(n862), .B(n252), .C(n251), .D(n846), .Y(n401) );
  OAI22X1 U109 ( .A(n862), .B(n187), .C(n252), .D(n846), .Y(n402) );
  OAI22X1 U127 ( .A(n862), .B(n236), .C(n187), .D(n846), .Y(n539) );
  XNOR2X1 U128 ( .A(n877), .B(n831), .Y(n254) );
  XNOR2X1 U129 ( .A(n877), .B(n221), .Y(n255) );
  XNOR2X1 U130 ( .A(n877), .B(n222), .Y(n256) );
  XNOR2X1 U131 ( .A(n877), .B(n223), .Y(n257) );
  XNOR2X1 U132 ( .A(n877), .B(n224), .Y(n258) );
  XNOR2X1 U133 ( .A(n877), .B(n225), .Y(n259) );
  XNOR2X1 U134 ( .A(n877), .B(n226), .Y(n260) );
  XNOR2X1 U135 ( .A(n877), .B(n227), .Y(n261) );
  XNOR2X1 U136 ( .A(n876), .B(b[8]), .Y(n262) );
  XNOR2X1 U137 ( .A(n876), .B(b[9]), .Y(n263) );
  XNOR2X1 U138 ( .A(n876), .B(b[10]), .Y(n264) );
  XNOR2X1 U139 ( .A(n876), .B(b[11]), .Y(n265) );
  XNOR2X1 U140 ( .A(n876), .B(b[12]), .Y(n266) );
  XNOR2X1 U141 ( .A(n876), .B(b[13]), .Y(n267) );
  XNOR2X1 U142 ( .A(n876), .B(b[14]), .Y(n268) );
  XNOR2X1 U143 ( .A(n876), .B(b[15]), .Y(n269) );
  OAI22X1 U144 ( .A(n255), .B(n861), .C(n254), .D(n845), .Y(n405) );
  OAI22X1 U145 ( .A(n256), .B(n861), .C(n255), .D(n845), .Y(n406) );
  OAI22X1 U146 ( .A(n257), .B(n861), .C(n256), .D(n845), .Y(n407) );
  OAI22X1 U147 ( .A(n258), .B(n861), .C(n257), .D(n845), .Y(n408) );
  OAI22X1 U148 ( .A(n259), .B(n861), .C(n258), .D(n845), .Y(n409) );
  OAI22X1 U149 ( .A(n260), .B(n861), .C(n259), .D(n845), .Y(n410) );
  OAI22X1 U150 ( .A(n261), .B(n861), .C(n260), .D(n845), .Y(n411) );
  OAI22X1 U151 ( .A(n262), .B(n861), .C(n261), .D(n845), .Y(n412) );
  OAI22X1 U152 ( .A(n263), .B(n861), .C(n262), .D(n845), .Y(n413) );
  OAI22X1 U153 ( .A(n264), .B(n860), .C(n263), .D(n844), .Y(n414) );
  OAI22X1 U154 ( .A(n265), .B(n860), .C(n264), .D(n844), .Y(n415) );
  OAI22X1 U155 ( .A(n266), .B(n860), .C(n265), .D(n844), .Y(n416) );
  OAI22X1 U156 ( .A(n267), .B(n860), .C(n266), .D(n844), .Y(n417) );
  OAI22X1 U157 ( .A(n268), .B(n860), .C(n267), .D(n844), .Y(n418) );
  OAI22X1 U158 ( .A(n269), .B(n860), .C(n268), .D(n844), .Y(n419) );
  OAI22X1 U159 ( .A(n188), .B(n860), .C(n269), .D(n844), .Y(n420) );
  OAI22X1 U160 ( .A(n860), .B(n253), .C(n188), .D(n844), .Y(n540) );
  XNOR2X1 U161 ( .A(n875), .B(n831), .Y(n271) );
  XNOR2X1 U162 ( .A(n875), .B(n221), .Y(n272) );
  XNOR2X1 U163 ( .A(n875), .B(n222), .Y(n273) );
  XNOR2X1 U164 ( .A(n875), .B(n223), .Y(n274) );
  XNOR2X1 U165 ( .A(n875), .B(n224), .Y(n275) );
  XNOR2X1 U166 ( .A(n875), .B(n225), .Y(n276) );
  XNOR2X1 U167 ( .A(n875), .B(n226), .Y(n277) );
  XNOR2X1 U168 ( .A(n875), .B(n227), .Y(n278) );
  XNOR2X1 U169 ( .A(n874), .B(b[8]), .Y(n279) );
  XNOR2X1 U170 ( .A(n874), .B(b[9]), .Y(n280) );
  XNOR2X1 U171 ( .A(n874), .B(b[10]), .Y(n281) );
  XNOR2X1 U172 ( .A(n874), .B(b[11]), .Y(n282) );
  XNOR2X1 U173 ( .A(n874), .B(b[12]), .Y(n283) );
  XNOR2X1 U174 ( .A(n874), .B(b[13]), .Y(n284) );
  XNOR2X1 U175 ( .A(n874), .B(b[14]), .Y(n285) );
  XNOR2X1 U176 ( .A(n874), .B(b[15]), .Y(n286) );
  OAI22X1 U177 ( .A(n272), .B(n859), .C(n271), .D(n843), .Y(n423) );
  OAI22X1 U178 ( .A(n273), .B(n859), .C(n272), .D(n843), .Y(n424) );
  OAI22X1 U179 ( .A(n274), .B(n859), .C(n273), .D(n843), .Y(n425) );
  OAI22X1 U180 ( .A(n275), .B(n859), .C(n274), .D(n843), .Y(n426) );
  OAI22X1 U181 ( .A(n276), .B(n859), .C(n275), .D(n843), .Y(n427) );
  OAI22X1 U182 ( .A(n277), .B(n859), .C(n276), .D(n843), .Y(n428) );
  OAI22X1 U183 ( .A(n278), .B(n859), .C(n277), .D(n843), .Y(n429) );
  OAI22X1 U184 ( .A(n279), .B(n859), .C(n278), .D(n843), .Y(n430) );
  OAI22X1 U185 ( .A(n280), .B(n859), .C(n279), .D(n843), .Y(n431) );
  OAI22X1 U186 ( .A(n281), .B(n858), .C(n280), .D(n842), .Y(n432) );
  OAI22X1 U187 ( .A(n282), .B(n858), .C(n281), .D(n842), .Y(n433) );
  OAI22X1 U188 ( .A(n283), .B(n858), .C(n282), .D(n842), .Y(n434) );
  OAI22X1 U189 ( .A(n284), .B(n858), .C(n283), .D(n842), .Y(n435) );
  OAI22X1 U190 ( .A(n285), .B(n858), .C(n284), .D(n842), .Y(n436) );
  OAI22X1 U191 ( .A(n286), .B(n858), .C(n285), .D(n842), .Y(n437) );
  OAI22X1 U192 ( .A(n189), .B(n858), .C(n286), .D(n842), .Y(n438) );
  OAI22X1 U193 ( .A(n858), .B(n270), .C(n189), .D(n842), .Y(n541) );
  XNOR2X1 U194 ( .A(n873), .B(n831), .Y(n288) );
  XNOR2X1 U195 ( .A(n873), .B(n221), .Y(n289) );
  XNOR2X1 U196 ( .A(n873), .B(n222), .Y(n290) );
  XNOR2X1 U197 ( .A(n873), .B(n223), .Y(n291) );
  XNOR2X1 U198 ( .A(n873), .B(n224), .Y(n292) );
  XNOR2X1 U199 ( .A(n873), .B(n225), .Y(n293) );
  XNOR2X1 U200 ( .A(n873), .B(n226), .Y(n294) );
  XNOR2X1 U201 ( .A(n873), .B(n227), .Y(n295) );
  XNOR2X1 U202 ( .A(n872), .B(b[8]), .Y(n296) );
  XNOR2X1 U203 ( .A(n872), .B(b[9]), .Y(n297) );
  XNOR2X1 U204 ( .A(n872), .B(b[10]), .Y(n298) );
  XNOR2X1 U205 ( .A(n872), .B(b[11]), .Y(n299) );
  XNOR2X1 U206 ( .A(n872), .B(b[12]), .Y(n300) );
  XNOR2X1 U207 ( .A(n872), .B(b[13]), .Y(n301) );
  XNOR2X1 U208 ( .A(n872), .B(b[14]), .Y(n302) );
  XNOR2X1 U209 ( .A(n872), .B(b[15]), .Y(n303) );
  OAI22X1 U218 ( .A(n289), .B(n857), .C(n288), .D(n841), .Y(n441) );
  OAI22X1 U219 ( .A(n290), .B(n857), .C(n289), .D(n841), .Y(n442) );
  OAI22X1 U220 ( .A(n291), .B(n857), .C(n290), .D(n841), .Y(n443) );
  OAI22X1 U221 ( .A(n292), .B(n857), .C(n291), .D(n841), .Y(n444) );
  OAI22X1 U222 ( .A(n293), .B(n857), .C(n292), .D(n841), .Y(n445) );
  OAI22X1 U223 ( .A(n294), .B(n857), .C(n293), .D(n841), .Y(n446) );
  OAI22X1 U224 ( .A(n295), .B(n857), .C(n294), .D(n841), .Y(n447) );
  OAI22X1 U225 ( .A(n296), .B(n857), .C(n295), .D(n841), .Y(n448) );
  OAI22X1 U226 ( .A(n297), .B(n857), .C(n296), .D(n841), .Y(n449) );
  OAI22X1 U227 ( .A(n298), .B(n856), .C(n297), .D(n840), .Y(n450) );
  OAI22X1 U228 ( .A(n299), .B(n856), .C(n298), .D(n840), .Y(n451) );
  OAI22X1 U229 ( .A(n300), .B(n856), .C(n299), .D(n840), .Y(n452) );
  OAI22X1 U230 ( .A(n301), .B(n856), .C(n300), .D(n840), .Y(n453) );
  OAI22X1 U231 ( .A(n302), .B(n856), .C(n301), .D(n840), .Y(n454) );
  OAI22X1 U232 ( .A(n303), .B(n856), .C(n302), .D(n840), .Y(n455) );
  OAI22X1 U233 ( .A(n190), .B(n856), .C(n303), .D(n840), .Y(n456) );
  OAI22X1 U234 ( .A(n856), .B(n287), .C(n190), .D(n840), .Y(n542) );
  XNOR2X1 U235 ( .A(n871), .B(n831), .Y(n305) );
  XNOR2X1 U236 ( .A(n871), .B(n221), .Y(n306) );
  XNOR2X1 U237 ( .A(n871), .B(n222), .Y(n307) );
  XNOR2X1 U238 ( .A(n871), .B(n223), .Y(n308) );
  XNOR2X1 U239 ( .A(n871), .B(n224), .Y(n309) );
  XNOR2X1 U240 ( .A(n871), .B(n225), .Y(n310) );
  XNOR2X1 U241 ( .A(n871), .B(n226), .Y(n311) );
  XNOR2X1 U242 ( .A(n871), .B(n227), .Y(n312) );
  XNOR2X1 U243 ( .A(n870), .B(b[8]), .Y(n313) );
  XNOR2X1 U244 ( .A(n870), .B(b[9]), .Y(n314) );
  XNOR2X1 U245 ( .A(n870), .B(b[10]), .Y(n315) );
  XNOR2X1 U246 ( .A(n870), .B(b[11]), .Y(n316) );
  XNOR2X1 U247 ( .A(n870), .B(b[12]), .Y(n317) );
  XNOR2X1 U248 ( .A(n870), .B(b[13]), .Y(n318) );
  XNOR2X1 U249 ( .A(n870), .B(b[14]), .Y(n319) );
  XNOR2X1 U250 ( .A(n870), .B(b[15]), .Y(n320) );
  OAI22X1 U251 ( .A(n306), .B(n855), .C(n305), .D(n839), .Y(n459) );
  OAI22X1 U252 ( .A(n307), .B(n855), .C(n306), .D(n839), .Y(n460) );
  OAI22X1 U253 ( .A(n308), .B(n855), .C(n307), .D(n839), .Y(n461) );
  OAI22X1 U254 ( .A(n309), .B(n855), .C(n308), .D(n839), .Y(n462) );
  OAI22X1 U255 ( .A(n310), .B(n855), .C(n309), .D(n839), .Y(n463) );
  OAI22X1 U256 ( .A(n311), .B(n855), .C(n310), .D(n839), .Y(n464) );
  OAI22X1 U257 ( .A(n312), .B(n855), .C(n311), .D(n839), .Y(n465) );
  OAI22X1 U258 ( .A(n313), .B(n855), .C(n312), .D(n839), .Y(n466) );
  OAI22X1 U259 ( .A(n314), .B(n855), .C(n313), .D(n839), .Y(n467) );
  OAI22X1 U260 ( .A(n315), .B(n854), .C(n314), .D(n838), .Y(n468) );
  OAI22X1 U261 ( .A(n316), .B(n854), .C(n315), .D(n838), .Y(n469) );
  OAI22X1 U262 ( .A(n317), .B(n854), .C(n316), .D(n838), .Y(n470) );
  OAI22X1 U263 ( .A(n318), .B(n854), .C(n317), .D(n838), .Y(n471) );
  OAI22X1 U264 ( .A(n319), .B(n854), .C(n318), .D(n838), .Y(n472) );
  OAI22X1 U265 ( .A(n320), .B(n854), .C(n319), .D(n838), .Y(n473) );
  OAI22X1 U266 ( .A(n191), .B(n854), .C(n320), .D(n838), .Y(n474) );
  OAI22X1 U267 ( .A(n854), .B(n304), .C(n191), .D(n838), .Y(n543) );
  XNOR2X1 U268 ( .A(n869), .B(n831), .Y(n322) );
  XNOR2X1 U269 ( .A(n869), .B(n221), .Y(n323) );
  XNOR2X1 U270 ( .A(n869), .B(n222), .Y(n324) );
  XNOR2X1 U271 ( .A(n869), .B(n223), .Y(n325) );
  XNOR2X1 U272 ( .A(n869), .B(n224), .Y(n326) );
  XNOR2X1 U273 ( .A(n869), .B(n225), .Y(n327) );
  XNOR2X1 U274 ( .A(n869), .B(n226), .Y(n328) );
  XNOR2X1 U275 ( .A(n869), .B(n227), .Y(n329) );
  XNOR2X1 U276 ( .A(n868), .B(b[8]), .Y(n330) );
  XNOR2X1 U277 ( .A(n868), .B(b[9]), .Y(n331) );
  XNOR2X1 U278 ( .A(n868), .B(b[10]), .Y(n332) );
  XNOR2X1 U279 ( .A(n868), .B(b[11]), .Y(n333) );
  XNOR2X1 U280 ( .A(n868), .B(b[12]), .Y(n334) );
  XNOR2X1 U281 ( .A(n868), .B(b[13]), .Y(n335) );
  XNOR2X1 U282 ( .A(n868), .B(b[14]), .Y(n336) );
  XNOR2X1 U283 ( .A(n868), .B(b[15]), .Y(n337) );
  OAI22X1 U284 ( .A(n323), .B(n853), .C(n322), .D(n837), .Y(n477) );
  OAI22X1 U285 ( .A(n324), .B(n853), .C(n323), .D(n837), .Y(n478) );
  OAI22X1 U286 ( .A(n325), .B(n853), .C(n324), .D(n837), .Y(n479) );
  OAI22X1 U287 ( .A(n326), .B(n853), .C(n325), .D(n837), .Y(n480) );
  OAI22X1 U288 ( .A(n327), .B(n853), .C(n326), .D(n837), .Y(n481) );
  OAI22X1 U289 ( .A(n328), .B(n853), .C(n327), .D(n837), .Y(n482) );
  OAI22X1 U290 ( .A(n329), .B(n853), .C(n328), .D(n837), .Y(n483) );
  OAI22X1 U291 ( .A(n330), .B(n853), .C(n329), .D(n837), .Y(n484) );
  OAI22X1 U292 ( .A(n331), .B(n853), .C(n330), .D(n837), .Y(n485) );
  OAI22X1 U293 ( .A(n332), .B(n852), .C(n331), .D(n836), .Y(n486) );
  OAI22X1 U294 ( .A(n333), .B(n852), .C(n332), .D(n836), .Y(n487) );
  OAI22X1 U295 ( .A(n334), .B(n852), .C(n333), .D(n836), .Y(n488) );
  OAI22X1 U296 ( .A(n335), .B(n852), .C(n334), .D(n836), .Y(n489) );
  OAI22X1 U297 ( .A(n336), .B(n852), .C(n335), .D(n836), .Y(n490) );
  OAI22X1 U298 ( .A(n337), .B(n852), .C(n336), .D(n836), .Y(n491) );
  OAI22X1 U299 ( .A(n192), .B(n852), .C(n337), .D(n836), .Y(n492) );
  OAI22X1 U300 ( .A(n852), .B(n321), .C(n192), .D(n836), .Y(n544) );
  XNOR2X1 U301 ( .A(n867), .B(n831), .Y(n339) );
  XNOR2X1 U302 ( .A(n867), .B(n221), .Y(n340) );
  XNOR2X1 U303 ( .A(n867), .B(n222), .Y(n341) );
  XNOR2X1 U304 ( .A(n867), .B(n223), .Y(n342) );
  XNOR2X1 U305 ( .A(n867), .B(n224), .Y(n343) );
  XNOR2X1 U306 ( .A(n867), .B(n225), .Y(n344) );
  XNOR2X1 U307 ( .A(n867), .B(n226), .Y(n345) );
  XNOR2X1 U308 ( .A(n867), .B(n227), .Y(n346) );
  XNOR2X1 U309 ( .A(n866), .B(b[8]), .Y(n347) );
  XNOR2X1 U310 ( .A(n866), .B(b[9]), .Y(n348) );
  XNOR2X1 U311 ( .A(n866), .B(b[10]), .Y(n349) );
  XNOR2X1 U312 ( .A(n866), .B(b[11]), .Y(n350) );
  XNOR2X1 U313 ( .A(n866), .B(b[12]), .Y(n351) );
  XNOR2X1 U314 ( .A(n866), .B(b[13]), .Y(n352) );
  XNOR2X1 U315 ( .A(n866), .B(b[14]), .Y(n353) );
  XNOR2X1 U316 ( .A(n866), .B(b[15]), .Y(n354) );
  OAI22X1 U317 ( .A(n340), .B(n851), .C(n339), .D(n835), .Y(n495) );
  OAI22X1 U318 ( .A(n341), .B(n851), .C(n340), .D(n835), .Y(n496) );
  OAI22X1 U319 ( .A(n342), .B(n851), .C(n341), .D(n835), .Y(n497) );
  OAI22X1 U320 ( .A(n343), .B(n851), .C(n342), .D(n835), .Y(n498) );
  OAI22X1 U321 ( .A(n344), .B(n851), .C(n343), .D(n835), .Y(n499) );
  OAI22X1 U322 ( .A(n345), .B(n851), .C(n344), .D(n835), .Y(n500) );
  OAI22X1 U323 ( .A(n346), .B(n851), .C(n345), .D(n835), .Y(n501) );
  OAI22X1 U324 ( .A(n347), .B(n851), .C(n346), .D(n835), .Y(n502) );
  OAI22X1 U325 ( .A(n348), .B(n851), .C(n347), .D(n835), .Y(n503) );
  OAI22X1 U326 ( .A(n349), .B(n850), .C(n348), .D(n834), .Y(n504) );
  OAI22X1 U327 ( .A(n350), .B(n850), .C(n349), .D(n834), .Y(n505) );
  OAI22X1 U328 ( .A(n351), .B(n850), .C(n350), .D(n834), .Y(n506) );
  OAI22X1 U329 ( .A(n352), .B(n850), .C(n351), .D(n834), .Y(n507) );
  OAI22X1 U330 ( .A(n353), .B(n850), .C(n352), .D(n834), .Y(n508) );
  OAI22X1 U331 ( .A(n354), .B(n850), .C(n353), .D(n834), .Y(n509) );
  OAI22X1 U332 ( .A(n193), .B(n850), .C(n354), .D(n834), .Y(n510) );
  OAI22X1 U333 ( .A(n850), .B(n338), .C(n193), .D(n834), .Y(n545) );
  XNOR2X1 U334 ( .A(n865), .B(n831), .Y(n356) );
  XNOR2X1 U335 ( .A(n865), .B(n221), .Y(n357) );
  XNOR2X1 U336 ( .A(n865), .B(n222), .Y(n358) );
  XNOR2X1 U337 ( .A(n865), .B(n223), .Y(n359) );
  XNOR2X1 U338 ( .A(n865), .B(n224), .Y(n360) );
  XNOR2X1 U339 ( .A(n865), .B(n225), .Y(n361) );
  XNOR2X1 U340 ( .A(n865), .B(n226), .Y(n362) );
  XNOR2X1 U341 ( .A(n865), .B(n227), .Y(n363) );
  XNOR2X1 U342 ( .A(n864), .B(b[8]), .Y(n364) );
  XNOR2X1 U343 ( .A(n864), .B(b[9]), .Y(n365) );
  XNOR2X1 U344 ( .A(n864), .B(b[10]), .Y(n366) );
  XNOR2X1 U345 ( .A(n864), .B(b[11]), .Y(n367) );
  XNOR2X1 U346 ( .A(n864), .B(b[12]), .Y(n368) );
  XNOR2X1 U347 ( .A(n864), .B(b[13]), .Y(n369) );
  XNOR2X1 U348 ( .A(n864), .B(b[14]), .Y(n370) );
  XNOR2X1 U349 ( .A(n864), .B(b[15]), .Y(n371) );
  OAI22X1 U350 ( .A(n357), .B(n849), .C(n356), .D(n833), .Y(n513) );
  OAI22X1 U351 ( .A(n358), .B(n849), .C(n357), .D(n833), .Y(n514) );
  OAI22X1 U352 ( .A(n359), .B(n849), .C(n358), .D(n833), .Y(n515) );
  OAI22X1 U353 ( .A(n360), .B(n849), .C(n359), .D(n833), .Y(n516) );
  OAI22X1 U354 ( .A(n361), .B(n849), .C(n360), .D(n833), .Y(n517) );
  OAI22X1 U355 ( .A(n362), .B(n849), .C(n361), .D(n833), .Y(n518) );
  OAI22X1 U356 ( .A(n363), .B(n849), .C(n362), .D(n833), .Y(n519) );
  OAI22X1 U357 ( .A(n364), .B(n849), .C(n363), .D(n833), .Y(n520) );
  OAI22X1 U358 ( .A(n365), .B(n849), .C(n364), .D(n833), .Y(n521) );
  OAI22X1 U359 ( .A(n366), .B(n848), .C(n365), .D(n832), .Y(n522) );
  OAI22X1 U360 ( .A(n367), .B(n848), .C(n366), .D(n832), .Y(n523) );
  OAI22X1 U361 ( .A(n368), .B(n848), .C(n367), .D(n832), .Y(n524) );
  OAI22X1 U362 ( .A(n369), .B(n848), .C(n368), .D(n832), .Y(n525) );
  OAI22X1 U363 ( .A(n370), .B(n848), .C(n369), .D(n832), .Y(n526) );
  OAI22X1 U364 ( .A(n371), .B(n848), .C(n370), .D(n832), .Y(n527) );
  OAI22X1 U365 ( .A(n178), .B(n848), .C(n371), .D(n832), .Y(n528) );
  OAI22X1 U366 ( .A(n848), .B(n355), .C(n178), .D(n832), .Y(n546) );
  INVX2 U367 ( .A(n221), .Y(n372) );
  INVX2 U368 ( .A(n222), .Y(n373) );
  INVX2 U369 ( .A(n223), .Y(n374) );
  INVX2 U370 ( .A(n224), .Y(n375) );
  INVX2 U371 ( .A(n225), .Y(n376) );
  INVX2 U372 ( .A(n226), .Y(n377) );
  INVX2 U373 ( .A(n227), .Y(n378) );
  INVX2 U374 ( .A(b[8]), .Y(n379) );
  INVX2 U375 ( .A(b[9]), .Y(n380) );
  INVX2 U376 ( .A(b[10]), .Y(n381) );
  INVX2 U377 ( .A(b[11]), .Y(n382) );
  INVX2 U378 ( .A(b[12]), .Y(n383) );
  INVX2 U379 ( .A(b[13]), .Y(n384) );
  INVX2 U380 ( .A(b[14]), .Y(n385) );
  INVX2 U381 ( .A(b[15]), .Y(n386) );
  NOR2X1 U382 ( .A(n372), .B(n203), .Y(n675) );
  NOR2X1 U383 ( .A(n373), .B(n203), .Y(n531) );
  NOR2X1 U384 ( .A(n374), .B(n203), .Y(n532) );
  NOR2X1 U385 ( .A(n375), .B(n203), .Y(n705) );
  NOR2X1 U386 ( .A(n376), .B(n203), .Y(n533) );
  NOR2X1 U387 ( .A(n377), .B(n203), .Y(n731) );
  NOR2X1 U388 ( .A(n378), .B(n203), .Y(n534) );
  NOR2X1 U389 ( .A(n379), .B(n203), .Y(n753) );
  NOR2X1 U390 ( .A(n380), .B(n203), .Y(n535) );
  NOR2X1 U391 ( .A(n381), .B(n203), .Y(n771) );
  NOR2X1 U392 ( .A(n382), .B(n203), .Y(n536) );
  NOR2X1 U393 ( .A(n383), .B(n203), .Y(n785) );
  NOR2X1 U394 ( .A(n384), .B(n203), .Y(n537) );
  NOR2X1 U395 ( .A(n385), .B(n203), .Y(n795) );
  NOR2X1 U396 ( .A(n386), .B(n203), .Y(n538) );
  HAX1 U397 ( .A(n389), .B(n405), .YC(n548), .YS(n547) );
  FAX1 U398 ( .A(n390), .B(n406), .C(n548), .YC(n550), .YS(n549) );
  HAX1 U399 ( .A(n391), .B(n541), .YC(n552), .YS(n551) );
  FAX1 U400 ( .A(n407), .B(n423), .C(n551), .YC(n554), .YS(n553) );
  FAX1 U401 ( .A(n392), .B(n424), .C(n408), .YC(n556), .YS(n555) );
  FAX1 U402 ( .A(n552), .B(n942), .C(n555), .YC(n558), .YS(n557) );
  HAX1 U403 ( .A(n393), .B(n542), .YC(n560), .YS(n559) );
  FAX1 U404 ( .A(n409), .B(n441), .C(n425), .YC(n562), .YS(n561) );
  FAX1 U405 ( .A(n559), .B(n556), .C(n561), .YC(n564), .YS(n563) );
  FAX1 U406 ( .A(n394), .B(n426), .C(n442), .YC(n566), .YS(n565) );
  FAX1 U407 ( .A(n410), .B(n560), .C(n945), .YC(n568), .YS(n567) );
  FAX1 U408 ( .A(n562), .B(n565), .C(n567), .YC(n570), .YS(n569) );
  HAX1 U409 ( .A(n395), .B(n543), .YC(n572), .YS(n571) );
  FAX1 U410 ( .A(n443), .B(n459), .C(n427), .YC(n574), .YS(n573) );
  FAX1 U411 ( .A(n411), .B(n571), .C(n566), .YC(n576), .YS(n575) );
  FAX1 U412 ( .A(n573), .B(n568), .C(n575), .YC(n578), .YS(n577) );
  FAX1 U413 ( .A(n396), .B(n412), .C(n428), .YC(n580), .YS(n579) );
  FAX1 U414 ( .A(n444), .B(n460), .C(n572), .YC(n582), .YS(n581) );
  FAX1 U415 ( .A(n940), .B(n574), .C(n579), .YC(n584), .YS(n583) );
  FAX1 U416 ( .A(n581), .B(n576), .C(n583), .YC(n586), .YS(n585) );
  HAX1 U417 ( .A(n397), .B(n544), .YC(n588), .YS(n587) );
  FAX1 U418 ( .A(n445), .B(n477), .C(n413), .YC(n590), .YS(n589) );
  FAX1 U419 ( .A(n429), .B(n461), .C(n587), .YC(n592), .YS(n591) );
  FAX1 U420 ( .A(n580), .B(n589), .C(n582), .YC(n594), .YS(n593) );
  FAX1 U421 ( .A(n591), .B(n584), .C(n593), .YC(n596), .YS(n595) );
  FAX1 U422 ( .A(n398), .B(n414), .C(n478), .YC(n598), .YS(n597) );
  FAX1 U423 ( .A(n430), .B(n462), .C(n446), .YC(n600), .YS(n599) );
  FAX1 U424 ( .A(n588), .B(n941), .C(n590), .YC(n602), .YS(n601) );
  FAX1 U425 ( .A(n597), .B(n599), .C(n592), .YC(n604), .YS(n603) );
  FAX1 U426 ( .A(n601), .B(n594), .C(n603), .YC(n606), .YS(n605) );
  HAX1 U427 ( .A(n399), .B(n545), .YC(n608), .YS(n607) );
  FAX1 U428 ( .A(n463), .B(n415), .C(n431), .YC(n610), .YS(n609) );
  FAX1 U429 ( .A(n447), .B(n495), .C(n479), .YC(n612), .YS(n611) );
  FAX1 U430 ( .A(n607), .B(n598), .C(n600), .YC(n614), .YS(n613) );
  FAX1 U431 ( .A(n611), .B(n609), .C(n602), .YC(n616), .YS(n615) );
  FAX1 U432 ( .A(n613), .B(n604), .C(n615), .YC(n618), .YS(n617) );
  FAX1 U433 ( .A(n400), .B(n416), .C(n432), .YC(n620), .YS(n619) );
  FAX1 U434 ( .A(n448), .B(n496), .C(n480), .YC(n622), .YS(n621) );
  FAX1 U435 ( .A(n464), .B(n608), .C(n944), .YC(n624), .YS(n623) );
  FAX1 U436 ( .A(n610), .B(n612), .C(n619), .YC(n626), .YS(n625) );
  FAX1 U437 ( .A(n621), .B(n623), .C(n614), .YC(n628), .YS(n627) );
  FAX1 U438 ( .A(n625), .B(n616), .C(n627), .YC(n630), .YS(n629) );
  HAX1 U439 ( .A(n401), .B(n546), .YC(n632), .YS(n631) );
  FAX1 U440 ( .A(n465), .B(n513), .C(n497), .YC(n634), .YS(n633) );
  FAX1 U441 ( .A(n417), .B(n481), .C(n449), .YC(n636), .YS(n635) );
  FAX1 U442 ( .A(n433), .B(n631), .C(n620), .YC(n638), .YS(n637) );
  FAX1 U443 ( .A(n622), .B(n635), .C(n633), .YC(n640), .YS(n639) );
  FAX1 U444 ( .A(n624), .B(n626), .C(n637), .YC(n642), .YS(n641) );
  FAX1 U445 ( .A(n639), .B(n628), .C(n641), .YC(n644), .YS(n643) );
  FAX1 U446 ( .A(n402), .B(n418), .C(n947), .YC(n646), .YS(n645) );
  FAX1 U447 ( .A(n434), .B(n514), .C(n498), .YC(n648), .YS(n647) );
  FAX1 U448 ( .A(n450), .B(n482), .C(n466), .YC(n650), .YS(n649) );
  FAX1 U449 ( .A(n632), .B(n634), .C(n636), .YC(n652), .YS(n651) );
  FAX1 U450 ( .A(n645), .B(n649), .C(n647), .YC(n654), .YS(n653) );
  FAX1 U451 ( .A(n638), .B(n640), .C(n651), .YC(n656), .YS(n655) );
  FAX1 U452 ( .A(n653), .B(n642), .C(n655), .YC(n658), .YS(n657) );
  INVX2 U453 ( .A(n675), .Y(n659) );
  FAX1 U454 ( .A(n659), .B(n499), .C(n451), .YC(n661), .YS(n660) );
  FAX1 U455 ( .A(n467), .B(n483), .C(n515), .YC(n663), .YS(n662) );
  FAX1 U456 ( .A(n419), .B(n435), .C(n403), .YC(n665), .YS(n664) );
  FAX1 U457 ( .A(n646), .B(n648), .C(n650), .YC(n667), .YS(n666) );
  FAX1 U458 ( .A(n660), .B(n662), .C(n664), .YC(n669), .YS(n668) );
  FAX1 U459 ( .A(n652), .B(n654), .C(n666), .YC(n671), .YS(n670) );
  FAX1 U460 ( .A(n668), .B(n656), .C(n670), .YC(n673), .YS(n672) );
  FAX1 U462 ( .A(n531), .B(n659), .C(n420), .YC(n677), .YS(n676) );
  FAX1 U463 ( .A(n436), .B(n516), .C(n452), .YC(n679), .YS(n678) );
  FAX1 U464 ( .A(n468), .B(n500), .C(n484), .YC(n681), .YS(n680) );
  FAX1 U465 ( .A(n661), .B(n663), .C(n676), .YC(n683), .YS(n682) );
  FAX1 U466 ( .A(n680), .B(n678), .C(n665), .YC(n685), .YS(n684) );
  FAX1 U467 ( .A(n667), .B(n682), .C(n669), .YC(n687), .YS(n686) );
  FAX1 U468 ( .A(n684), .B(n671), .C(n686), .YC(n689), .YS(n688) );
  FAX1 U469 ( .A(n675), .B(n532), .C(n469), .YC(n691), .YS(n690) );
  FAX1 U470 ( .A(n485), .B(n501), .C(n517), .YC(n693), .YS(n692) );
  FAX1 U471 ( .A(n437), .B(n453), .C(n421), .YC(n695), .YS(n694) );
  FAX1 U472 ( .A(n677), .B(n679), .C(n681), .YC(n697), .YS(n696) );
  FAX1 U473 ( .A(n690), .B(n692), .C(n694), .YC(n699), .YS(n698) );
  FAX1 U474 ( .A(n683), .B(n696), .C(n685), .YC(n701), .YS(n700) );
  FAX1 U475 ( .A(n698), .B(n687), .C(n700), .YC(n703), .YS(n702) );
  INVX2 U476 ( .A(n705), .Y(n704) );
  FAX1 U477 ( .A(n704), .B(n438), .C(n454), .YC(n707), .YS(n706) );
  FAX1 U478 ( .A(n518), .B(n470), .C(n486), .YC(n709), .YS(n708) );
  FAX1 U479 ( .A(n502), .B(n691), .C(n693), .YC(n711), .YS(n710) );
  FAX1 U480 ( .A(n706), .B(n708), .C(n695), .YC(n713), .YS(n712) );
  FAX1 U481 ( .A(n697), .B(n710), .C(n699), .YC(n715), .YS(n714) );
  FAX1 U482 ( .A(n712), .B(n701), .C(n714), .YC(n717), .YS(n716) );
  FAX1 U483 ( .A(n705), .B(n533), .C(n471), .YC(n719), .YS(n718) );
  FAX1 U484 ( .A(n487), .B(n519), .C(n455), .YC(n721), .YS(n720) );
  FAX1 U485 ( .A(n503), .B(n439), .C(n707), .YC(n723), .YS(n722) );
  FAX1 U486 ( .A(n709), .B(n718), .C(n720), .YC(n725), .YS(n724) );
  FAX1 U487 ( .A(n711), .B(n722), .C(n713), .YC(n727), .YS(n726) );
  FAX1 U488 ( .A(n724), .B(n715), .C(n726), .YC(n729), .YS(n728) );
  INVX2 U489 ( .A(n731), .Y(n730) );
  FAX1 U490 ( .A(n730), .B(n456), .C(n472), .YC(n733), .YS(n732) );
  FAX1 U491 ( .A(n520), .B(n504), .C(n488), .YC(n735), .YS(n734) );
  FAX1 U492 ( .A(n719), .B(n721), .C(n732), .YC(n737), .YS(n736) );
  FAX1 U493 ( .A(n734), .B(n723), .C(n725), .YC(n739), .YS(n738) );
  FAX1 U494 ( .A(n736), .B(n727), .C(n738), .YC(n741), .YS(n740) );
  FAX1 U495 ( .A(n731), .B(n534), .C(n489), .YC(n743), .YS(n742) );
  FAX1 U496 ( .A(n505), .B(n521), .C(n473), .YC(n745), .YS(n744) );
  FAX1 U497 ( .A(n457), .B(n733), .C(n735), .YC(n747), .YS(n746) );
  FAX1 U498 ( .A(n742), .B(n744), .C(n737), .YC(n749), .YS(n748) );
  FAX1 U499 ( .A(n746), .B(n739), .C(n748), .YC(n751), .YS(n750) );
  INVX2 U500 ( .A(n753), .Y(n752) );
  FAX1 U501 ( .A(n752), .B(n474), .C(n490), .YC(n755), .YS(n754) );
  FAX1 U502 ( .A(n506), .B(n522), .C(n743), .YC(n757), .YS(n756) );
  FAX1 U503 ( .A(n745), .B(n754), .C(n756), .YC(n759), .YS(n758) );
  FAX1 U504 ( .A(n747), .B(n749), .C(n758), .YC(n761), .YS(n760) );
  FAX1 U505 ( .A(n753), .B(n535), .C(n491), .YC(n763), .YS(n762) );
  FAX1 U506 ( .A(n523), .B(n507), .C(n475), .YC(n765), .YS(n764) );
  FAX1 U507 ( .A(n755), .B(n762), .C(n764), .YC(n767), .YS(n766) );
  FAX1 U508 ( .A(n757), .B(n766), .C(n759), .YC(n769), .YS(n768) );
  INVX2 U509 ( .A(n771), .Y(n770) );
  FAX1 U510 ( .A(n770), .B(n492), .C(n508), .YC(n773), .YS(n772) );
  FAX1 U511 ( .A(n524), .B(n763), .C(n772), .YC(n775), .YS(n774) );
  FAX1 U512 ( .A(n765), .B(n774), .C(n767), .YC(n777), .YS(n776) );
  FAX1 U513 ( .A(n771), .B(n536), .C(n509), .YC(n779), .YS(n778) );
  FAX1 U514 ( .A(n525), .B(n493), .C(n773), .YC(n781), .YS(n780) );
  FAX1 U515 ( .A(n778), .B(n775), .C(n780), .YC(n783), .YS(n782) );
  INVX2 U516 ( .A(n785), .Y(n784) );
  FAX1 U517 ( .A(n784), .B(n510), .C(n526), .YC(n787), .YS(n786) );
  FAX1 U518 ( .A(n779), .B(n786), .C(n781), .YC(n789), .YS(n788) );
  FAX1 U519 ( .A(n785), .B(n537), .C(n527), .YC(n791), .YS(n790) );
  FAX1 U520 ( .A(n511), .B(n787), .C(n790), .YC(n793), .YS(n792) );
  INVX2 U521 ( .A(n795), .Y(n794) );
  FAX1 U522 ( .A(n794), .B(n528), .C(n791), .YC(n797), .YS(n796) );
  HAX1 U523 ( .A(n539), .B(n387), .YC(n799), .YS(product[1]) );
  FAX1 U524 ( .A(n388), .B(n799), .C(n943), .YC(n800), .YS(product[2]) );
  FAX1 U525 ( .A(n540), .B(n547), .C(n800), .YC(n801), .YS(product[3]) );
  FAX1 U526 ( .A(n939), .B(n549), .C(n801), .YC(n802), .YS(product[4]) );
  FAX1 U527 ( .A(n550), .B(n553), .C(n802), .YC(n803), .YS(product[5]) );
  FAX1 U528 ( .A(n554), .B(n557), .C(n803), .YC(n804), .YS(product[6]) );
  FAX1 U529 ( .A(n558), .B(n563), .C(n804), .YC(n805), .YS(product[7]) );
  FAX1 U530 ( .A(n564), .B(n569), .C(n805), .YC(n806), .YS(product[8]) );
  FAX1 U531 ( .A(n570), .B(n577), .C(n806), .YC(n807), .YS(product[9]) );
  FAX1 U532 ( .A(n578), .B(n585), .C(n807), .YC(n808), .YS(product[10]) );
  FAX1 U533 ( .A(n586), .B(n595), .C(n808), .YC(n809), .YS(product[11]) );
  FAX1 U534 ( .A(n596), .B(n605), .C(n809), .YC(n810), .YS(product[12]) );
  FAX1 U535 ( .A(n606), .B(n617), .C(n810), .YC(n811), .YS(product[13]) );
  FAX1 U536 ( .A(n618), .B(n629), .C(n811), .YC(n812), .YS(product[14]) );
  FAX1 U537 ( .A(n630), .B(n643), .C(n812), .YC(n813), .YS(product[15]) );
  FAX1 U538 ( .A(n644), .B(n657), .C(n813), .YC(n814), .YS(product[16]) );
  FAX1 U539 ( .A(n658), .B(n672), .C(n814), .YC(n815), .YS(product[17]) );
  FAX1 U540 ( .A(n673), .B(n688), .C(n815), .YC(n816), .YS(product[18]) );
  FAX1 U541 ( .A(n689), .B(n702), .C(n816), .YC(n817), .YS(product[19]) );
  FAX1 U542 ( .A(n703), .B(n716), .C(n817), .YC(n818), .YS(product[20]) );
  FAX1 U543 ( .A(n717), .B(n728), .C(n818), .YC(n819), .YS(product[21]) );
  FAX1 U544 ( .A(n729), .B(n740), .C(n819), .YC(n820), .YS(product[22]) );
  FAX1 U545 ( .A(n741), .B(n750), .C(n820), .YC(n821), .YS(product[23]) );
  FAX1 U546 ( .A(n751), .B(n760), .C(n821), .YC(n822), .YS(product[24]) );
  FAX1 U547 ( .A(n761), .B(n768), .C(n822), .YC(n823), .YS(product[25]) );
  FAX1 U548 ( .A(n776), .B(n769), .C(n823), .YC(n824), .YS(product[26]) );
  FAX1 U549 ( .A(n782), .B(n777), .C(n824), .YC(n825), .YS(product[27]) );
  FAX1 U550 ( .A(n788), .B(n783), .C(n825), .YC(n826), .YS(product[28]) );
  FAX1 U551 ( .A(n792), .B(n789), .C(n826), .YC(n827), .YS(product[29]) );
  FAX1 U552 ( .A(n796), .B(n793), .C(n827), .YC(n828), .YS(product[30]) );
  XOR2X1 U553 ( .A(n797), .B(n798), .Y(n829) );
  XOR2X1 U554 ( .A(n828), .B(n829), .Y(product[31]) );
  AND2X2 U607 ( .A(n830), .B(n134), .Y(n939) );
  AND2X2 U608 ( .A(n830), .B(n86), .Y(n940) );
  AND2X2 U609 ( .A(n830), .B(n60), .Y(n941) );
  AND2X2 U610 ( .A(n830), .B(n118), .Y(n942) );
  AND2X2 U611 ( .A(n831), .B(n150), .Y(n943) );
  AND2X2 U612 ( .A(n830), .B(n26), .Y(n944) );
  AND2X2 U613 ( .A(n830), .B(n102), .Y(n945) );
  AND2X2 U614 ( .A(n831), .B(a[0]), .Y(product[0]) );
  AND2X2 U615 ( .A(n830), .B(a[15]), .Y(n947) );
  BUFX2 U616 ( .A(n205), .Y(n845) );
  BUFX2 U617 ( .A(n206), .Y(n843) );
  BUFX2 U618 ( .A(n207), .Y(n841) );
  BUFX2 U619 ( .A(n208), .Y(n839) );
  BUFX2 U620 ( .A(n209), .Y(n837) );
  BUFX2 U621 ( .A(n210), .Y(n835) );
  BUFX2 U622 ( .A(n211), .Y(n833) );
  BUFX2 U623 ( .A(n204), .Y(n847) );
  BUFX2 U624 ( .A(n196), .Y(n861) );
  BUFX2 U625 ( .A(n197), .Y(n859) );
  BUFX2 U626 ( .A(n198), .Y(n857) );
  BUFX2 U627 ( .A(n199), .Y(n855) );
  BUFX2 U628 ( .A(n200), .Y(n853) );
  BUFX2 U629 ( .A(n201), .Y(n851) );
  BUFX2 U630 ( .A(n202), .Y(n849) );
  BUFX2 U631 ( .A(n196), .Y(n860) );
  BUFX2 U632 ( .A(n197), .Y(n858) );
  BUFX2 U633 ( .A(n198), .Y(n856) );
  BUFX2 U634 ( .A(n199), .Y(n854) );
  BUFX2 U635 ( .A(n200), .Y(n852) );
  BUFX2 U636 ( .A(n201), .Y(n850) );
  BUFX2 U637 ( .A(n202), .Y(n848) );
  BUFX2 U638 ( .A(n195), .Y(n862) );
  BUFX2 U639 ( .A(n205), .Y(n844) );
  BUFX2 U640 ( .A(n206), .Y(n842) );
  BUFX2 U641 ( .A(n207), .Y(n840) );
  BUFX2 U642 ( .A(n208), .Y(n838) );
  BUFX2 U643 ( .A(n209), .Y(n836) );
  BUFX2 U644 ( .A(n211), .Y(n832) );
  BUFX2 U645 ( .A(n210), .Y(n834) );
  BUFX2 U646 ( .A(n204), .Y(n846) );
  BUFX2 U647 ( .A(n195), .Y(n863) );
  BUFX2 U648 ( .A(b[0]), .Y(n831) );
  BUFX2 U649 ( .A(a[1]), .Y(n879) );
  BUFX2 U650 ( .A(a[5]), .Y(n875) );
  BUFX2 U651 ( .A(a[3]), .Y(n877) );
  BUFX2 U652 ( .A(a[7]), .Y(n873) );
  BUFX2 U653 ( .A(a[9]), .Y(n871) );
  BUFX2 U654 ( .A(a[11]), .Y(n869) );
  BUFX2 U655 ( .A(a[13]), .Y(n867) );
  BUFX2 U656 ( .A(a[15]), .Y(n865) );
  BUFX2 U657 ( .A(a[1]), .Y(n878) );
  BUFX2 U658 ( .A(a[3]), .Y(n876) );
  BUFX2 U659 ( .A(a[5]), .Y(n874) );
  BUFX2 U660 ( .A(a[7]), .Y(n872) );
  BUFX2 U661 ( .A(a[9]), .Y(n870) );
  BUFX2 U662 ( .A(a[11]), .Y(n868) );
  BUFX2 U663 ( .A(a[13]), .Y(n866) );
  BUFX2 U664 ( .A(a[15]), .Y(n864) );
  BUFX2 U665 ( .A(n178), .Y(n203) );
  BUFX2 U666 ( .A(b[0]), .Y(n830) );
  BUFX2 U667 ( .A(b[1]), .Y(n221) );
  BUFX2 U668 ( .A(b[2]), .Y(n222) );
  BUFX2 U669 ( .A(b[3]), .Y(n223) );
  BUFX2 U670 ( .A(b[4]), .Y(n224) );
  BUFX2 U671 ( .A(b[5]), .Y(n225) );
  BUFX2 U672 ( .A(b[6]), .Y(n226) );
  BUFX2 U673 ( .A(b[7]), .Y(n227) );
endmodule


module alu_DW_mult_uns_6 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176;

  NOR2X1 U17 ( .A(n1), .B(n9), .Y(product[0]) );
  NOR2X1 U18 ( .A(n1), .B(n10), .Y(n17) );
  NOR2X1 U19 ( .A(n1), .B(n11), .Y(n18) );
  NOR2X1 U20 ( .A(n1), .B(n12), .Y(n19) );
  NOR2X1 U21 ( .A(n1), .B(n13), .Y(n20) );
  NOR2X1 U22 ( .A(n1), .B(n14), .Y(n21) );
  NOR2X1 U23 ( .A(n1), .B(n15), .Y(n22) );
  NOR2X1 U24 ( .A(n1), .B(n16), .Y(n23) );
  NOR2X1 U25 ( .A(n2), .B(n9), .Y(n24) );
  NOR2X1 U26 ( .A(n2), .B(n10), .Y(n25) );
  NOR2X1 U27 ( .A(n2), .B(n11), .Y(n26) );
  NOR2X1 U28 ( .A(n2), .B(n12), .Y(n27) );
  NOR2X1 U29 ( .A(n2), .B(n13), .Y(n28) );
  NOR2X1 U30 ( .A(n2), .B(n14), .Y(n29) );
  NOR2X1 U31 ( .A(n2), .B(n15), .Y(n30) );
  NOR2X1 U32 ( .A(n2), .B(n16), .Y(n31) );
  NOR2X1 U33 ( .A(n3), .B(n9), .Y(n32) );
  NOR2X1 U34 ( .A(n3), .B(n10), .Y(n33) );
  NOR2X1 U35 ( .A(n3), .B(n11), .Y(n34) );
  NOR2X1 U36 ( .A(n3), .B(n12), .Y(n35) );
  NOR2X1 U37 ( .A(n3), .B(n13), .Y(n36) );
  NOR2X1 U38 ( .A(n3), .B(n14), .Y(n37) );
  NOR2X1 U39 ( .A(n3), .B(n15), .Y(n38) );
  NOR2X1 U40 ( .A(n3), .B(n16), .Y(n39) );
  NOR2X1 U41 ( .A(n4), .B(n9), .Y(n40) );
  NOR2X1 U42 ( .A(n4), .B(n10), .Y(n41) );
  NOR2X1 U43 ( .A(n4), .B(n11), .Y(n42) );
  NOR2X1 U44 ( .A(n4), .B(n12), .Y(n43) );
  NOR2X1 U45 ( .A(n4), .B(n13), .Y(n44) );
  NOR2X1 U46 ( .A(n4), .B(n14), .Y(n45) );
  NOR2X1 U47 ( .A(n4), .B(n15), .Y(n46) );
  NOR2X1 U48 ( .A(n4), .B(n16), .Y(n47) );
  NOR2X1 U49 ( .A(n5), .B(n9), .Y(n48) );
  NOR2X1 U50 ( .A(n5), .B(n10), .Y(n49) );
  NOR2X1 U51 ( .A(n5), .B(n11), .Y(n50) );
  NOR2X1 U52 ( .A(n5), .B(n12), .Y(n51) );
  NOR2X1 U53 ( .A(n5), .B(n13), .Y(n52) );
  NOR2X1 U54 ( .A(n5), .B(n14), .Y(n53) );
  NOR2X1 U55 ( .A(n5), .B(n15), .Y(n54) );
  NOR2X1 U56 ( .A(n5), .B(n16), .Y(n55) );
  NOR2X1 U57 ( .A(n6), .B(n9), .Y(n56) );
  NOR2X1 U58 ( .A(n6), .B(n10), .Y(n57) );
  NOR2X1 U59 ( .A(n6), .B(n11), .Y(n58) );
  NOR2X1 U60 ( .A(n6), .B(n12), .Y(n59) );
  NOR2X1 U61 ( .A(n6), .B(n13), .Y(n60) );
  NOR2X1 U62 ( .A(n6), .B(n14), .Y(n61) );
  NOR2X1 U63 ( .A(n6), .B(n15), .Y(n62) );
  NOR2X1 U64 ( .A(n6), .B(n16), .Y(n63) );
  NOR2X1 U65 ( .A(n7), .B(n9), .Y(n64) );
  NOR2X1 U66 ( .A(n7), .B(n10), .Y(n65) );
  NOR2X1 U67 ( .A(n7), .B(n11), .Y(n66) );
  NOR2X1 U68 ( .A(n7), .B(n12), .Y(n67) );
  NOR2X1 U69 ( .A(n7), .B(n13), .Y(n68) );
  NOR2X1 U70 ( .A(n7), .B(n14), .Y(n69) );
  NOR2X1 U71 ( .A(n7), .B(n15), .Y(n70) );
  NOR2X1 U72 ( .A(n7), .B(n16), .Y(n71) );
  NOR2X1 U73 ( .A(n8), .B(n9), .Y(n72) );
  NOR2X1 U74 ( .A(n8), .B(n10), .Y(n73) );
  NOR2X1 U75 ( .A(n8), .B(n11), .Y(n74) );
  NOR2X1 U76 ( .A(n8), .B(n12), .Y(n75) );
  NOR2X1 U77 ( .A(n8), .B(n13), .Y(n76) );
  NOR2X1 U78 ( .A(n8), .B(n14), .Y(n77) );
  NOR2X1 U79 ( .A(n8), .B(n15), .Y(n78) );
  NOR2X1 U80 ( .A(n8), .B(n16), .Y(n79) );
  HAX1 U81 ( .A(n18), .B(n25), .YC(n81), .YS(n80) );
  HAX1 U82 ( .A(n33), .B(n40), .YC(n83), .YS(n82) );
  FAX1 U83 ( .A(n19), .B(n26), .C(n81), .YC(n85), .YS(n84) );
  HAX1 U84 ( .A(n41), .B(n48), .YC(n87), .YS(n86) );
  FAX1 U85 ( .A(n20), .B(n34), .C(n27), .YC(n89), .YS(n88) );
  FAX1 U86 ( .A(n83), .B(n86), .C(n88), .YC(n91), .YS(n90) );
  HAX1 U87 ( .A(n49), .B(n56), .YC(n93), .YS(n92) );
  FAX1 U88 ( .A(n21), .B(n42), .C(n35), .YC(n95), .YS(n94) );
  FAX1 U89 ( .A(n28), .B(n87), .C(n92), .YC(n97), .YS(n96) );
  FAX1 U90 ( .A(n89), .B(n94), .C(n96), .YC(n99), .YS(n98) );
  HAX1 U91 ( .A(n57), .B(n64), .YC(n101), .YS(n100) );
  FAX1 U92 ( .A(n22), .B(n50), .C(n29), .YC(n103), .YS(n102) );
  FAX1 U93 ( .A(n36), .B(n43), .C(n93), .YC(n105), .YS(n104) );
  FAX1 U94 ( .A(n100), .B(n95), .C(n102), .YC(n107), .YS(n106) );
  FAX1 U95 ( .A(n97), .B(n104), .C(n106), .YC(n109), .YS(n108) );
  HAX1 U96 ( .A(n65), .B(n72), .YC(n111), .YS(n110) );
  FAX1 U97 ( .A(n23), .B(n58), .C(n30), .YC(n113), .YS(n112) );
  FAX1 U98 ( .A(n37), .B(n51), .C(n44), .YC(n115), .YS(n114) );
  FAX1 U99 ( .A(n101), .B(n110), .C(n103), .YC(n117), .YS(n116) );
  FAX1 U100 ( .A(n114), .B(n112), .C(n105), .YC(n119), .YS(n118) );
  FAX1 U101 ( .A(n107), .B(n116), .C(n118), .YC(n121), .YS(n120) );
  HAX1 U102 ( .A(n66), .B(n73), .YC(n123), .YS(n122) );
  FAX1 U103 ( .A(n52), .B(n59), .C(n31), .YC(n125), .YS(n124) );
  FAX1 U104 ( .A(n38), .B(n45), .C(n111), .YC(n127), .YS(n126) );
  FAX1 U105 ( .A(n122), .B(n113), .C(n115), .YC(n129), .YS(n128) );
  FAX1 U106 ( .A(n124), .B(n126), .C(n117), .YC(n131), .YS(n130) );
  FAX1 U107 ( .A(n128), .B(n119), .C(n130), .YC(n133), .YS(n132) );
  FAX1 U108 ( .A(n39), .B(n74), .C(n67), .YC(n135), .YS(n134) );
  FAX1 U109 ( .A(n60), .B(n53), .C(n46), .YC(n137), .YS(n136) );
  FAX1 U110 ( .A(n123), .B(n125), .C(n136), .YC(n139), .YS(n138) );
  FAX1 U111 ( .A(n134), .B(n127), .C(n129), .YC(n141), .YS(n140) );
  FAX1 U112 ( .A(n138), .B(n131), .C(n140), .YC(n143), .YS(n142) );
  FAX1 U113 ( .A(n47), .B(n75), .C(n68), .YC(n145), .YS(n144) );
  FAX1 U114 ( .A(n54), .B(n61), .C(n135), .YC(n147), .YS(n146) );
  FAX1 U115 ( .A(n137), .B(n144), .C(n139), .YC(n149), .YS(n148) );
  FAX1 U116 ( .A(n146), .B(n141), .C(n148), .YC(n151), .YS(n150) );
  FAX1 U117 ( .A(n55), .B(n76), .C(n69), .YC(n153), .YS(n152) );
  FAX1 U118 ( .A(n62), .B(n145), .C(n152), .YC(n155), .YS(n154) );
  FAX1 U119 ( .A(n147), .B(n154), .C(n149), .YC(n157), .YS(n156) );
  FAX1 U120 ( .A(n63), .B(n77), .C(n70), .YC(n159), .YS(n158) );
  FAX1 U121 ( .A(n153), .B(n158), .C(n155), .YC(n161), .YS(n160) );
  FAX1 U122 ( .A(n71), .B(n78), .C(n159), .YC(n163), .YS(n162) );
  HAX1 U123 ( .A(n24), .B(n17), .YC(n164), .YS(product[1]) );
  FAX1 U124 ( .A(n32), .B(n164), .C(n80), .YC(n165), .YS(product[2]) );
  FAX1 U125 ( .A(n82), .B(n165), .C(n84), .YC(n166), .YS(product[3]) );
  FAX1 U126 ( .A(n85), .B(n90), .C(n166), .YC(n167), .YS(product[4]) );
  FAX1 U127 ( .A(n91), .B(n98), .C(n167), .YC(n168), .YS(product[5]) );
  FAX1 U128 ( .A(n99), .B(n108), .C(n168), .YC(n169), .YS(product[6]) );
  FAX1 U129 ( .A(n109), .B(n120), .C(n169), .YC(n170), .YS(product[7]) );
  FAX1 U130 ( .A(n121), .B(n132), .C(n170), .YC(n171), .YS(product[8]) );
  FAX1 U131 ( .A(n133), .B(n142), .C(n171), .YC(n172), .YS(product[9]) );
  FAX1 U132 ( .A(n143), .B(n150), .C(n172), .YC(n173), .YS(product[10]) );
  FAX1 U133 ( .A(n151), .B(n156), .C(n173), .YC(n174), .YS(product[11]) );
  FAX1 U134 ( .A(n160), .B(n157), .C(n174), .YC(n175), .YS(product[12]) );
  FAX1 U135 ( .A(n162), .B(n161), .C(n175), .YC(n176), .YS(product[13]) );
  FAX1 U136 ( .A(n79), .B(n163), .C(n176), .YC(product[15]), .YS(product[14])
         );
  INVX2 U140 ( .A(b[0]), .Y(n9) );
  INVX2 U141 ( .A(b[1]), .Y(n10) );
  INVX2 U142 ( .A(b[2]), .Y(n11) );
  INVX2 U143 ( .A(b[3]), .Y(n12) );
  INVX2 U144 ( .A(b[4]), .Y(n13) );
  INVX2 U145 ( .A(b[5]), .Y(n14) );
  INVX2 U146 ( .A(b[6]), .Y(n15) );
  INVX2 U147 ( .A(b[7]), .Y(n16) );
  INVX2 U148 ( .A(a[0]), .Y(n1) );
  INVX2 U149 ( .A(a[1]), .Y(n2) );
  INVX2 U150 ( .A(a[2]), .Y(n3) );
  INVX2 U151 ( .A(a[3]), .Y(n4) );
  INVX2 U152 ( .A(a[4]), .Y(n5) );
  INVX2 U153 ( .A(a[5]), .Y(n6) );
  INVX2 U154 ( .A(a[6]), .Y(n7) );
  INVX2 U155 ( .A(a[7]), .Y(n8) );
endmodule


module alu_DW_mult_uns_7 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n15, n25, n26, n50, n60, n80, n85, n86, n101, n102, n117, n118, n133,
         n134, n149, n150, n160, n165, n176, n178, n187, n188, n189, n190,
         n191, n192, n193, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n221, n222, n223, n224, n225,
         n226, n227, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n940,
         n941, n942, n943, n944, n945, n946, n947;

  NAND2X1 OR_NOTi ( .A(n176), .B(n878), .Y(n236) );
  INVX1 U1 ( .A(n831), .Y(n176) );
  OAI21X1 AO21i ( .A(n165), .B(a[0]), .C(a[1]), .Y(n403) );
  INVX1 U12 ( .A(n846), .Y(n165) );
  NAND2X1 OR_NOTi1 ( .A(n160), .B(n876), .Y(n253) );
  INVX1 U13 ( .A(n831), .Y(n160) );
  OAI21X1 AO21i1 ( .A(n149), .B(n150), .C(a[3]), .Y(n421) );
  INVX1 U23 ( .A(n860), .Y(n150) );
  INVX1 U15 ( .A(n844), .Y(n149) );
  NAND2X1 OR_NOTi2 ( .A(n160), .B(n874), .Y(n270) );
  OAI21X1 AO21i2 ( .A(n133), .B(n134), .C(a[5]), .Y(n439) );
  INVX1 U25 ( .A(n858), .Y(n134) );
  INVX1 U18 ( .A(n842), .Y(n133) );
  NAND2X1 OR_NOTi3 ( .A(n160), .B(n872), .Y(n287) );
  OAI21X1 AO21i3 ( .A(n117), .B(n118), .C(a[7]), .Y(n457) );
  INVX1 U27 ( .A(n856), .Y(n118) );
  INVX1 U111 ( .A(n840), .Y(n117) );
  NAND2X1 OR_NOTi4 ( .A(n80), .B(n870), .Y(n304) );
  OAI21X1 AO21i4 ( .A(n101), .B(n102), .C(a[9]), .Y(n475) );
  INVX1 U29 ( .A(n854), .Y(n102) );
  INVX1 U114 ( .A(n838), .Y(n101) );
  NAND2X1 OR_NOTi5 ( .A(n80), .B(n868), .Y(n321) );
  OAI21X1 AO21i5 ( .A(n85), .B(n86), .C(a[11]), .Y(n493) );
  INVX1 U211 ( .A(n852), .Y(n86) );
  INVX1 U117 ( .A(n836), .Y(n85) );
  NAND2X1 OR_NOTi6 ( .A(n80), .B(n866), .Y(n338) );
  INVX1 U118 ( .A(n830), .Y(n80) );
  OAI21X1 AO21i6 ( .A(n50), .B(n60), .C(a[13]), .Y(n511) );
  INVX1 U213 ( .A(n850), .Y(n60) );
  INVX1 U120 ( .A(n834), .Y(n50) );
  NAND2X1 OR_NOTi7 ( .A(n176), .B(n864), .Y(n355) );
  OAI21X1 AO21i7 ( .A(n25), .B(n26), .C(a[15]), .Y(n529) );
  INVX1 U215 ( .A(n848), .Y(n26) );
  INVX1 U123 ( .A(n832), .Y(n25) );
  XOR2X1 U217 ( .A(n538), .B(n795), .Y(n15) );
  XOR2X1 U125 ( .A(n529), .B(n15), .Y(n798) );
  INVX2 U4 ( .A(a[0]), .Y(n195) );
  XOR2X1 U5 ( .A(a[0]), .B(a[1]), .Y(n212) );
  NAND2X1 U6 ( .A(n195), .B(n212), .Y(n204) );
  XNOR2X1 U7 ( .A(a[2]), .B(a[1]), .Y(n196) );
  XOR2X1 U8 ( .A(a[2]), .B(a[3]), .Y(n213) );
  NAND2X1 U9 ( .A(n213), .B(n196), .Y(n205) );
  XNOR2X1 U10 ( .A(a[4]), .B(a[3]), .Y(n197) );
  XOR2X1 U20 ( .A(a[4]), .B(a[5]), .Y(n214) );
  NAND2X1 U30 ( .A(n214), .B(n197), .Y(n206) );
  XNOR2X1 U38 ( .A(a[6]), .B(a[5]), .Y(n198) );
  XOR2X1 U39 ( .A(a[6]), .B(a[7]), .Y(n215) );
  NAND2X1 U40 ( .A(n215), .B(n198), .Y(n207) );
  XNOR2X1 U41 ( .A(a[8]), .B(a[7]), .Y(n199) );
  XOR2X1 U42 ( .A(a[8]), .B(a[9]), .Y(n216) );
  NAND2X1 U43 ( .A(n216), .B(n199), .Y(n208) );
  XNOR2X1 U44 ( .A(a[10]), .B(a[9]), .Y(n200) );
  XOR2X1 U45 ( .A(a[10]), .B(a[11]), .Y(n217) );
  NAND2X1 U46 ( .A(n217), .B(n200), .Y(n209) );
  XNOR2X1 U47 ( .A(a[12]), .B(a[11]), .Y(n201) );
  XOR2X1 U48 ( .A(a[12]), .B(a[13]), .Y(n218) );
  NAND2X1 U49 ( .A(n218), .B(n201), .Y(n210) );
  XNOR2X1 U50 ( .A(a[14]), .B(a[13]), .Y(n202) );
  XOR2X1 U51 ( .A(a[14]), .B(a[15]), .Y(n219) );
  NAND2X1 U52 ( .A(n219), .B(n202), .Y(n211) );
  INVX2 U53 ( .A(a[15]), .Y(n178) );
  INVX2 U54 ( .A(n879), .Y(n187) );
  INVX2 U55 ( .A(n877), .Y(n188) );
  INVX2 U56 ( .A(n875), .Y(n189) );
  INVX2 U57 ( .A(n873), .Y(n190) );
  INVX2 U58 ( .A(n871), .Y(n191) );
  INVX2 U59 ( .A(n869), .Y(n192) );
  INVX2 U60 ( .A(n867), .Y(n193) );
  XNOR2X1 U78 ( .A(n879), .B(n831), .Y(n237) );
  XNOR2X1 U79 ( .A(n879), .B(n221), .Y(n238) );
  XNOR2X1 U80 ( .A(n879), .B(n222), .Y(n239) );
  XNOR2X1 U81 ( .A(n879), .B(n223), .Y(n240) );
  XNOR2X1 U82 ( .A(n879), .B(n224), .Y(n241) );
  XNOR2X1 U83 ( .A(n879), .B(n225), .Y(n242) );
  XNOR2X1 U84 ( .A(n879), .B(n226), .Y(n243) );
  XNOR2X1 U85 ( .A(n879), .B(n227), .Y(n244) );
  XNOR2X1 U86 ( .A(n878), .B(b[8]), .Y(n245) );
  XNOR2X1 U87 ( .A(n878), .B(b[9]), .Y(n246) );
  XNOR2X1 U88 ( .A(n878), .B(b[10]), .Y(n247) );
  XNOR2X1 U89 ( .A(n878), .B(b[11]), .Y(n248) );
  XNOR2X1 U90 ( .A(n878), .B(b[12]), .Y(n249) );
  XNOR2X1 U91 ( .A(n878), .B(b[13]), .Y(n250) );
  XNOR2X1 U92 ( .A(n878), .B(b[14]), .Y(n251) );
  XNOR2X1 U93 ( .A(n878), .B(b[15]), .Y(n252) );
  OAI22X1 U94 ( .A(n863), .B(n238), .C(n237), .D(n847), .Y(n387) );
  OAI22X1 U95 ( .A(n863), .B(n239), .C(n238), .D(n847), .Y(n388) );
  OAI22X1 U96 ( .A(n863), .B(n240), .C(n239), .D(n847), .Y(n389) );
  OAI22X1 U97 ( .A(n863), .B(n241), .C(n240), .D(n847), .Y(n390) );
  OAI22X1 U98 ( .A(n863), .B(n242), .C(n241), .D(n847), .Y(n391) );
  OAI22X1 U99 ( .A(n863), .B(n243), .C(n242), .D(n847), .Y(n392) );
  OAI22X1 U100 ( .A(n863), .B(n244), .C(n243), .D(n847), .Y(n393) );
  OAI22X1 U101 ( .A(n863), .B(n245), .C(n244), .D(n847), .Y(n394) );
  OAI22X1 U102 ( .A(n863), .B(n246), .C(n245), .D(n847), .Y(n395) );
  OAI22X1 U103 ( .A(n862), .B(n247), .C(n246), .D(n846), .Y(n396) );
  OAI22X1 U104 ( .A(n862), .B(n248), .C(n247), .D(n846), .Y(n397) );
  OAI22X1 U105 ( .A(n862), .B(n249), .C(n248), .D(n846), .Y(n398) );
  OAI22X1 U106 ( .A(n862), .B(n250), .C(n249), .D(n846), .Y(n399) );
  OAI22X1 U107 ( .A(n862), .B(n251), .C(n250), .D(n846), .Y(n400) );
  OAI22X1 U108 ( .A(n862), .B(n252), .C(n251), .D(n846), .Y(n401) );
  OAI22X1 U109 ( .A(n862), .B(n187), .C(n252), .D(n846), .Y(n402) );
  OAI22X1 U127 ( .A(n862), .B(n236), .C(n187), .D(n846), .Y(n539) );
  XNOR2X1 U128 ( .A(n877), .B(n831), .Y(n254) );
  XNOR2X1 U129 ( .A(n877), .B(n221), .Y(n255) );
  XNOR2X1 U130 ( .A(n877), .B(n222), .Y(n256) );
  XNOR2X1 U131 ( .A(n877), .B(n223), .Y(n257) );
  XNOR2X1 U132 ( .A(n877), .B(n224), .Y(n258) );
  XNOR2X1 U133 ( .A(n877), .B(n225), .Y(n259) );
  XNOR2X1 U134 ( .A(n877), .B(n226), .Y(n260) );
  XNOR2X1 U135 ( .A(n877), .B(n227), .Y(n261) );
  XNOR2X1 U136 ( .A(n876), .B(b[8]), .Y(n262) );
  XNOR2X1 U137 ( .A(n876), .B(b[9]), .Y(n263) );
  XNOR2X1 U138 ( .A(n876), .B(b[10]), .Y(n264) );
  XNOR2X1 U139 ( .A(n876), .B(b[11]), .Y(n265) );
  XNOR2X1 U140 ( .A(n876), .B(b[12]), .Y(n266) );
  XNOR2X1 U141 ( .A(n876), .B(b[13]), .Y(n267) );
  XNOR2X1 U142 ( .A(n876), .B(b[14]), .Y(n268) );
  XNOR2X1 U143 ( .A(n876), .B(b[15]), .Y(n269) );
  OAI22X1 U144 ( .A(n255), .B(n861), .C(n254), .D(n845), .Y(n405) );
  OAI22X1 U145 ( .A(n256), .B(n861), .C(n255), .D(n845), .Y(n406) );
  OAI22X1 U146 ( .A(n257), .B(n861), .C(n256), .D(n845), .Y(n407) );
  OAI22X1 U147 ( .A(n258), .B(n861), .C(n257), .D(n845), .Y(n408) );
  OAI22X1 U148 ( .A(n259), .B(n861), .C(n258), .D(n845), .Y(n409) );
  OAI22X1 U149 ( .A(n260), .B(n861), .C(n259), .D(n845), .Y(n410) );
  OAI22X1 U150 ( .A(n261), .B(n861), .C(n260), .D(n845), .Y(n411) );
  OAI22X1 U151 ( .A(n262), .B(n861), .C(n261), .D(n845), .Y(n412) );
  OAI22X1 U152 ( .A(n263), .B(n861), .C(n262), .D(n845), .Y(n413) );
  OAI22X1 U153 ( .A(n264), .B(n860), .C(n263), .D(n844), .Y(n414) );
  OAI22X1 U154 ( .A(n265), .B(n860), .C(n264), .D(n844), .Y(n415) );
  OAI22X1 U155 ( .A(n266), .B(n860), .C(n265), .D(n844), .Y(n416) );
  OAI22X1 U156 ( .A(n267), .B(n860), .C(n266), .D(n844), .Y(n417) );
  OAI22X1 U157 ( .A(n268), .B(n860), .C(n267), .D(n844), .Y(n418) );
  OAI22X1 U158 ( .A(n269), .B(n860), .C(n268), .D(n844), .Y(n419) );
  OAI22X1 U159 ( .A(n188), .B(n860), .C(n269), .D(n844), .Y(n420) );
  OAI22X1 U160 ( .A(n860), .B(n253), .C(n188), .D(n844), .Y(n540) );
  XNOR2X1 U161 ( .A(n875), .B(n831), .Y(n271) );
  XNOR2X1 U162 ( .A(n875), .B(n221), .Y(n272) );
  XNOR2X1 U163 ( .A(n875), .B(n222), .Y(n273) );
  XNOR2X1 U164 ( .A(n875), .B(n223), .Y(n274) );
  XNOR2X1 U165 ( .A(n875), .B(n224), .Y(n275) );
  XNOR2X1 U166 ( .A(n875), .B(n225), .Y(n276) );
  XNOR2X1 U167 ( .A(n875), .B(n226), .Y(n277) );
  XNOR2X1 U168 ( .A(n875), .B(n227), .Y(n278) );
  XNOR2X1 U169 ( .A(n874), .B(b[8]), .Y(n279) );
  XNOR2X1 U170 ( .A(n874), .B(b[9]), .Y(n280) );
  XNOR2X1 U171 ( .A(n874), .B(b[10]), .Y(n281) );
  XNOR2X1 U172 ( .A(n874), .B(b[11]), .Y(n282) );
  XNOR2X1 U173 ( .A(n874), .B(b[12]), .Y(n283) );
  XNOR2X1 U174 ( .A(n874), .B(b[13]), .Y(n284) );
  XNOR2X1 U175 ( .A(n874), .B(b[14]), .Y(n285) );
  XNOR2X1 U176 ( .A(n874), .B(b[15]), .Y(n286) );
  OAI22X1 U177 ( .A(n272), .B(n859), .C(n271), .D(n843), .Y(n423) );
  OAI22X1 U178 ( .A(n273), .B(n859), .C(n272), .D(n843), .Y(n424) );
  OAI22X1 U179 ( .A(n274), .B(n859), .C(n273), .D(n843), .Y(n425) );
  OAI22X1 U180 ( .A(n275), .B(n859), .C(n274), .D(n843), .Y(n426) );
  OAI22X1 U181 ( .A(n276), .B(n859), .C(n275), .D(n843), .Y(n427) );
  OAI22X1 U182 ( .A(n277), .B(n859), .C(n276), .D(n843), .Y(n428) );
  OAI22X1 U183 ( .A(n278), .B(n859), .C(n277), .D(n843), .Y(n429) );
  OAI22X1 U184 ( .A(n279), .B(n859), .C(n278), .D(n843), .Y(n430) );
  OAI22X1 U185 ( .A(n280), .B(n859), .C(n279), .D(n843), .Y(n431) );
  OAI22X1 U186 ( .A(n281), .B(n858), .C(n280), .D(n842), .Y(n432) );
  OAI22X1 U187 ( .A(n282), .B(n858), .C(n281), .D(n842), .Y(n433) );
  OAI22X1 U188 ( .A(n283), .B(n858), .C(n282), .D(n842), .Y(n434) );
  OAI22X1 U189 ( .A(n284), .B(n858), .C(n283), .D(n842), .Y(n435) );
  OAI22X1 U190 ( .A(n285), .B(n858), .C(n284), .D(n842), .Y(n436) );
  OAI22X1 U191 ( .A(n286), .B(n858), .C(n285), .D(n842), .Y(n437) );
  OAI22X1 U192 ( .A(n189), .B(n858), .C(n286), .D(n842), .Y(n438) );
  OAI22X1 U193 ( .A(n858), .B(n270), .C(n189), .D(n842), .Y(n541) );
  XNOR2X1 U194 ( .A(n873), .B(n831), .Y(n288) );
  XNOR2X1 U195 ( .A(n873), .B(n221), .Y(n289) );
  XNOR2X1 U196 ( .A(n873), .B(n222), .Y(n290) );
  XNOR2X1 U197 ( .A(n873), .B(n223), .Y(n291) );
  XNOR2X1 U198 ( .A(n873), .B(n224), .Y(n292) );
  XNOR2X1 U199 ( .A(n873), .B(n225), .Y(n293) );
  XNOR2X1 U200 ( .A(n873), .B(n226), .Y(n294) );
  XNOR2X1 U201 ( .A(n873), .B(n227), .Y(n295) );
  XNOR2X1 U202 ( .A(n872), .B(b[8]), .Y(n296) );
  XNOR2X1 U203 ( .A(n872), .B(b[9]), .Y(n297) );
  XNOR2X1 U204 ( .A(n872), .B(b[10]), .Y(n298) );
  XNOR2X1 U205 ( .A(n872), .B(b[11]), .Y(n299) );
  XNOR2X1 U206 ( .A(n872), .B(b[12]), .Y(n300) );
  XNOR2X1 U207 ( .A(n872), .B(b[13]), .Y(n301) );
  XNOR2X1 U208 ( .A(n872), .B(b[14]), .Y(n302) );
  XNOR2X1 U209 ( .A(n872), .B(b[15]), .Y(n303) );
  OAI22X1 U218 ( .A(n289), .B(n857), .C(n288), .D(n841), .Y(n441) );
  OAI22X1 U219 ( .A(n290), .B(n857), .C(n289), .D(n841), .Y(n442) );
  OAI22X1 U220 ( .A(n291), .B(n857), .C(n290), .D(n841), .Y(n443) );
  OAI22X1 U221 ( .A(n292), .B(n857), .C(n291), .D(n841), .Y(n444) );
  OAI22X1 U222 ( .A(n293), .B(n857), .C(n292), .D(n841), .Y(n445) );
  OAI22X1 U223 ( .A(n294), .B(n857), .C(n293), .D(n841), .Y(n446) );
  OAI22X1 U224 ( .A(n295), .B(n857), .C(n294), .D(n841), .Y(n447) );
  OAI22X1 U225 ( .A(n296), .B(n857), .C(n295), .D(n841), .Y(n448) );
  OAI22X1 U226 ( .A(n297), .B(n857), .C(n296), .D(n841), .Y(n449) );
  OAI22X1 U227 ( .A(n298), .B(n856), .C(n297), .D(n840), .Y(n450) );
  OAI22X1 U228 ( .A(n299), .B(n856), .C(n298), .D(n840), .Y(n451) );
  OAI22X1 U229 ( .A(n300), .B(n856), .C(n299), .D(n840), .Y(n452) );
  OAI22X1 U230 ( .A(n301), .B(n856), .C(n300), .D(n840), .Y(n453) );
  OAI22X1 U231 ( .A(n302), .B(n856), .C(n301), .D(n840), .Y(n454) );
  OAI22X1 U232 ( .A(n303), .B(n856), .C(n302), .D(n840), .Y(n455) );
  OAI22X1 U233 ( .A(n190), .B(n856), .C(n303), .D(n840), .Y(n456) );
  OAI22X1 U234 ( .A(n856), .B(n287), .C(n190), .D(n840), .Y(n542) );
  XNOR2X1 U235 ( .A(n871), .B(n831), .Y(n305) );
  XNOR2X1 U236 ( .A(n871), .B(n221), .Y(n306) );
  XNOR2X1 U237 ( .A(n871), .B(n222), .Y(n307) );
  XNOR2X1 U238 ( .A(n871), .B(n223), .Y(n308) );
  XNOR2X1 U239 ( .A(n871), .B(n224), .Y(n309) );
  XNOR2X1 U240 ( .A(n871), .B(n225), .Y(n310) );
  XNOR2X1 U241 ( .A(n871), .B(n226), .Y(n311) );
  XNOR2X1 U242 ( .A(n871), .B(n227), .Y(n312) );
  XNOR2X1 U243 ( .A(n870), .B(b[8]), .Y(n313) );
  XNOR2X1 U244 ( .A(n870), .B(b[9]), .Y(n314) );
  XNOR2X1 U245 ( .A(n870), .B(b[10]), .Y(n315) );
  XNOR2X1 U246 ( .A(n870), .B(b[11]), .Y(n316) );
  XNOR2X1 U247 ( .A(n870), .B(b[12]), .Y(n317) );
  XNOR2X1 U248 ( .A(n870), .B(b[13]), .Y(n318) );
  XNOR2X1 U249 ( .A(n870), .B(b[14]), .Y(n319) );
  XNOR2X1 U250 ( .A(n870), .B(b[15]), .Y(n320) );
  OAI22X1 U251 ( .A(n306), .B(n855), .C(n305), .D(n839), .Y(n459) );
  OAI22X1 U252 ( .A(n307), .B(n855), .C(n306), .D(n839), .Y(n460) );
  OAI22X1 U253 ( .A(n308), .B(n855), .C(n307), .D(n839), .Y(n461) );
  OAI22X1 U254 ( .A(n309), .B(n855), .C(n308), .D(n839), .Y(n462) );
  OAI22X1 U255 ( .A(n310), .B(n855), .C(n309), .D(n839), .Y(n463) );
  OAI22X1 U256 ( .A(n311), .B(n855), .C(n310), .D(n839), .Y(n464) );
  OAI22X1 U257 ( .A(n312), .B(n855), .C(n311), .D(n839), .Y(n465) );
  OAI22X1 U258 ( .A(n313), .B(n855), .C(n312), .D(n839), .Y(n466) );
  OAI22X1 U259 ( .A(n314), .B(n855), .C(n313), .D(n839), .Y(n467) );
  OAI22X1 U260 ( .A(n315), .B(n854), .C(n314), .D(n838), .Y(n468) );
  OAI22X1 U261 ( .A(n316), .B(n854), .C(n315), .D(n838), .Y(n469) );
  OAI22X1 U262 ( .A(n317), .B(n854), .C(n316), .D(n838), .Y(n470) );
  OAI22X1 U263 ( .A(n318), .B(n854), .C(n317), .D(n838), .Y(n471) );
  OAI22X1 U264 ( .A(n319), .B(n854), .C(n318), .D(n838), .Y(n472) );
  OAI22X1 U265 ( .A(n320), .B(n854), .C(n319), .D(n838), .Y(n473) );
  OAI22X1 U266 ( .A(n191), .B(n854), .C(n320), .D(n838), .Y(n474) );
  OAI22X1 U267 ( .A(n854), .B(n304), .C(n191), .D(n838), .Y(n543) );
  XNOR2X1 U268 ( .A(n869), .B(n831), .Y(n322) );
  XNOR2X1 U269 ( .A(n869), .B(n221), .Y(n323) );
  XNOR2X1 U270 ( .A(n869), .B(n222), .Y(n324) );
  XNOR2X1 U271 ( .A(n869), .B(n223), .Y(n325) );
  XNOR2X1 U272 ( .A(n869), .B(n224), .Y(n326) );
  XNOR2X1 U273 ( .A(n869), .B(n225), .Y(n327) );
  XNOR2X1 U274 ( .A(n869), .B(n226), .Y(n328) );
  XNOR2X1 U275 ( .A(n869), .B(n227), .Y(n329) );
  XNOR2X1 U276 ( .A(n868), .B(b[8]), .Y(n330) );
  XNOR2X1 U277 ( .A(n868), .B(b[9]), .Y(n331) );
  XNOR2X1 U278 ( .A(n868), .B(b[10]), .Y(n332) );
  XNOR2X1 U279 ( .A(n868), .B(b[11]), .Y(n333) );
  XNOR2X1 U280 ( .A(n868), .B(b[12]), .Y(n334) );
  XNOR2X1 U281 ( .A(n868), .B(b[13]), .Y(n335) );
  XNOR2X1 U282 ( .A(n868), .B(b[14]), .Y(n336) );
  XNOR2X1 U283 ( .A(n868), .B(b[15]), .Y(n337) );
  OAI22X1 U284 ( .A(n323), .B(n853), .C(n322), .D(n837), .Y(n477) );
  OAI22X1 U285 ( .A(n324), .B(n853), .C(n323), .D(n837), .Y(n478) );
  OAI22X1 U286 ( .A(n325), .B(n853), .C(n324), .D(n837), .Y(n479) );
  OAI22X1 U287 ( .A(n326), .B(n853), .C(n325), .D(n837), .Y(n480) );
  OAI22X1 U288 ( .A(n327), .B(n853), .C(n326), .D(n837), .Y(n481) );
  OAI22X1 U289 ( .A(n328), .B(n853), .C(n327), .D(n837), .Y(n482) );
  OAI22X1 U290 ( .A(n329), .B(n853), .C(n328), .D(n837), .Y(n483) );
  OAI22X1 U291 ( .A(n330), .B(n853), .C(n329), .D(n837), .Y(n484) );
  OAI22X1 U292 ( .A(n331), .B(n853), .C(n330), .D(n837), .Y(n485) );
  OAI22X1 U293 ( .A(n332), .B(n852), .C(n331), .D(n836), .Y(n486) );
  OAI22X1 U294 ( .A(n333), .B(n852), .C(n332), .D(n836), .Y(n487) );
  OAI22X1 U295 ( .A(n334), .B(n852), .C(n333), .D(n836), .Y(n488) );
  OAI22X1 U296 ( .A(n335), .B(n852), .C(n334), .D(n836), .Y(n489) );
  OAI22X1 U297 ( .A(n336), .B(n852), .C(n335), .D(n836), .Y(n490) );
  OAI22X1 U298 ( .A(n337), .B(n852), .C(n336), .D(n836), .Y(n491) );
  OAI22X1 U299 ( .A(n192), .B(n852), .C(n337), .D(n836), .Y(n492) );
  OAI22X1 U300 ( .A(n852), .B(n321), .C(n192), .D(n836), .Y(n544) );
  XNOR2X1 U301 ( .A(n867), .B(n831), .Y(n339) );
  XNOR2X1 U302 ( .A(n867), .B(n221), .Y(n340) );
  XNOR2X1 U303 ( .A(n867), .B(n222), .Y(n341) );
  XNOR2X1 U304 ( .A(n867), .B(n223), .Y(n342) );
  XNOR2X1 U305 ( .A(n867), .B(n224), .Y(n343) );
  XNOR2X1 U306 ( .A(n867), .B(n225), .Y(n344) );
  XNOR2X1 U307 ( .A(n867), .B(n226), .Y(n345) );
  XNOR2X1 U308 ( .A(n867), .B(n227), .Y(n346) );
  XNOR2X1 U309 ( .A(n866), .B(b[8]), .Y(n347) );
  XNOR2X1 U310 ( .A(n866), .B(b[9]), .Y(n348) );
  XNOR2X1 U311 ( .A(n866), .B(b[10]), .Y(n349) );
  XNOR2X1 U312 ( .A(n866), .B(b[11]), .Y(n350) );
  XNOR2X1 U313 ( .A(n866), .B(b[12]), .Y(n351) );
  XNOR2X1 U314 ( .A(n866), .B(b[13]), .Y(n352) );
  XNOR2X1 U315 ( .A(n866), .B(b[14]), .Y(n353) );
  XNOR2X1 U316 ( .A(n866), .B(b[15]), .Y(n354) );
  OAI22X1 U317 ( .A(n340), .B(n851), .C(n339), .D(n835), .Y(n495) );
  OAI22X1 U318 ( .A(n341), .B(n851), .C(n340), .D(n835), .Y(n496) );
  OAI22X1 U319 ( .A(n342), .B(n851), .C(n341), .D(n835), .Y(n497) );
  OAI22X1 U320 ( .A(n343), .B(n851), .C(n342), .D(n835), .Y(n498) );
  OAI22X1 U321 ( .A(n344), .B(n851), .C(n343), .D(n835), .Y(n499) );
  OAI22X1 U322 ( .A(n345), .B(n851), .C(n344), .D(n835), .Y(n500) );
  OAI22X1 U323 ( .A(n346), .B(n851), .C(n345), .D(n835), .Y(n501) );
  OAI22X1 U324 ( .A(n347), .B(n851), .C(n346), .D(n835), .Y(n502) );
  OAI22X1 U325 ( .A(n348), .B(n851), .C(n347), .D(n835), .Y(n503) );
  OAI22X1 U326 ( .A(n349), .B(n850), .C(n348), .D(n834), .Y(n504) );
  OAI22X1 U327 ( .A(n350), .B(n850), .C(n349), .D(n834), .Y(n505) );
  OAI22X1 U328 ( .A(n351), .B(n850), .C(n350), .D(n834), .Y(n506) );
  OAI22X1 U329 ( .A(n352), .B(n850), .C(n351), .D(n834), .Y(n507) );
  OAI22X1 U330 ( .A(n353), .B(n850), .C(n352), .D(n834), .Y(n508) );
  OAI22X1 U331 ( .A(n354), .B(n850), .C(n353), .D(n834), .Y(n509) );
  OAI22X1 U332 ( .A(n193), .B(n850), .C(n354), .D(n834), .Y(n510) );
  OAI22X1 U333 ( .A(n850), .B(n338), .C(n193), .D(n834), .Y(n545) );
  XNOR2X1 U334 ( .A(n865), .B(n831), .Y(n356) );
  XNOR2X1 U335 ( .A(n865), .B(n221), .Y(n357) );
  XNOR2X1 U336 ( .A(n865), .B(n222), .Y(n358) );
  XNOR2X1 U337 ( .A(n865), .B(n223), .Y(n359) );
  XNOR2X1 U338 ( .A(n865), .B(n224), .Y(n360) );
  XNOR2X1 U339 ( .A(n865), .B(n225), .Y(n361) );
  XNOR2X1 U340 ( .A(n865), .B(n226), .Y(n362) );
  XNOR2X1 U341 ( .A(n865), .B(n227), .Y(n363) );
  XNOR2X1 U342 ( .A(n864), .B(b[8]), .Y(n364) );
  XNOR2X1 U343 ( .A(n864), .B(b[9]), .Y(n365) );
  XNOR2X1 U344 ( .A(n864), .B(b[10]), .Y(n366) );
  XNOR2X1 U345 ( .A(n864), .B(b[11]), .Y(n367) );
  XNOR2X1 U346 ( .A(n864), .B(b[12]), .Y(n368) );
  XNOR2X1 U347 ( .A(n864), .B(b[13]), .Y(n369) );
  XNOR2X1 U348 ( .A(n864), .B(b[14]), .Y(n370) );
  XNOR2X1 U349 ( .A(n864), .B(b[15]), .Y(n371) );
  OAI22X1 U350 ( .A(n357), .B(n849), .C(n356), .D(n833), .Y(n513) );
  OAI22X1 U351 ( .A(n358), .B(n849), .C(n357), .D(n833), .Y(n514) );
  OAI22X1 U352 ( .A(n359), .B(n849), .C(n358), .D(n833), .Y(n515) );
  OAI22X1 U353 ( .A(n360), .B(n849), .C(n359), .D(n833), .Y(n516) );
  OAI22X1 U354 ( .A(n361), .B(n849), .C(n360), .D(n833), .Y(n517) );
  OAI22X1 U355 ( .A(n362), .B(n849), .C(n361), .D(n833), .Y(n518) );
  OAI22X1 U356 ( .A(n363), .B(n849), .C(n362), .D(n833), .Y(n519) );
  OAI22X1 U357 ( .A(n364), .B(n849), .C(n363), .D(n833), .Y(n520) );
  OAI22X1 U358 ( .A(n365), .B(n849), .C(n364), .D(n833), .Y(n521) );
  OAI22X1 U359 ( .A(n366), .B(n848), .C(n365), .D(n832), .Y(n522) );
  OAI22X1 U360 ( .A(n367), .B(n848), .C(n366), .D(n832), .Y(n523) );
  OAI22X1 U361 ( .A(n368), .B(n848), .C(n367), .D(n832), .Y(n524) );
  OAI22X1 U362 ( .A(n369), .B(n848), .C(n368), .D(n832), .Y(n525) );
  OAI22X1 U363 ( .A(n370), .B(n848), .C(n369), .D(n832), .Y(n526) );
  OAI22X1 U364 ( .A(n371), .B(n848), .C(n370), .D(n832), .Y(n527) );
  OAI22X1 U365 ( .A(n178), .B(n848), .C(n371), .D(n832), .Y(n528) );
  OAI22X1 U366 ( .A(n848), .B(n355), .C(n178), .D(n832), .Y(n546) );
  INVX2 U367 ( .A(n221), .Y(n372) );
  INVX2 U368 ( .A(n222), .Y(n373) );
  INVX2 U369 ( .A(n223), .Y(n374) );
  INVX2 U370 ( .A(n224), .Y(n375) );
  INVX2 U371 ( .A(n225), .Y(n376) );
  INVX2 U372 ( .A(n226), .Y(n377) );
  INVX2 U373 ( .A(n227), .Y(n378) );
  INVX2 U374 ( .A(b[8]), .Y(n379) );
  INVX2 U375 ( .A(b[9]), .Y(n380) );
  INVX2 U376 ( .A(b[10]), .Y(n381) );
  INVX2 U377 ( .A(b[11]), .Y(n382) );
  INVX2 U378 ( .A(b[12]), .Y(n383) );
  INVX2 U379 ( .A(b[13]), .Y(n384) );
  INVX2 U380 ( .A(b[14]), .Y(n385) );
  INVX2 U381 ( .A(b[15]), .Y(n386) );
  NOR2X1 U382 ( .A(n372), .B(n203), .Y(n675) );
  NOR2X1 U383 ( .A(n373), .B(n203), .Y(n531) );
  NOR2X1 U384 ( .A(n374), .B(n203), .Y(n532) );
  NOR2X1 U385 ( .A(n375), .B(n203), .Y(n705) );
  NOR2X1 U386 ( .A(n376), .B(n203), .Y(n533) );
  NOR2X1 U387 ( .A(n377), .B(n203), .Y(n731) );
  NOR2X1 U388 ( .A(n378), .B(n203), .Y(n534) );
  NOR2X1 U389 ( .A(n379), .B(n203), .Y(n753) );
  NOR2X1 U390 ( .A(n380), .B(n203), .Y(n535) );
  NOR2X1 U391 ( .A(n381), .B(n203), .Y(n771) );
  NOR2X1 U392 ( .A(n382), .B(n203), .Y(n536) );
  NOR2X1 U393 ( .A(n383), .B(n203), .Y(n785) );
  NOR2X1 U394 ( .A(n384), .B(n203), .Y(n537) );
  NOR2X1 U395 ( .A(n385), .B(n203), .Y(n795) );
  NOR2X1 U396 ( .A(n386), .B(n203), .Y(n538) );
  HAX1 U397 ( .A(n389), .B(n405), .YC(n548), .YS(n547) );
  FAX1 U398 ( .A(n390), .B(n406), .C(n548), .YC(n550), .YS(n549) );
  HAX1 U399 ( .A(n391), .B(n541), .YC(n552), .YS(n551) );
  FAX1 U400 ( .A(n407), .B(n423), .C(n551), .YC(n554), .YS(n553) );
  FAX1 U401 ( .A(n392), .B(n424), .C(n408), .YC(n556), .YS(n555) );
  FAX1 U402 ( .A(n552), .B(n943), .C(n555), .YC(n558), .YS(n557) );
  HAX1 U403 ( .A(n393), .B(n542), .YC(n560), .YS(n559) );
  FAX1 U404 ( .A(n409), .B(n441), .C(n425), .YC(n562), .YS(n561) );
  FAX1 U405 ( .A(n559), .B(n556), .C(n561), .YC(n564), .YS(n563) );
  FAX1 U406 ( .A(n394), .B(n426), .C(n442), .YC(n566), .YS(n565) );
  FAX1 U407 ( .A(n410), .B(n560), .C(n946), .YC(n568), .YS(n567) );
  FAX1 U408 ( .A(n562), .B(n565), .C(n567), .YC(n570), .YS(n569) );
  HAX1 U409 ( .A(n395), .B(n543), .YC(n572), .YS(n571) );
  FAX1 U410 ( .A(n443), .B(n459), .C(n427), .YC(n574), .YS(n573) );
  FAX1 U411 ( .A(n411), .B(n571), .C(n566), .YC(n576), .YS(n575) );
  FAX1 U412 ( .A(n573), .B(n568), .C(n575), .YC(n578), .YS(n577) );
  FAX1 U413 ( .A(n396), .B(n412), .C(n428), .YC(n580), .YS(n579) );
  FAX1 U414 ( .A(n444), .B(n460), .C(n572), .YC(n582), .YS(n581) );
  FAX1 U415 ( .A(n941), .B(n574), .C(n579), .YC(n584), .YS(n583) );
  FAX1 U416 ( .A(n581), .B(n576), .C(n583), .YC(n586), .YS(n585) );
  HAX1 U417 ( .A(n397), .B(n544), .YC(n588), .YS(n587) );
  FAX1 U418 ( .A(n445), .B(n477), .C(n413), .YC(n590), .YS(n589) );
  FAX1 U419 ( .A(n429), .B(n461), .C(n587), .YC(n592), .YS(n591) );
  FAX1 U420 ( .A(n580), .B(n589), .C(n582), .YC(n594), .YS(n593) );
  FAX1 U421 ( .A(n591), .B(n584), .C(n593), .YC(n596), .YS(n595) );
  FAX1 U422 ( .A(n398), .B(n414), .C(n478), .YC(n598), .YS(n597) );
  FAX1 U423 ( .A(n430), .B(n462), .C(n446), .YC(n600), .YS(n599) );
  FAX1 U424 ( .A(n588), .B(n942), .C(n590), .YC(n602), .YS(n601) );
  FAX1 U425 ( .A(n597), .B(n599), .C(n592), .YC(n604), .YS(n603) );
  FAX1 U426 ( .A(n601), .B(n594), .C(n603), .YC(n606), .YS(n605) );
  HAX1 U427 ( .A(n399), .B(n545), .YC(n608), .YS(n607) );
  FAX1 U428 ( .A(n463), .B(n415), .C(n431), .YC(n610), .YS(n609) );
  FAX1 U429 ( .A(n447), .B(n495), .C(n479), .YC(n612), .YS(n611) );
  FAX1 U430 ( .A(n607), .B(n598), .C(n600), .YC(n614), .YS(n613) );
  FAX1 U431 ( .A(n611), .B(n609), .C(n602), .YC(n616), .YS(n615) );
  FAX1 U432 ( .A(n613), .B(n604), .C(n615), .YC(n618), .YS(n617) );
  FAX1 U433 ( .A(n400), .B(n416), .C(n432), .YC(n620), .YS(n619) );
  FAX1 U434 ( .A(n448), .B(n496), .C(n480), .YC(n622), .YS(n621) );
  FAX1 U435 ( .A(n464), .B(n608), .C(n945), .YC(n624), .YS(n623) );
  FAX1 U436 ( .A(n610), .B(n612), .C(n619), .YC(n626), .YS(n625) );
  FAX1 U437 ( .A(n621), .B(n623), .C(n614), .YC(n628), .YS(n627) );
  FAX1 U438 ( .A(n625), .B(n616), .C(n627), .YC(n630), .YS(n629) );
  HAX1 U439 ( .A(n401), .B(n546), .YC(n632), .YS(n631) );
  FAX1 U440 ( .A(n465), .B(n513), .C(n497), .YC(n634), .YS(n633) );
  FAX1 U441 ( .A(n417), .B(n481), .C(n449), .YC(n636), .YS(n635) );
  FAX1 U442 ( .A(n433), .B(n631), .C(n620), .YC(n638), .YS(n637) );
  FAX1 U443 ( .A(n622), .B(n635), .C(n633), .YC(n640), .YS(n639) );
  FAX1 U444 ( .A(n624), .B(n626), .C(n637), .YC(n642), .YS(n641) );
  FAX1 U445 ( .A(n639), .B(n628), .C(n641), .YC(n644), .YS(n643) );
  FAX1 U446 ( .A(n402), .B(n418), .C(n947), .YC(n646), .YS(n645) );
  FAX1 U447 ( .A(n434), .B(n514), .C(n498), .YC(n648), .YS(n647) );
  FAX1 U448 ( .A(n450), .B(n482), .C(n466), .YC(n650), .YS(n649) );
  FAX1 U449 ( .A(n632), .B(n634), .C(n636), .YC(n652), .YS(n651) );
  FAX1 U450 ( .A(n645), .B(n649), .C(n647), .YC(n654), .YS(n653) );
  FAX1 U451 ( .A(n638), .B(n640), .C(n651), .YC(n656), .YS(n655) );
  FAX1 U452 ( .A(n653), .B(n642), .C(n655), .YC(n658), .YS(n657) );
  INVX2 U453 ( .A(n675), .Y(n659) );
  FAX1 U454 ( .A(n659), .B(n499), .C(n451), .YC(n661), .YS(n660) );
  FAX1 U455 ( .A(n467), .B(n483), .C(n515), .YC(n663), .YS(n662) );
  FAX1 U456 ( .A(n419), .B(n435), .C(n403), .YC(n665), .YS(n664) );
  FAX1 U457 ( .A(n646), .B(n648), .C(n650), .YC(n667), .YS(n666) );
  FAX1 U458 ( .A(n660), .B(n662), .C(n664), .YC(n669), .YS(n668) );
  FAX1 U459 ( .A(n652), .B(n654), .C(n666), .YC(n671), .YS(n670) );
  FAX1 U460 ( .A(n668), .B(n656), .C(n670), .YC(n673), .YS(n672) );
  FAX1 U462 ( .A(n531), .B(n659), .C(n420), .YC(n677), .YS(n676) );
  FAX1 U463 ( .A(n436), .B(n516), .C(n452), .YC(n679), .YS(n678) );
  FAX1 U464 ( .A(n468), .B(n500), .C(n484), .YC(n681), .YS(n680) );
  FAX1 U465 ( .A(n661), .B(n663), .C(n676), .YC(n683), .YS(n682) );
  FAX1 U466 ( .A(n680), .B(n678), .C(n665), .YC(n685), .YS(n684) );
  FAX1 U467 ( .A(n667), .B(n682), .C(n669), .YC(n687), .YS(n686) );
  FAX1 U468 ( .A(n684), .B(n671), .C(n686), .YC(n689), .YS(n688) );
  FAX1 U469 ( .A(n675), .B(n532), .C(n469), .YC(n691), .YS(n690) );
  FAX1 U470 ( .A(n485), .B(n501), .C(n517), .YC(n693), .YS(n692) );
  FAX1 U471 ( .A(n437), .B(n453), .C(n421), .YC(n695), .YS(n694) );
  FAX1 U472 ( .A(n677), .B(n679), .C(n681), .YC(n697), .YS(n696) );
  FAX1 U473 ( .A(n690), .B(n692), .C(n694), .YC(n699), .YS(n698) );
  FAX1 U474 ( .A(n683), .B(n696), .C(n685), .YC(n701), .YS(n700) );
  FAX1 U475 ( .A(n698), .B(n687), .C(n700), .YC(n703), .YS(n702) );
  INVX2 U476 ( .A(n705), .Y(n704) );
  FAX1 U477 ( .A(n704), .B(n438), .C(n454), .YC(n707), .YS(n706) );
  FAX1 U478 ( .A(n518), .B(n470), .C(n486), .YC(n709), .YS(n708) );
  FAX1 U479 ( .A(n502), .B(n691), .C(n693), .YC(n711), .YS(n710) );
  FAX1 U480 ( .A(n706), .B(n708), .C(n695), .YC(n713), .YS(n712) );
  FAX1 U481 ( .A(n697), .B(n710), .C(n699), .YC(n715), .YS(n714) );
  FAX1 U482 ( .A(n712), .B(n701), .C(n714), .YC(n717), .YS(n716) );
  FAX1 U483 ( .A(n705), .B(n533), .C(n471), .YC(n719), .YS(n718) );
  FAX1 U484 ( .A(n487), .B(n519), .C(n455), .YC(n721), .YS(n720) );
  FAX1 U485 ( .A(n503), .B(n439), .C(n707), .YC(n723), .YS(n722) );
  FAX1 U486 ( .A(n709), .B(n718), .C(n720), .YC(n725), .YS(n724) );
  FAX1 U487 ( .A(n711), .B(n722), .C(n713), .YC(n727), .YS(n726) );
  FAX1 U488 ( .A(n724), .B(n715), .C(n726), .YC(n729), .YS(n728) );
  INVX2 U489 ( .A(n731), .Y(n730) );
  FAX1 U490 ( .A(n730), .B(n456), .C(n472), .YC(n733), .YS(n732) );
  FAX1 U491 ( .A(n520), .B(n504), .C(n488), .YC(n735), .YS(n734) );
  FAX1 U492 ( .A(n719), .B(n721), .C(n732), .YC(n737), .YS(n736) );
  FAX1 U493 ( .A(n734), .B(n723), .C(n725), .YC(n739), .YS(n738) );
  FAX1 U494 ( .A(n736), .B(n727), .C(n738), .YC(n741), .YS(n740) );
  FAX1 U495 ( .A(n731), .B(n534), .C(n489), .YC(n743), .YS(n742) );
  FAX1 U496 ( .A(n505), .B(n521), .C(n473), .YC(n745), .YS(n744) );
  FAX1 U497 ( .A(n457), .B(n733), .C(n735), .YC(n747), .YS(n746) );
  FAX1 U498 ( .A(n742), .B(n744), .C(n737), .YC(n749), .YS(n748) );
  FAX1 U499 ( .A(n746), .B(n739), .C(n748), .YC(n751), .YS(n750) );
  INVX2 U500 ( .A(n753), .Y(n752) );
  FAX1 U501 ( .A(n752), .B(n474), .C(n490), .YC(n755), .YS(n754) );
  FAX1 U502 ( .A(n506), .B(n522), .C(n743), .YC(n757), .YS(n756) );
  FAX1 U503 ( .A(n745), .B(n754), .C(n756), .YC(n759), .YS(n758) );
  FAX1 U504 ( .A(n747), .B(n749), .C(n758), .YC(n761), .YS(n760) );
  FAX1 U505 ( .A(n753), .B(n535), .C(n491), .YC(n763), .YS(n762) );
  FAX1 U506 ( .A(n523), .B(n507), .C(n475), .YC(n765), .YS(n764) );
  FAX1 U507 ( .A(n755), .B(n762), .C(n764), .YC(n767), .YS(n766) );
  FAX1 U508 ( .A(n757), .B(n766), .C(n759), .YC(n769), .YS(n768) );
  INVX2 U509 ( .A(n771), .Y(n770) );
  FAX1 U510 ( .A(n770), .B(n492), .C(n508), .YC(n773), .YS(n772) );
  FAX1 U511 ( .A(n524), .B(n763), .C(n772), .YC(n775), .YS(n774) );
  FAX1 U512 ( .A(n765), .B(n774), .C(n767), .YC(n777), .YS(n776) );
  FAX1 U513 ( .A(n771), .B(n536), .C(n509), .YC(n779), .YS(n778) );
  FAX1 U514 ( .A(n525), .B(n493), .C(n773), .YC(n781), .YS(n780) );
  FAX1 U515 ( .A(n778), .B(n775), .C(n780), .YC(n783), .YS(n782) );
  INVX2 U516 ( .A(n785), .Y(n784) );
  FAX1 U517 ( .A(n784), .B(n510), .C(n526), .YC(n787), .YS(n786) );
  FAX1 U518 ( .A(n779), .B(n786), .C(n781), .YC(n789), .YS(n788) );
  FAX1 U519 ( .A(n785), .B(n537), .C(n527), .YC(n791), .YS(n790) );
  FAX1 U520 ( .A(n511), .B(n787), .C(n790), .YC(n793), .YS(n792) );
  INVX2 U521 ( .A(n795), .Y(n794) );
  FAX1 U522 ( .A(n794), .B(n528), .C(n791), .YC(n797), .YS(n796) );
  HAX1 U523 ( .A(n539), .B(n387), .YC(n799), .YS(product[1]) );
  FAX1 U524 ( .A(n388), .B(n799), .C(n944), .YC(n800), .YS(product[2]) );
  FAX1 U525 ( .A(n540), .B(n547), .C(n800), .YC(n801), .YS(product[3]) );
  FAX1 U526 ( .A(n940), .B(n549), .C(n801), .YC(n802), .YS(product[4]) );
  FAX1 U527 ( .A(n550), .B(n553), .C(n802), .YC(n803), .YS(product[5]) );
  FAX1 U528 ( .A(n554), .B(n557), .C(n803), .YC(n804), .YS(product[6]) );
  FAX1 U529 ( .A(n558), .B(n563), .C(n804), .YC(n805), .YS(product[7]) );
  FAX1 U530 ( .A(n564), .B(n569), .C(n805), .YC(n806), .YS(product[8]) );
  FAX1 U531 ( .A(n570), .B(n577), .C(n806), .YC(n807), .YS(product[9]) );
  FAX1 U532 ( .A(n578), .B(n585), .C(n807), .YC(n808), .YS(product[10]) );
  FAX1 U533 ( .A(n586), .B(n595), .C(n808), .YC(n809), .YS(product[11]) );
  FAX1 U534 ( .A(n596), .B(n605), .C(n809), .YC(n810), .YS(product[12]) );
  FAX1 U535 ( .A(n606), .B(n617), .C(n810), .YC(n811), .YS(product[13]) );
  FAX1 U536 ( .A(n618), .B(n629), .C(n811), .YC(n812), .YS(product[14]) );
  FAX1 U537 ( .A(n630), .B(n643), .C(n812), .YC(n813), .YS(product[15]) );
  FAX1 U538 ( .A(n644), .B(n657), .C(n813), .YC(n814), .YS(product[16]) );
  FAX1 U539 ( .A(n658), .B(n672), .C(n814), .YC(n815), .YS(product[17]) );
  FAX1 U540 ( .A(n673), .B(n688), .C(n815), .YC(n816), .YS(product[18]) );
  FAX1 U541 ( .A(n689), .B(n702), .C(n816), .YC(n817), .YS(product[19]) );
  FAX1 U542 ( .A(n703), .B(n716), .C(n817), .YC(n818), .YS(product[20]) );
  FAX1 U543 ( .A(n717), .B(n728), .C(n818), .YC(n819), .YS(product[21]) );
  FAX1 U544 ( .A(n729), .B(n740), .C(n819), .YC(n820), .YS(product[22]) );
  FAX1 U545 ( .A(n741), .B(n750), .C(n820), .YC(n821), .YS(product[23]) );
  FAX1 U546 ( .A(n751), .B(n760), .C(n821), .YC(n822), .YS(product[24]) );
  FAX1 U547 ( .A(n761), .B(n768), .C(n822), .YC(n823), .YS(product[25]) );
  FAX1 U548 ( .A(n776), .B(n769), .C(n823), .YC(n824), .YS(product[26]) );
  FAX1 U549 ( .A(n782), .B(n777), .C(n824), .YC(n825), .YS(product[27]) );
  FAX1 U550 ( .A(n788), .B(n783), .C(n825), .YC(n826), .YS(product[28]) );
  FAX1 U551 ( .A(n792), .B(n789), .C(n826), .YC(n827), .YS(product[29]) );
  FAX1 U552 ( .A(n796), .B(n793), .C(n827), .YC(n828), .YS(product[30]) );
  XOR2X1 U553 ( .A(n797), .B(n798), .Y(n829) );
  XOR2X1 U554 ( .A(n828), .B(n829), .Y(product[31]) );
  AND2X2 U607 ( .A(n831), .B(a[0]), .Y(product[0]) );
  AND2X2 U608 ( .A(n830), .B(n134), .Y(n940) );
  AND2X2 U609 ( .A(n830), .B(n86), .Y(n941) );
  AND2X2 U610 ( .A(n830), .B(n60), .Y(n942) );
  AND2X2 U611 ( .A(n830), .B(n118), .Y(n943) );
  AND2X2 U612 ( .A(n831), .B(n150), .Y(n944) );
  AND2X2 U613 ( .A(n830), .B(n26), .Y(n945) );
  AND2X2 U614 ( .A(n830), .B(n102), .Y(n946) );
  AND2X2 U615 ( .A(n830), .B(a[15]), .Y(n947) );
  BUFX2 U616 ( .A(n205), .Y(n845) );
  BUFX2 U617 ( .A(n206), .Y(n843) );
  BUFX2 U618 ( .A(n207), .Y(n841) );
  BUFX2 U619 ( .A(n208), .Y(n839) );
  BUFX2 U620 ( .A(n209), .Y(n837) );
  BUFX2 U621 ( .A(n210), .Y(n835) );
  BUFX2 U622 ( .A(n211), .Y(n833) );
  BUFX2 U623 ( .A(n204), .Y(n847) );
  BUFX2 U624 ( .A(n196), .Y(n861) );
  BUFX2 U625 ( .A(n197), .Y(n859) );
  BUFX2 U626 ( .A(n198), .Y(n857) );
  BUFX2 U627 ( .A(n199), .Y(n855) );
  BUFX2 U628 ( .A(n200), .Y(n853) );
  BUFX2 U629 ( .A(n201), .Y(n851) );
  BUFX2 U630 ( .A(n202), .Y(n849) );
  BUFX2 U631 ( .A(n196), .Y(n860) );
  BUFX2 U632 ( .A(n197), .Y(n858) );
  BUFX2 U633 ( .A(n198), .Y(n856) );
  BUFX2 U634 ( .A(n199), .Y(n854) );
  BUFX2 U635 ( .A(n200), .Y(n852) );
  BUFX2 U636 ( .A(n201), .Y(n850) );
  BUFX2 U637 ( .A(n202), .Y(n848) );
  BUFX2 U638 ( .A(n195), .Y(n862) );
  BUFX2 U639 ( .A(n205), .Y(n844) );
  BUFX2 U640 ( .A(n206), .Y(n842) );
  BUFX2 U641 ( .A(n207), .Y(n840) );
  BUFX2 U642 ( .A(n208), .Y(n838) );
  BUFX2 U643 ( .A(n209), .Y(n836) );
  BUFX2 U644 ( .A(n211), .Y(n832) );
  BUFX2 U645 ( .A(n210), .Y(n834) );
  BUFX2 U646 ( .A(n204), .Y(n846) );
  BUFX2 U647 ( .A(n195), .Y(n863) );
  BUFX2 U648 ( .A(b[0]), .Y(n831) );
  BUFX2 U649 ( .A(a[1]), .Y(n879) );
  BUFX2 U650 ( .A(a[5]), .Y(n875) );
  BUFX2 U651 ( .A(a[3]), .Y(n877) );
  BUFX2 U652 ( .A(a[7]), .Y(n873) );
  BUFX2 U653 ( .A(a[9]), .Y(n871) );
  BUFX2 U654 ( .A(a[11]), .Y(n869) );
  BUFX2 U655 ( .A(a[13]), .Y(n867) );
  BUFX2 U656 ( .A(a[15]), .Y(n865) );
  BUFX2 U657 ( .A(a[1]), .Y(n878) );
  BUFX2 U658 ( .A(a[3]), .Y(n876) );
  BUFX2 U659 ( .A(a[5]), .Y(n874) );
  BUFX2 U660 ( .A(a[7]), .Y(n872) );
  BUFX2 U661 ( .A(a[9]), .Y(n870) );
  BUFX2 U662 ( .A(a[11]), .Y(n868) );
  BUFX2 U663 ( .A(a[13]), .Y(n866) );
  BUFX2 U664 ( .A(a[15]), .Y(n864) );
  BUFX2 U665 ( .A(n178), .Y(n203) );
  BUFX2 U666 ( .A(b[0]), .Y(n830) );
  BUFX2 U667 ( .A(b[1]), .Y(n221) );
  BUFX2 U668 ( .A(b[2]), .Y(n222) );
  BUFX2 U669 ( .A(b[3]), .Y(n223) );
  BUFX2 U670 ( .A(b[4]), .Y(n224) );
  BUFX2 U671 ( .A(b[5]), .Y(n225) );
  BUFX2 U672 ( .A(b[6]), .Y(n226) );
  BUFX2 U673 ( .A(b[7]), .Y(n227) );
endmodule


module alu_DW_mult_uns_8 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n15, n25, n26, n50, n60, n80, n85, n86, n101, n102, n117, n118, n133,
         n134, n149, n150, n160, n165, n176, n178, n187, n188, n189, n190,
         n191, n192, n193, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n940, n941, n942, n943,
         n944, n945, n946, n947;

  NAND2X1 OR_NOTi ( .A(n176), .B(n878), .Y(n236) );
  INVX1 U1 ( .A(n831), .Y(n176) );
  OAI21X1 AO21i ( .A(n165), .B(a[0]), .C(a[1]), .Y(n403) );
  INVX1 U12 ( .A(n846), .Y(n165) );
  NAND2X1 OR_NOTi1 ( .A(n160), .B(n876), .Y(n253) );
  INVX1 U13 ( .A(n831), .Y(n160) );
  OAI21X1 AO21i1 ( .A(n149), .B(n150), .C(a[3]), .Y(n421) );
  INVX1 U23 ( .A(n860), .Y(n150) );
  INVX1 U15 ( .A(n844), .Y(n149) );
  NAND2X1 OR_NOTi2 ( .A(n160), .B(n874), .Y(n270) );
  OAI21X1 AO21i2 ( .A(n133), .B(n134), .C(a[5]), .Y(n439) );
  INVX1 U25 ( .A(n858), .Y(n134) );
  INVX1 U18 ( .A(n842), .Y(n133) );
  NAND2X1 OR_NOTi3 ( .A(n160), .B(n872), .Y(n287) );
  OAI21X1 AO21i3 ( .A(n117), .B(n118), .C(a[7]), .Y(n457) );
  INVX1 U27 ( .A(n856), .Y(n118) );
  INVX1 U111 ( .A(n840), .Y(n117) );
  NAND2X1 OR_NOTi4 ( .A(n80), .B(n870), .Y(n304) );
  OAI21X1 AO21i4 ( .A(n101), .B(n102), .C(a[9]), .Y(n475) );
  INVX1 U29 ( .A(n854), .Y(n102) );
  INVX1 U114 ( .A(n838), .Y(n101) );
  NAND2X1 OR_NOTi5 ( .A(n80), .B(n868), .Y(n321) );
  OAI21X1 AO21i5 ( .A(n85), .B(n86), .C(a[11]), .Y(n493) );
  INVX1 U211 ( .A(n852), .Y(n86) );
  INVX1 U117 ( .A(n836), .Y(n85) );
  NAND2X1 OR_NOTi6 ( .A(n80), .B(n866), .Y(n338) );
  INVX1 U118 ( .A(n830), .Y(n80) );
  OAI21X1 AO21i6 ( .A(n50), .B(n60), .C(a[13]), .Y(n511) );
  INVX1 U213 ( .A(n850), .Y(n60) );
  INVX1 U120 ( .A(n834), .Y(n50) );
  NAND2X1 OR_NOTi7 ( .A(n176), .B(n864), .Y(n355) );
  OAI21X1 AO21i7 ( .A(n25), .B(n26), .C(a[15]), .Y(n529) );
  INVX1 U215 ( .A(n848), .Y(n26) );
  INVX1 U123 ( .A(n832), .Y(n25) );
  XOR2X1 U217 ( .A(n538), .B(n795), .Y(n15) );
  XOR2X1 U125 ( .A(n529), .B(n15), .Y(n798) );
  INVX2 U4 ( .A(a[0]), .Y(n195) );
  XOR2X1 U5 ( .A(a[0]), .B(a[1]), .Y(n212) );
  NAND2X1 U6 ( .A(n195), .B(n212), .Y(n204) );
  XNOR2X1 U7 ( .A(a[2]), .B(a[1]), .Y(n196) );
  XOR2X1 U8 ( .A(a[2]), .B(a[3]), .Y(n213) );
  NAND2X1 U9 ( .A(n213), .B(n196), .Y(n205) );
  XNOR2X1 U10 ( .A(a[4]), .B(a[3]), .Y(n197) );
  XOR2X1 U20 ( .A(a[4]), .B(a[5]), .Y(n214) );
  NAND2X1 U30 ( .A(n214), .B(n197), .Y(n206) );
  XNOR2X1 U38 ( .A(a[6]), .B(a[5]), .Y(n198) );
  XOR2X1 U39 ( .A(a[6]), .B(a[7]), .Y(n215) );
  NAND2X1 U40 ( .A(n215), .B(n198), .Y(n207) );
  XNOR2X1 U41 ( .A(a[8]), .B(a[7]), .Y(n199) );
  XOR2X1 U42 ( .A(a[8]), .B(a[9]), .Y(n216) );
  NAND2X1 U43 ( .A(n216), .B(n199), .Y(n208) );
  XNOR2X1 U44 ( .A(a[10]), .B(a[9]), .Y(n200) );
  XOR2X1 U45 ( .A(a[10]), .B(a[11]), .Y(n217) );
  NAND2X1 U46 ( .A(n217), .B(n200), .Y(n209) );
  XNOR2X1 U47 ( .A(a[12]), .B(a[11]), .Y(n201) );
  XOR2X1 U48 ( .A(a[12]), .B(a[13]), .Y(n218) );
  NAND2X1 U49 ( .A(n218), .B(n201), .Y(n210) );
  XNOR2X1 U50 ( .A(a[14]), .B(a[13]), .Y(n202) );
  XOR2X1 U51 ( .A(a[14]), .B(a[15]), .Y(n219) );
  NAND2X1 U52 ( .A(n219), .B(n202), .Y(n211) );
  INVX2 U53 ( .A(a[15]), .Y(n178) );
  INVX2 U54 ( .A(n879), .Y(n187) );
  INVX2 U55 ( .A(n877), .Y(n188) );
  INVX2 U56 ( .A(n875), .Y(n189) );
  INVX2 U57 ( .A(n873), .Y(n190) );
  INVX2 U58 ( .A(n871), .Y(n191) );
  INVX2 U59 ( .A(n869), .Y(n192) );
  INVX2 U60 ( .A(n867), .Y(n193) );
  XNOR2X1 U78 ( .A(n879), .B(n831), .Y(n237) );
  XNOR2X1 U79 ( .A(n879), .B(n221), .Y(n238) );
  XNOR2X1 U80 ( .A(n879), .B(n222), .Y(n239) );
  XNOR2X1 U81 ( .A(n879), .B(n223), .Y(n240) );
  XNOR2X1 U82 ( .A(n879), .B(n224), .Y(n241) );
  XNOR2X1 U83 ( .A(n879), .B(n225), .Y(n242) );
  XNOR2X1 U84 ( .A(n879), .B(n226), .Y(n243) );
  XNOR2X1 U85 ( .A(n879), .B(n227), .Y(n244) );
  XNOR2X1 U86 ( .A(n878), .B(n228), .Y(n245) );
  XNOR2X1 U87 ( .A(n878), .B(n229), .Y(n246) );
  XNOR2X1 U88 ( .A(n878), .B(n230), .Y(n247) );
  XNOR2X1 U89 ( .A(n878), .B(n231), .Y(n248) );
  XNOR2X1 U90 ( .A(n878), .B(n232), .Y(n249) );
  XNOR2X1 U91 ( .A(n878), .B(n233), .Y(n250) );
  XNOR2X1 U92 ( .A(n878), .B(n234), .Y(n251) );
  XNOR2X1 U93 ( .A(n878), .B(n235), .Y(n252) );
  OAI22X1 U94 ( .A(n863), .B(n238), .C(n237), .D(n847), .Y(n387) );
  OAI22X1 U95 ( .A(n863), .B(n239), .C(n238), .D(n847), .Y(n388) );
  OAI22X1 U96 ( .A(n863), .B(n240), .C(n239), .D(n847), .Y(n389) );
  OAI22X1 U97 ( .A(n863), .B(n241), .C(n240), .D(n847), .Y(n390) );
  OAI22X1 U98 ( .A(n863), .B(n242), .C(n241), .D(n847), .Y(n391) );
  OAI22X1 U99 ( .A(n863), .B(n243), .C(n242), .D(n847), .Y(n392) );
  OAI22X1 U100 ( .A(n863), .B(n244), .C(n243), .D(n847), .Y(n393) );
  OAI22X1 U101 ( .A(n863), .B(n245), .C(n244), .D(n847), .Y(n394) );
  OAI22X1 U102 ( .A(n863), .B(n246), .C(n245), .D(n847), .Y(n395) );
  OAI22X1 U103 ( .A(n862), .B(n247), .C(n246), .D(n846), .Y(n396) );
  OAI22X1 U104 ( .A(n862), .B(n248), .C(n247), .D(n846), .Y(n397) );
  OAI22X1 U105 ( .A(n862), .B(n249), .C(n248), .D(n846), .Y(n398) );
  OAI22X1 U106 ( .A(n862), .B(n250), .C(n249), .D(n846), .Y(n399) );
  OAI22X1 U107 ( .A(n862), .B(n251), .C(n250), .D(n846), .Y(n400) );
  OAI22X1 U108 ( .A(n862), .B(n252), .C(n251), .D(n846), .Y(n401) );
  OAI22X1 U109 ( .A(n862), .B(n187), .C(n252), .D(n846), .Y(n402) );
  OAI22X1 U127 ( .A(n862), .B(n236), .C(n187), .D(n846), .Y(n539) );
  XNOR2X1 U128 ( .A(n877), .B(n831), .Y(n254) );
  XNOR2X1 U129 ( .A(n877), .B(n221), .Y(n255) );
  XNOR2X1 U130 ( .A(n877), .B(n222), .Y(n256) );
  XNOR2X1 U131 ( .A(n877), .B(n223), .Y(n257) );
  XNOR2X1 U132 ( .A(n877), .B(n224), .Y(n258) );
  XNOR2X1 U133 ( .A(n877), .B(n225), .Y(n259) );
  XNOR2X1 U134 ( .A(n877), .B(n226), .Y(n260) );
  XNOR2X1 U135 ( .A(n877), .B(n227), .Y(n261) );
  XNOR2X1 U136 ( .A(n876), .B(n228), .Y(n262) );
  XNOR2X1 U137 ( .A(n876), .B(n229), .Y(n263) );
  XNOR2X1 U138 ( .A(n876), .B(n230), .Y(n264) );
  XNOR2X1 U139 ( .A(n876), .B(n231), .Y(n265) );
  XNOR2X1 U140 ( .A(n876), .B(n232), .Y(n266) );
  XNOR2X1 U141 ( .A(n876), .B(n233), .Y(n267) );
  XNOR2X1 U142 ( .A(n876), .B(n234), .Y(n268) );
  XNOR2X1 U143 ( .A(n876), .B(n235), .Y(n269) );
  OAI22X1 U144 ( .A(n255), .B(n861), .C(n254), .D(n845), .Y(n405) );
  OAI22X1 U145 ( .A(n256), .B(n861), .C(n255), .D(n845), .Y(n406) );
  OAI22X1 U146 ( .A(n257), .B(n861), .C(n256), .D(n845), .Y(n407) );
  OAI22X1 U147 ( .A(n258), .B(n861), .C(n257), .D(n845), .Y(n408) );
  OAI22X1 U148 ( .A(n259), .B(n861), .C(n258), .D(n845), .Y(n409) );
  OAI22X1 U149 ( .A(n260), .B(n861), .C(n259), .D(n845), .Y(n410) );
  OAI22X1 U150 ( .A(n261), .B(n861), .C(n260), .D(n845), .Y(n411) );
  OAI22X1 U151 ( .A(n262), .B(n861), .C(n261), .D(n845), .Y(n412) );
  OAI22X1 U152 ( .A(n263), .B(n861), .C(n262), .D(n845), .Y(n413) );
  OAI22X1 U153 ( .A(n264), .B(n860), .C(n263), .D(n844), .Y(n414) );
  OAI22X1 U154 ( .A(n265), .B(n860), .C(n264), .D(n844), .Y(n415) );
  OAI22X1 U155 ( .A(n266), .B(n860), .C(n265), .D(n844), .Y(n416) );
  OAI22X1 U156 ( .A(n267), .B(n860), .C(n266), .D(n844), .Y(n417) );
  OAI22X1 U157 ( .A(n268), .B(n860), .C(n267), .D(n844), .Y(n418) );
  OAI22X1 U158 ( .A(n269), .B(n860), .C(n268), .D(n844), .Y(n419) );
  OAI22X1 U159 ( .A(n188), .B(n860), .C(n269), .D(n844), .Y(n420) );
  OAI22X1 U160 ( .A(n860), .B(n253), .C(n188), .D(n844), .Y(n540) );
  XNOR2X1 U161 ( .A(n875), .B(n831), .Y(n271) );
  XNOR2X1 U162 ( .A(n875), .B(n221), .Y(n272) );
  XNOR2X1 U163 ( .A(n875), .B(n222), .Y(n273) );
  XNOR2X1 U164 ( .A(n875), .B(n223), .Y(n274) );
  XNOR2X1 U165 ( .A(n875), .B(n224), .Y(n275) );
  XNOR2X1 U166 ( .A(n875), .B(n225), .Y(n276) );
  XNOR2X1 U167 ( .A(n875), .B(n226), .Y(n277) );
  XNOR2X1 U168 ( .A(n875), .B(n227), .Y(n278) );
  XNOR2X1 U169 ( .A(n874), .B(n228), .Y(n279) );
  XNOR2X1 U170 ( .A(n874), .B(n229), .Y(n280) );
  XNOR2X1 U171 ( .A(n874), .B(n230), .Y(n281) );
  XNOR2X1 U172 ( .A(n874), .B(n231), .Y(n282) );
  XNOR2X1 U173 ( .A(n874), .B(n232), .Y(n283) );
  XNOR2X1 U174 ( .A(n874), .B(n233), .Y(n284) );
  XNOR2X1 U175 ( .A(n874), .B(n234), .Y(n285) );
  XNOR2X1 U176 ( .A(n874), .B(n235), .Y(n286) );
  OAI22X1 U177 ( .A(n272), .B(n859), .C(n271), .D(n843), .Y(n423) );
  OAI22X1 U178 ( .A(n273), .B(n859), .C(n272), .D(n843), .Y(n424) );
  OAI22X1 U179 ( .A(n274), .B(n859), .C(n273), .D(n843), .Y(n425) );
  OAI22X1 U180 ( .A(n275), .B(n859), .C(n274), .D(n843), .Y(n426) );
  OAI22X1 U181 ( .A(n276), .B(n859), .C(n275), .D(n843), .Y(n427) );
  OAI22X1 U182 ( .A(n277), .B(n859), .C(n276), .D(n843), .Y(n428) );
  OAI22X1 U183 ( .A(n278), .B(n859), .C(n277), .D(n843), .Y(n429) );
  OAI22X1 U184 ( .A(n279), .B(n859), .C(n278), .D(n843), .Y(n430) );
  OAI22X1 U185 ( .A(n280), .B(n859), .C(n279), .D(n843), .Y(n431) );
  OAI22X1 U186 ( .A(n281), .B(n858), .C(n280), .D(n842), .Y(n432) );
  OAI22X1 U187 ( .A(n282), .B(n858), .C(n281), .D(n842), .Y(n433) );
  OAI22X1 U188 ( .A(n283), .B(n858), .C(n282), .D(n842), .Y(n434) );
  OAI22X1 U189 ( .A(n284), .B(n858), .C(n283), .D(n842), .Y(n435) );
  OAI22X1 U190 ( .A(n285), .B(n858), .C(n284), .D(n842), .Y(n436) );
  OAI22X1 U191 ( .A(n286), .B(n858), .C(n285), .D(n842), .Y(n437) );
  OAI22X1 U192 ( .A(n189), .B(n858), .C(n286), .D(n842), .Y(n438) );
  OAI22X1 U193 ( .A(n858), .B(n270), .C(n189), .D(n842), .Y(n541) );
  XNOR2X1 U194 ( .A(n873), .B(n831), .Y(n288) );
  XNOR2X1 U195 ( .A(n873), .B(n221), .Y(n289) );
  XNOR2X1 U196 ( .A(n873), .B(n222), .Y(n290) );
  XNOR2X1 U197 ( .A(n873), .B(n223), .Y(n291) );
  XNOR2X1 U198 ( .A(n873), .B(n224), .Y(n292) );
  XNOR2X1 U199 ( .A(n873), .B(n225), .Y(n293) );
  XNOR2X1 U200 ( .A(n873), .B(n226), .Y(n294) );
  XNOR2X1 U201 ( .A(n873), .B(n227), .Y(n295) );
  XNOR2X1 U202 ( .A(n872), .B(n228), .Y(n296) );
  XNOR2X1 U203 ( .A(n872), .B(n229), .Y(n297) );
  XNOR2X1 U204 ( .A(n872), .B(n230), .Y(n298) );
  XNOR2X1 U205 ( .A(n872), .B(n231), .Y(n299) );
  XNOR2X1 U206 ( .A(n872), .B(n232), .Y(n300) );
  XNOR2X1 U207 ( .A(n872), .B(n233), .Y(n301) );
  XNOR2X1 U208 ( .A(n872), .B(n234), .Y(n302) );
  XNOR2X1 U209 ( .A(n872), .B(n235), .Y(n303) );
  OAI22X1 U218 ( .A(n289), .B(n857), .C(n288), .D(n841), .Y(n441) );
  OAI22X1 U219 ( .A(n290), .B(n857), .C(n289), .D(n841), .Y(n442) );
  OAI22X1 U220 ( .A(n291), .B(n857), .C(n290), .D(n841), .Y(n443) );
  OAI22X1 U221 ( .A(n292), .B(n857), .C(n291), .D(n841), .Y(n444) );
  OAI22X1 U222 ( .A(n293), .B(n857), .C(n292), .D(n841), .Y(n445) );
  OAI22X1 U223 ( .A(n294), .B(n857), .C(n293), .D(n841), .Y(n446) );
  OAI22X1 U224 ( .A(n295), .B(n857), .C(n294), .D(n841), .Y(n447) );
  OAI22X1 U225 ( .A(n296), .B(n857), .C(n295), .D(n841), .Y(n448) );
  OAI22X1 U226 ( .A(n297), .B(n857), .C(n296), .D(n841), .Y(n449) );
  OAI22X1 U227 ( .A(n298), .B(n856), .C(n297), .D(n840), .Y(n450) );
  OAI22X1 U228 ( .A(n299), .B(n856), .C(n298), .D(n840), .Y(n451) );
  OAI22X1 U229 ( .A(n300), .B(n856), .C(n299), .D(n840), .Y(n452) );
  OAI22X1 U230 ( .A(n301), .B(n856), .C(n300), .D(n840), .Y(n453) );
  OAI22X1 U231 ( .A(n302), .B(n856), .C(n301), .D(n840), .Y(n454) );
  OAI22X1 U232 ( .A(n303), .B(n856), .C(n302), .D(n840), .Y(n455) );
  OAI22X1 U233 ( .A(n190), .B(n856), .C(n303), .D(n840), .Y(n456) );
  OAI22X1 U234 ( .A(n856), .B(n287), .C(n190), .D(n840), .Y(n542) );
  XNOR2X1 U235 ( .A(n871), .B(n831), .Y(n305) );
  XNOR2X1 U236 ( .A(n871), .B(n221), .Y(n306) );
  XNOR2X1 U237 ( .A(n871), .B(n222), .Y(n307) );
  XNOR2X1 U238 ( .A(n871), .B(n223), .Y(n308) );
  XNOR2X1 U239 ( .A(n871), .B(n224), .Y(n309) );
  XNOR2X1 U240 ( .A(n871), .B(n225), .Y(n310) );
  XNOR2X1 U241 ( .A(n871), .B(n226), .Y(n311) );
  XNOR2X1 U242 ( .A(n871), .B(n227), .Y(n312) );
  XNOR2X1 U243 ( .A(n870), .B(n228), .Y(n313) );
  XNOR2X1 U244 ( .A(n870), .B(n229), .Y(n314) );
  XNOR2X1 U245 ( .A(n870), .B(n230), .Y(n315) );
  XNOR2X1 U246 ( .A(n870), .B(n231), .Y(n316) );
  XNOR2X1 U247 ( .A(n870), .B(n232), .Y(n317) );
  XNOR2X1 U248 ( .A(n870), .B(n233), .Y(n318) );
  XNOR2X1 U249 ( .A(n870), .B(n234), .Y(n319) );
  XNOR2X1 U250 ( .A(n870), .B(n235), .Y(n320) );
  OAI22X1 U251 ( .A(n306), .B(n855), .C(n305), .D(n839), .Y(n459) );
  OAI22X1 U252 ( .A(n307), .B(n855), .C(n306), .D(n839), .Y(n460) );
  OAI22X1 U253 ( .A(n308), .B(n855), .C(n307), .D(n839), .Y(n461) );
  OAI22X1 U254 ( .A(n309), .B(n855), .C(n308), .D(n839), .Y(n462) );
  OAI22X1 U255 ( .A(n310), .B(n855), .C(n309), .D(n839), .Y(n463) );
  OAI22X1 U256 ( .A(n311), .B(n855), .C(n310), .D(n839), .Y(n464) );
  OAI22X1 U257 ( .A(n312), .B(n855), .C(n311), .D(n839), .Y(n465) );
  OAI22X1 U258 ( .A(n313), .B(n855), .C(n312), .D(n839), .Y(n466) );
  OAI22X1 U259 ( .A(n314), .B(n855), .C(n313), .D(n839), .Y(n467) );
  OAI22X1 U260 ( .A(n315), .B(n854), .C(n314), .D(n838), .Y(n468) );
  OAI22X1 U261 ( .A(n316), .B(n854), .C(n315), .D(n838), .Y(n469) );
  OAI22X1 U262 ( .A(n317), .B(n854), .C(n316), .D(n838), .Y(n470) );
  OAI22X1 U263 ( .A(n318), .B(n854), .C(n317), .D(n838), .Y(n471) );
  OAI22X1 U264 ( .A(n319), .B(n854), .C(n318), .D(n838), .Y(n472) );
  OAI22X1 U265 ( .A(n320), .B(n854), .C(n319), .D(n838), .Y(n473) );
  OAI22X1 U266 ( .A(n191), .B(n854), .C(n320), .D(n838), .Y(n474) );
  OAI22X1 U267 ( .A(n854), .B(n304), .C(n191), .D(n838), .Y(n543) );
  XNOR2X1 U268 ( .A(n869), .B(n831), .Y(n322) );
  XNOR2X1 U269 ( .A(n869), .B(n221), .Y(n323) );
  XNOR2X1 U270 ( .A(n869), .B(n222), .Y(n324) );
  XNOR2X1 U271 ( .A(n869), .B(n223), .Y(n325) );
  XNOR2X1 U272 ( .A(n869), .B(n224), .Y(n326) );
  XNOR2X1 U273 ( .A(n869), .B(n225), .Y(n327) );
  XNOR2X1 U274 ( .A(n869), .B(n226), .Y(n328) );
  XNOR2X1 U275 ( .A(n869), .B(n227), .Y(n329) );
  XNOR2X1 U276 ( .A(n868), .B(n228), .Y(n330) );
  XNOR2X1 U277 ( .A(n868), .B(n229), .Y(n331) );
  XNOR2X1 U278 ( .A(n868), .B(n230), .Y(n332) );
  XNOR2X1 U279 ( .A(n868), .B(n231), .Y(n333) );
  XNOR2X1 U280 ( .A(n868), .B(n232), .Y(n334) );
  XNOR2X1 U281 ( .A(n868), .B(n233), .Y(n335) );
  XNOR2X1 U282 ( .A(n868), .B(n234), .Y(n336) );
  XNOR2X1 U283 ( .A(n868), .B(n235), .Y(n337) );
  OAI22X1 U284 ( .A(n323), .B(n853), .C(n322), .D(n837), .Y(n477) );
  OAI22X1 U285 ( .A(n324), .B(n853), .C(n323), .D(n837), .Y(n478) );
  OAI22X1 U286 ( .A(n325), .B(n853), .C(n324), .D(n837), .Y(n479) );
  OAI22X1 U287 ( .A(n326), .B(n853), .C(n325), .D(n837), .Y(n480) );
  OAI22X1 U288 ( .A(n327), .B(n853), .C(n326), .D(n837), .Y(n481) );
  OAI22X1 U289 ( .A(n328), .B(n853), .C(n327), .D(n837), .Y(n482) );
  OAI22X1 U290 ( .A(n329), .B(n853), .C(n328), .D(n837), .Y(n483) );
  OAI22X1 U291 ( .A(n330), .B(n853), .C(n329), .D(n837), .Y(n484) );
  OAI22X1 U292 ( .A(n331), .B(n853), .C(n330), .D(n837), .Y(n485) );
  OAI22X1 U293 ( .A(n332), .B(n852), .C(n331), .D(n836), .Y(n486) );
  OAI22X1 U294 ( .A(n333), .B(n852), .C(n332), .D(n836), .Y(n487) );
  OAI22X1 U295 ( .A(n334), .B(n852), .C(n333), .D(n836), .Y(n488) );
  OAI22X1 U296 ( .A(n335), .B(n852), .C(n334), .D(n836), .Y(n489) );
  OAI22X1 U297 ( .A(n336), .B(n852), .C(n335), .D(n836), .Y(n490) );
  OAI22X1 U298 ( .A(n337), .B(n852), .C(n336), .D(n836), .Y(n491) );
  OAI22X1 U299 ( .A(n192), .B(n852), .C(n337), .D(n836), .Y(n492) );
  OAI22X1 U300 ( .A(n852), .B(n321), .C(n192), .D(n836), .Y(n544) );
  XNOR2X1 U301 ( .A(n867), .B(n831), .Y(n339) );
  XNOR2X1 U302 ( .A(n867), .B(n221), .Y(n340) );
  XNOR2X1 U303 ( .A(n867), .B(n222), .Y(n341) );
  XNOR2X1 U304 ( .A(n867), .B(n223), .Y(n342) );
  XNOR2X1 U305 ( .A(n867), .B(n224), .Y(n343) );
  XNOR2X1 U306 ( .A(n867), .B(n225), .Y(n344) );
  XNOR2X1 U307 ( .A(n867), .B(n226), .Y(n345) );
  XNOR2X1 U308 ( .A(n867), .B(n227), .Y(n346) );
  XNOR2X1 U309 ( .A(n866), .B(n228), .Y(n347) );
  XNOR2X1 U310 ( .A(n866), .B(n229), .Y(n348) );
  XNOR2X1 U311 ( .A(n866), .B(n230), .Y(n349) );
  XNOR2X1 U312 ( .A(n866), .B(n231), .Y(n350) );
  XNOR2X1 U313 ( .A(n866), .B(n232), .Y(n351) );
  XNOR2X1 U314 ( .A(n866), .B(n233), .Y(n352) );
  XNOR2X1 U315 ( .A(n866), .B(n234), .Y(n353) );
  XNOR2X1 U316 ( .A(n866), .B(n235), .Y(n354) );
  OAI22X1 U317 ( .A(n340), .B(n851), .C(n339), .D(n835), .Y(n495) );
  OAI22X1 U318 ( .A(n341), .B(n851), .C(n340), .D(n835), .Y(n496) );
  OAI22X1 U319 ( .A(n342), .B(n851), .C(n341), .D(n835), .Y(n497) );
  OAI22X1 U320 ( .A(n343), .B(n851), .C(n342), .D(n835), .Y(n498) );
  OAI22X1 U321 ( .A(n344), .B(n851), .C(n343), .D(n835), .Y(n499) );
  OAI22X1 U322 ( .A(n345), .B(n851), .C(n344), .D(n835), .Y(n500) );
  OAI22X1 U323 ( .A(n346), .B(n851), .C(n345), .D(n835), .Y(n501) );
  OAI22X1 U324 ( .A(n347), .B(n851), .C(n346), .D(n835), .Y(n502) );
  OAI22X1 U325 ( .A(n348), .B(n851), .C(n347), .D(n835), .Y(n503) );
  OAI22X1 U326 ( .A(n349), .B(n850), .C(n348), .D(n834), .Y(n504) );
  OAI22X1 U327 ( .A(n350), .B(n850), .C(n349), .D(n834), .Y(n505) );
  OAI22X1 U328 ( .A(n351), .B(n850), .C(n350), .D(n834), .Y(n506) );
  OAI22X1 U329 ( .A(n352), .B(n850), .C(n351), .D(n834), .Y(n507) );
  OAI22X1 U330 ( .A(n353), .B(n850), .C(n352), .D(n834), .Y(n508) );
  OAI22X1 U331 ( .A(n354), .B(n850), .C(n353), .D(n834), .Y(n509) );
  OAI22X1 U332 ( .A(n193), .B(n850), .C(n354), .D(n834), .Y(n510) );
  OAI22X1 U333 ( .A(n850), .B(n338), .C(n193), .D(n834), .Y(n545) );
  XNOR2X1 U334 ( .A(n865), .B(n831), .Y(n356) );
  XNOR2X1 U335 ( .A(n865), .B(n221), .Y(n357) );
  XNOR2X1 U336 ( .A(n865), .B(n222), .Y(n358) );
  XNOR2X1 U337 ( .A(n865), .B(n223), .Y(n359) );
  XNOR2X1 U338 ( .A(n865), .B(n224), .Y(n360) );
  XNOR2X1 U339 ( .A(n865), .B(n225), .Y(n361) );
  XNOR2X1 U340 ( .A(n865), .B(n226), .Y(n362) );
  XNOR2X1 U341 ( .A(n865), .B(n227), .Y(n363) );
  XNOR2X1 U342 ( .A(n864), .B(n228), .Y(n364) );
  XNOR2X1 U343 ( .A(n864), .B(n229), .Y(n365) );
  XNOR2X1 U344 ( .A(n864), .B(n230), .Y(n366) );
  XNOR2X1 U345 ( .A(n864), .B(n231), .Y(n367) );
  XNOR2X1 U346 ( .A(n864), .B(n232), .Y(n368) );
  XNOR2X1 U347 ( .A(n864), .B(n233), .Y(n369) );
  XNOR2X1 U348 ( .A(n864), .B(n234), .Y(n370) );
  XNOR2X1 U349 ( .A(n864), .B(n235), .Y(n371) );
  OAI22X1 U350 ( .A(n357), .B(n849), .C(n356), .D(n833), .Y(n513) );
  OAI22X1 U351 ( .A(n358), .B(n849), .C(n357), .D(n833), .Y(n514) );
  OAI22X1 U352 ( .A(n359), .B(n849), .C(n358), .D(n833), .Y(n515) );
  OAI22X1 U353 ( .A(n360), .B(n849), .C(n359), .D(n833), .Y(n516) );
  OAI22X1 U354 ( .A(n361), .B(n849), .C(n360), .D(n833), .Y(n517) );
  OAI22X1 U355 ( .A(n362), .B(n849), .C(n361), .D(n833), .Y(n518) );
  OAI22X1 U356 ( .A(n363), .B(n849), .C(n362), .D(n833), .Y(n519) );
  OAI22X1 U357 ( .A(n364), .B(n849), .C(n363), .D(n833), .Y(n520) );
  OAI22X1 U358 ( .A(n365), .B(n849), .C(n364), .D(n833), .Y(n521) );
  OAI22X1 U359 ( .A(n366), .B(n848), .C(n365), .D(n832), .Y(n522) );
  OAI22X1 U360 ( .A(n367), .B(n848), .C(n366), .D(n832), .Y(n523) );
  OAI22X1 U361 ( .A(n368), .B(n848), .C(n367), .D(n832), .Y(n524) );
  OAI22X1 U362 ( .A(n369), .B(n848), .C(n368), .D(n832), .Y(n525) );
  OAI22X1 U363 ( .A(n370), .B(n848), .C(n369), .D(n832), .Y(n526) );
  OAI22X1 U364 ( .A(n371), .B(n848), .C(n370), .D(n832), .Y(n527) );
  OAI22X1 U365 ( .A(n178), .B(n848), .C(n371), .D(n832), .Y(n528) );
  OAI22X1 U366 ( .A(n848), .B(n355), .C(n178), .D(n832), .Y(n546) );
  INVX2 U367 ( .A(n221), .Y(n372) );
  INVX2 U368 ( .A(n222), .Y(n373) );
  INVX2 U369 ( .A(n223), .Y(n374) );
  INVX2 U370 ( .A(n224), .Y(n375) );
  INVX2 U371 ( .A(n225), .Y(n376) );
  INVX2 U372 ( .A(n226), .Y(n377) );
  INVX2 U373 ( .A(n227), .Y(n378) );
  INVX2 U374 ( .A(n228), .Y(n379) );
  INVX2 U375 ( .A(n229), .Y(n380) );
  INVX2 U376 ( .A(n230), .Y(n381) );
  INVX2 U377 ( .A(n231), .Y(n382) );
  INVX2 U378 ( .A(n232), .Y(n383) );
  INVX2 U379 ( .A(n233), .Y(n384) );
  INVX2 U380 ( .A(n234), .Y(n385) );
  INVX2 U381 ( .A(n235), .Y(n386) );
  NOR2X1 U382 ( .A(n372), .B(n203), .Y(n675) );
  NOR2X1 U383 ( .A(n373), .B(n203), .Y(n531) );
  NOR2X1 U384 ( .A(n374), .B(n203), .Y(n532) );
  NOR2X1 U385 ( .A(n375), .B(n203), .Y(n705) );
  NOR2X1 U386 ( .A(n376), .B(n203), .Y(n533) );
  NOR2X1 U387 ( .A(n377), .B(n203), .Y(n731) );
  NOR2X1 U388 ( .A(n378), .B(n203), .Y(n534) );
  NOR2X1 U389 ( .A(n379), .B(n203), .Y(n753) );
  NOR2X1 U390 ( .A(n380), .B(n203), .Y(n535) );
  NOR2X1 U391 ( .A(n381), .B(n203), .Y(n771) );
  NOR2X1 U392 ( .A(n382), .B(n203), .Y(n536) );
  NOR2X1 U393 ( .A(n383), .B(n203), .Y(n785) );
  NOR2X1 U394 ( .A(n384), .B(n203), .Y(n537) );
  NOR2X1 U395 ( .A(n385), .B(n203), .Y(n795) );
  NOR2X1 U396 ( .A(n386), .B(n203), .Y(n538) );
  HAX1 U397 ( .A(n389), .B(n405), .YC(n548), .YS(n547) );
  FAX1 U398 ( .A(n390), .B(n406), .C(n548), .YC(n550), .YS(n549) );
  HAX1 U399 ( .A(n391), .B(n541), .YC(n552), .YS(n551) );
  FAX1 U400 ( .A(n407), .B(n423), .C(n551), .YC(n554), .YS(n553) );
  FAX1 U401 ( .A(n392), .B(n424), .C(n408), .YC(n556), .YS(n555) );
  FAX1 U402 ( .A(n552), .B(n943), .C(n555), .YC(n558), .YS(n557) );
  HAX1 U403 ( .A(n393), .B(n542), .YC(n560), .YS(n559) );
  FAX1 U404 ( .A(n409), .B(n441), .C(n425), .YC(n562), .YS(n561) );
  FAX1 U405 ( .A(n559), .B(n556), .C(n561), .YC(n564), .YS(n563) );
  FAX1 U406 ( .A(n394), .B(n426), .C(n442), .YC(n566), .YS(n565) );
  FAX1 U407 ( .A(n410), .B(n560), .C(n946), .YC(n568), .YS(n567) );
  FAX1 U408 ( .A(n562), .B(n565), .C(n567), .YC(n570), .YS(n569) );
  HAX1 U409 ( .A(n395), .B(n543), .YC(n572), .YS(n571) );
  FAX1 U410 ( .A(n443), .B(n459), .C(n427), .YC(n574), .YS(n573) );
  FAX1 U411 ( .A(n411), .B(n571), .C(n566), .YC(n576), .YS(n575) );
  FAX1 U412 ( .A(n573), .B(n568), .C(n575), .YC(n578), .YS(n577) );
  FAX1 U413 ( .A(n396), .B(n412), .C(n428), .YC(n580), .YS(n579) );
  FAX1 U414 ( .A(n444), .B(n460), .C(n572), .YC(n582), .YS(n581) );
  FAX1 U415 ( .A(n941), .B(n574), .C(n579), .YC(n584), .YS(n583) );
  FAX1 U416 ( .A(n581), .B(n576), .C(n583), .YC(n586), .YS(n585) );
  HAX1 U417 ( .A(n397), .B(n544), .YC(n588), .YS(n587) );
  FAX1 U418 ( .A(n445), .B(n477), .C(n413), .YC(n590), .YS(n589) );
  FAX1 U419 ( .A(n429), .B(n461), .C(n587), .YC(n592), .YS(n591) );
  FAX1 U420 ( .A(n580), .B(n589), .C(n582), .YC(n594), .YS(n593) );
  FAX1 U421 ( .A(n591), .B(n584), .C(n593), .YC(n596), .YS(n595) );
  FAX1 U422 ( .A(n398), .B(n414), .C(n478), .YC(n598), .YS(n597) );
  FAX1 U423 ( .A(n430), .B(n462), .C(n446), .YC(n600), .YS(n599) );
  FAX1 U424 ( .A(n588), .B(n942), .C(n590), .YC(n602), .YS(n601) );
  FAX1 U425 ( .A(n597), .B(n599), .C(n592), .YC(n604), .YS(n603) );
  FAX1 U426 ( .A(n601), .B(n594), .C(n603), .YC(n606), .YS(n605) );
  HAX1 U427 ( .A(n399), .B(n545), .YC(n608), .YS(n607) );
  FAX1 U428 ( .A(n463), .B(n415), .C(n431), .YC(n610), .YS(n609) );
  FAX1 U429 ( .A(n447), .B(n495), .C(n479), .YC(n612), .YS(n611) );
  FAX1 U430 ( .A(n607), .B(n598), .C(n600), .YC(n614), .YS(n613) );
  FAX1 U431 ( .A(n611), .B(n609), .C(n602), .YC(n616), .YS(n615) );
  FAX1 U432 ( .A(n613), .B(n604), .C(n615), .YC(n618), .YS(n617) );
  FAX1 U433 ( .A(n400), .B(n416), .C(n432), .YC(n620), .YS(n619) );
  FAX1 U434 ( .A(n448), .B(n496), .C(n480), .YC(n622), .YS(n621) );
  FAX1 U435 ( .A(n464), .B(n608), .C(n945), .YC(n624), .YS(n623) );
  FAX1 U436 ( .A(n610), .B(n612), .C(n619), .YC(n626), .YS(n625) );
  FAX1 U437 ( .A(n621), .B(n623), .C(n614), .YC(n628), .YS(n627) );
  FAX1 U438 ( .A(n625), .B(n616), .C(n627), .YC(n630), .YS(n629) );
  HAX1 U439 ( .A(n401), .B(n546), .YC(n632), .YS(n631) );
  FAX1 U440 ( .A(n465), .B(n513), .C(n497), .YC(n634), .YS(n633) );
  FAX1 U441 ( .A(n417), .B(n481), .C(n449), .YC(n636), .YS(n635) );
  FAX1 U442 ( .A(n433), .B(n631), .C(n620), .YC(n638), .YS(n637) );
  FAX1 U443 ( .A(n622), .B(n635), .C(n633), .YC(n640), .YS(n639) );
  FAX1 U444 ( .A(n624), .B(n626), .C(n637), .YC(n642), .YS(n641) );
  FAX1 U445 ( .A(n639), .B(n628), .C(n641), .YC(n644), .YS(n643) );
  FAX1 U446 ( .A(n402), .B(n418), .C(n947), .YC(n646), .YS(n645) );
  FAX1 U447 ( .A(n434), .B(n514), .C(n498), .YC(n648), .YS(n647) );
  FAX1 U448 ( .A(n450), .B(n482), .C(n466), .YC(n650), .YS(n649) );
  FAX1 U449 ( .A(n632), .B(n634), .C(n636), .YC(n652), .YS(n651) );
  FAX1 U450 ( .A(n645), .B(n649), .C(n647), .YC(n654), .YS(n653) );
  FAX1 U451 ( .A(n638), .B(n640), .C(n651), .YC(n656), .YS(n655) );
  FAX1 U452 ( .A(n653), .B(n642), .C(n655), .YC(n658), .YS(n657) );
  INVX2 U453 ( .A(n675), .Y(n659) );
  FAX1 U454 ( .A(n659), .B(n499), .C(n451), .YC(n661), .YS(n660) );
  FAX1 U455 ( .A(n467), .B(n483), .C(n515), .YC(n663), .YS(n662) );
  FAX1 U456 ( .A(n419), .B(n435), .C(n403), .YC(n665), .YS(n664) );
  FAX1 U457 ( .A(n646), .B(n648), .C(n650), .YC(n667), .YS(n666) );
  FAX1 U458 ( .A(n660), .B(n662), .C(n664), .YC(n669), .YS(n668) );
  FAX1 U459 ( .A(n652), .B(n654), .C(n666), .YC(n671), .YS(n670) );
  FAX1 U460 ( .A(n668), .B(n656), .C(n670), .YC(n673), .YS(n672) );
  FAX1 U462 ( .A(n531), .B(n659), .C(n420), .YC(n677), .YS(n676) );
  FAX1 U463 ( .A(n436), .B(n516), .C(n452), .YC(n679), .YS(n678) );
  FAX1 U464 ( .A(n468), .B(n500), .C(n484), .YC(n681), .YS(n680) );
  FAX1 U465 ( .A(n661), .B(n663), .C(n676), .YC(n683), .YS(n682) );
  FAX1 U466 ( .A(n680), .B(n678), .C(n665), .YC(n685), .YS(n684) );
  FAX1 U467 ( .A(n667), .B(n682), .C(n669), .YC(n687), .YS(n686) );
  FAX1 U468 ( .A(n684), .B(n671), .C(n686), .YC(n689), .YS(n688) );
  FAX1 U469 ( .A(n675), .B(n532), .C(n469), .YC(n691), .YS(n690) );
  FAX1 U470 ( .A(n485), .B(n501), .C(n517), .YC(n693), .YS(n692) );
  FAX1 U471 ( .A(n437), .B(n453), .C(n421), .YC(n695), .YS(n694) );
  FAX1 U472 ( .A(n677), .B(n679), .C(n681), .YC(n697), .YS(n696) );
  FAX1 U473 ( .A(n690), .B(n692), .C(n694), .YC(n699), .YS(n698) );
  FAX1 U474 ( .A(n683), .B(n696), .C(n685), .YC(n701), .YS(n700) );
  FAX1 U475 ( .A(n698), .B(n687), .C(n700), .YC(n703), .YS(n702) );
  INVX2 U476 ( .A(n705), .Y(n704) );
  FAX1 U477 ( .A(n704), .B(n438), .C(n454), .YC(n707), .YS(n706) );
  FAX1 U478 ( .A(n518), .B(n470), .C(n486), .YC(n709), .YS(n708) );
  FAX1 U479 ( .A(n502), .B(n691), .C(n693), .YC(n711), .YS(n710) );
  FAX1 U480 ( .A(n706), .B(n708), .C(n695), .YC(n713), .YS(n712) );
  FAX1 U481 ( .A(n697), .B(n710), .C(n699), .YC(n715), .YS(n714) );
  FAX1 U482 ( .A(n712), .B(n701), .C(n714), .YC(n717), .YS(n716) );
  FAX1 U483 ( .A(n705), .B(n533), .C(n471), .YC(n719), .YS(n718) );
  FAX1 U484 ( .A(n487), .B(n519), .C(n455), .YC(n721), .YS(n720) );
  FAX1 U485 ( .A(n503), .B(n439), .C(n707), .YC(n723), .YS(n722) );
  FAX1 U486 ( .A(n709), .B(n718), .C(n720), .YC(n725), .YS(n724) );
  FAX1 U487 ( .A(n711), .B(n722), .C(n713), .YC(n727), .YS(n726) );
  FAX1 U488 ( .A(n724), .B(n715), .C(n726), .YC(n729), .YS(n728) );
  INVX2 U489 ( .A(n731), .Y(n730) );
  FAX1 U490 ( .A(n730), .B(n456), .C(n472), .YC(n733), .YS(n732) );
  FAX1 U491 ( .A(n520), .B(n504), .C(n488), .YC(n735), .YS(n734) );
  FAX1 U492 ( .A(n719), .B(n721), .C(n732), .YC(n737), .YS(n736) );
  FAX1 U493 ( .A(n734), .B(n723), .C(n725), .YC(n739), .YS(n738) );
  FAX1 U494 ( .A(n736), .B(n727), .C(n738), .YC(n741), .YS(n740) );
  FAX1 U495 ( .A(n731), .B(n534), .C(n489), .YC(n743), .YS(n742) );
  FAX1 U496 ( .A(n505), .B(n521), .C(n473), .YC(n745), .YS(n744) );
  FAX1 U497 ( .A(n457), .B(n733), .C(n735), .YC(n747), .YS(n746) );
  FAX1 U498 ( .A(n742), .B(n744), .C(n737), .YC(n749), .YS(n748) );
  FAX1 U499 ( .A(n746), .B(n739), .C(n748), .YC(n751), .YS(n750) );
  INVX2 U500 ( .A(n753), .Y(n752) );
  FAX1 U501 ( .A(n752), .B(n474), .C(n490), .YC(n755), .YS(n754) );
  FAX1 U502 ( .A(n506), .B(n522), .C(n743), .YC(n757), .YS(n756) );
  FAX1 U503 ( .A(n745), .B(n754), .C(n756), .YC(n759), .YS(n758) );
  FAX1 U504 ( .A(n747), .B(n749), .C(n758), .YC(n761), .YS(n760) );
  FAX1 U505 ( .A(n753), .B(n535), .C(n491), .YC(n763), .YS(n762) );
  FAX1 U506 ( .A(n523), .B(n507), .C(n475), .YC(n765), .YS(n764) );
  FAX1 U507 ( .A(n755), .B(n762), .C(n764), .YC(n767), .YS(n766) );
  FAX1 U508 ( .A(n757), .B(n766), .C(n759), .YC(n769), .YS(n768) );
  INVX2 U509 ( .A(n771), .Y(n770) );
  FAX1 U510 ( .A(n770), .B(n492), .C(n508), .YC(n773), .YS(n772) );
  FAX1 U511 ( .A(n524), .B(n763), .C(n772), .YC(n775), .YS(n774) );
  FAX1 U512 ( .A(n765), .B(n774), .C(n767), .YC(n777), .YS(n776) );
  FAX1 U513 ( .A(n771), .B(n536), .C(n509), .YC(n779), .YS(n778) );
  FAX1 U514 ( .A(n525), .B(n493), .C(n773), .YC(n781), .YS(n780) );
  FAX1 U515 ( .A(n778), .B(n775), .C(n780), .YC(n783), .YS(n782) );
  INVX2 U516 ( .A(n785), .Y(n784) );
  FAX1 U517 ( .A(n784), .B(n510), .C(n526), .YC(n787), .YS(n786) );
  FAX1 U518 ( .A(n779), .B(n786), .C(n781), .YC(n789), .YS(n788) );
  FAX1 U519 ( .A(n785), .B(n537), .C(n527), .YC(n791), .YS(n790) );
  FAX1 U520 ( .A(n511), .B(n787), .C(n790), .YC(n793), .YS(n792) );
  INVX2 U521 ( .A(n795), .Y(n794) );
  FAX1 U522 ( .A(n794), .B(n528), .C(n791), .YC(n797), .YS(n796) );
  HAX1 U523 ( .A(n539), .B(n387), .YC(n799), .YS(product[1]) );
  FAX1 U524 ( .A(n388), .B(n799), .C(n944), .YC(n800), .YS(product[2]) );
  FAX1 U525 ( .A(n540), .B(n547), .C(n800), .YC(n801), .YS(product[3]) );
  FAX1 U526 ( .A(n940), .B(n549), .C(n801), .YC(n802), .YS(product[4]) );
  FAX1 U527 ( .A(n550), .B(n553), .C(n802), .YC(n803), .YS(product[5]) );
  FAX1 U528 ( .A(n554), .B(n557), .C(n803), .YC(n804), .YS(product[6]) );
  FAX1 U529 ( .A(n558), .B(n563), .C(n804), .YC(n805), .YS(product[7]) );
  FAX1 U530 ( .A(n564), .B(n569), .C(n805), .YC(n806), .YS(product[8]) );
  FAX1 U531 ( .A(n570), .B(n577), .C(n806), .YC(n807), .YS(product[9]) );
  FAX1 U532 ( .A(n578), .B(n585), .C(n807), .YC(n808), .YS(product[10]) );
  FAX1 U533 ( .A(n586), .B(n595), .C(n808), .YC(n809), .YS(product[11]) );
  FAX1 U534 ( .A(n596), .B(n605), .C(n809), .YC(n810), .YS(product[12]) );
  FAX1 U535 ( .A(n606), .B(n617), .C(n810), .YC(n811), .YS(product[13]) );
  FAX1 U536 ( .A(n618), .B(n629), .C(n811), .YC(n812), .YS(product[14]) );
  FAX1 U537 ( .A(n630), .B(n643), .C(n812), .YC(n813), .YS(product[15]) );
  FAX1 U538 ( .A(n644), .B(n657), .C(n813), .YC(n814), .YS(product[16]) );
  FAX1 U539 ( .A(n658), .B(n672), .C(n814), .YC(n815), .YS(product[17]) );
  FAX1 U540 ( .A(n673), .B(n688), .C(n815), .YC(n816), .YS(product[18]) );
  FAX1 U541 ( .A(n689), .B(n702), .C(n816), .YC(n817), .YS(product[19]) );
  FAX1 U542 ( .A(n703), .B(n716), .C(n817), .YC(n818), .YS(product[20]) );
  FAX1 U543 ( .A(n717), .B(n728), .C(n818), .YC(n819), .YS(product[21]) );
  FAX1 U544 ( .A(n729), .B(n740), .C(n819), .YC(n820), .YS(product[22]) );
  FAX1 U545 ( .A(n741), .B(n750), .C(n820), .YC(n821), .YS(product[23]) );
  FAX1 U546 ( .A(n751), .B(n760), .C(n821), .YC(n822), .YS(product[24]) );
  FAX1 U547 ( .A(n761), .B(n768), .C(n822), .YC(n823), .YS(product[25]) );
  FAX1 U548 ( .A(n776), .B(n769), .C(n823), .YC(n824), .YS(product[26]) );
  FAX1 U549 ( .A(n782), .B(n777), .C(n824), .YC(n825), .YS(product[27]) );
  FAX1 U550 ( .A(n788), .B(n783), .C(n825), .YC(n826), .YS(product[28]) );
  FAX1 U551 ( .A(n792), .B(n789), .C(n826), .YC(n827), .YS(product[29]) );
  FAX1 U552 ( .A(n796), .B(n793), .C(n827), .YC(n828), .YS(product[30]) );
  XOR2X1 U553 ( .A(n797), .B(n798), .Y(n829) );
  XOR2X1 U554 ( .A(n828), .B(n829), .Y(product[31]) );
  AND2X2 U607 ( .A(n831), .B(a[0]), .Y(product[0]) );
  AND2X2 U608 ( .A(n830), .B(n134), .Y(n940) );
  AND2X2 U609 ( .A(n830), .B(n86), .Y(n941) );
  AND2X2 U610 ( .A(n830), .B(n60), .Y(n942) );
  AND2X2 U611 ( .A(n830), .B(n118), .Y(n943) );
  AND2X2 U612 ( .A(n831), .B(n150), .Y(n944) );
  AND2X2 U613 ( .A(n830), .B(n26), .Y(n945) );
  AND2X2 U614 ( .A(n830), .B(n102), .Y(n946) );
  AND2X2 U615 ( .A(n830), .B(a[15]), .Y(n947) );
  BUFX2 U616 ( .A(n205), .Y(n845) );
  BUFX2 U617 ( .A(n206), .Y(n843) );
  BUFX2 U618 ( .A(n207), .Y(n841) );
  BUFX2 U619 ( .A(n208), .Y(n839) );
  BUFX2 U620 ( .A(n209), .Y(n837) );
  BUFX2 U621 ( .A(n210), .Y(n835) );
  BUFX2 U622 ( .A(n211), .Y(n833) );
  BUFX2 U623 ( .A(n204), .Y(n847) );
  BUFX2 U624 ( .A(n196), .Y(n861) );
  BUFX2 U625 ( .A(n197), .Y(n859) );
  BUFX2 U626 ( .A(n198), .Y(n857) );
  BUFX2 U627 ( .A(n199), .Y(n855) );
  BUFX2 U628 ( .A(n200), .Y(n853) );
  BUFX2 U629 ( .A(n201), .Y(n851) );
  BUFX2 U630 ( .A(n202), .Y(n849) );
  BUFX2 U631 ( .A(n196), .Y(n860) );
  BUFX2 U632 ( .A(n197), .Y(n858) );
  BUFX2 U633 ( .A(n198), .Y(n856) );
  BUFX2 U634 ( .A(n199), .Y(n854) );
  BUFX2 U635 ( .A(n200), .Y(n852) );
  BUFX2 U636 ( .A(n201), .Y(n850) );
  BUFX2 U637 ( .A(n202), .Y(n848) );
  BUFX2 U638 ( .A(n195), .Y(n862) );
  BUFX2 U639 ( .A(n205), .Y(n844) );
  BUFX2 U640 ( .A(n206), .Y(n842) );
  BUFX2 U641 ( .A(n207), .Y(n840) );
  BUFX2 U642 ( .A(n208), .Y(n838) );
  BUFX2 U643 ( .A(n209), .Y(n836) );
  BUFX2 U644 ( .A(n211), .Y(n832) );
  BUFX2 U645 ( .A(n210), .Y(n834) );
  BUFX2 U646 ( .A(n204), .Y(n846) );
  BUFX2 U647 ( .A(n195), .Y(n863) );
  BUFX2 U648 ( .A(b[0]), .Y(n831) );
  BUFX2 U649 ( .A(a[1]), .Y(n879) );
  BUFX2 U650 ( .A(a[5]), .Y(n875) );
  BUFX2 U651 ( .A(a[3]), .Y(n877) );
  BUFX2 U652 ( .A(a[7]), .Y(n873) );
  BUFX2 U653 ( .A(a[9]), .Y(n871) );
  BUFX2 U654 ( .A(a[11]), .Y(n869) );
  BUFX2 U655 ( .A(a[13]), .Y(n867) );
  BUFX2 U656 ( .A(a[15]), .Y(n865) );
  BUFX2 U657 ( .A(a[1]), .Y(n878) );
  BUFX2 U658 ( .A(a[3]), .Y(n876) );
  BUFX2 U659 ( .A(a[5]), .Y(n874) );
  BUFX2 U660 ( .A(a[7]), .Y(n872) );
  BUFX2 U661 ( .A(a[9]), .Y(n870) );
  BUFX2 U662 ( .A(a[11]), .Y(n868) );
  BUFX2 U663 ( .A(a[13]), .Y(n866) );
  BUFX2 U664 ( .A(a[15]), .Y(n864) );
  BUFX2 U665 ( .A(n178), .Y(n203) );
  BUFX2 U666 ( .A(b[0]), .Y(n830) );
  BUFX2 U667 ( .A(b[1]), .Y(n221) );
  BUFX2 U668 ( .A(b[2]), .Y(n222) );
  BUFX2 U669 ( .A(b[3]), .Y(n223) );
  BUFX2 U670 ( .A(b[4]), .Y(n224) );
  BUFX2 U671 ( .A(b[5]), .Y(n225) );
  BUFX2 U672 ( .A(b[6]), .Y(n226) );
  BUFX2 U673 ( .A(b[7]), .Y(n227) );
  BUFX2 U674 ( .A(b[8]), .Y(n228) );
  BUFX2 U675 ( .A(b[9]), .Y(n229) );
  BUFX2 U676 ( .A(b[10]), .Y(n230) );
  BUFX2 U677 ( .A(b[11]), .Y(n231) );
  BUFX2 U678 ( .A(b[12]), .Y(n232) );
  BUFX2 U679 ( .A(b[13]), .Y(n233) );
  BUFX2 U680 ( .A(b[14]), .Y(n234) );
  BUFX2 U681 ( .A(b[15]), .Y(n235) );
endmodule


module alu ( reg_A, reg_B, ctrl_ww, alu_op, result );
  input [0:127] reg_A;
  input [0:127] reg_B;
  input [0:1] ctrl_ww;
  input [0:4] alu_op;
  output [0:127] result;
  wire   n228_1_, n228_2_, n228_3_, n228_6_, slice455_4_, slice455_5_,
         slice455_7_, slice455_8_, slice455_9_, slice455_10_, slice455_11_,
         slice455_12_, slice455_13_, slice455_14_, slice455_15_, slice455_16_,
         n203_1_, n203_4_, slice356_2_, slice356_3_, slice356_5_, slice356_6_,
         slice356_7_, slice356_8_, slice356_9_, slice356_10_, slice356_11_,
         slice356_12_, slice356_13_, slice356_14_, slice356_15_, slice356_16_,
         n208_1_, n208_2_, n208_3_, n208_6_, slice376_4_, slice376_5_,
         slice376_7_, slice376_8_, slice376_9_, slice376_10_, slice376_11_,
         slice376_12_, slice376_13_, slice376_14_, slice376_15_, slice376_16_,
         slice376_17_, slice376_18_, slice376_19_, slice376_20_, slice376_21_,
         slice376_22_, slice376_23_, slice376_24_, slice376_25_, slice376_26_,
         slice376_27_, slice376_28_, slice376_29_, slice376_30_, slice376_31_,
         slice376_32_, n213_1_, n213_2_, n213_3_, n213_6_, slice396_4_,
         slice396_5_, slice396_7_, slice396_8_, slice396_9_, slice396_10_,
         slice396_11_, slice396_12_, slice396_13_, slice396_14_, slice396_15_,
         slice396_16_, slice396_17_, slice396_18_, slice396_19_, slice396_20_,
         slice396_21_, slice396_22_, slice396_23_, slice396_24_, slice396_25_,
         slice396_26_, slice396_27_, slice396_28_, slice396_29_, slice396_30_,
         slice396_31_, slice396_32_, n218_1_, n218_2_, n218_3_, n218_6_,
         slice416_4_, slice416_5_, slice416_7_, slice416_8_, slice416_9_,
         slice416_10_, slice416_11_, slice416_12_, slice416_13_, slice416_14_,
         slice416_15_, slice416_16_, slice673_1_, slice673_2_, slice673_3_,
         slice673_4_, slice673_5_, slice673_6_, slice673_7_, slice673_8_,
         slice673_9_, slice673_10_, slice673_11_, slice673_12_, slice673_13_,
         slice673_14_, slice673_15_, slice673_16_, n313_1_, n313_2_, n313_3_,
         n313_6_, slice693_4_, slice693_5_, slice693_7_, slice693_8_,
         slice693_9_, slice693_10_, slice693_11_, slice693_12_, slice693_13_,
         slice693_14_, slice693_15_, slice693_16_, n328_1_, n328_2_, n328_3_,
         n328_6_, slice753_4_, slice753_5_, slice753_7_, slice753_8_,
         slice753_9_, slice753_10_, slice753_11_, slice753_12_, slice753_13_,
         slice753_14_, slice753_15_, slice753_16_, n333_1_, n333_2_, n333_3_,
         n333_6_, slice773_4_, slice773_5_, slice773_7_, slice773_8_,
         slice773_9_, slice773_10_, slice773_11_, slice773_12_, slice773_13_,
         slice773_14_, slice773_15_, slice773_16_, n338_1_, n338_2_, n338_3_,
         n338_6_, slice793_4_, slice793_5_, slice793_7_, slice793_8_,
         slice793_9_, slice793_10_, slice793_11_, slice793_12_, slice793_13_,
         slice793_14_, slice793_15_, slice793_16_, U69_U1_Z_0, U69_U1_Z_1,
         U69_U1_Z_2, U69_U1_Z_3, U69_U1_Z_4, U69_U1_Z_5, U69_U1_Z_6,
         U69_U1_Z_7, U69_U1_Z_8, U69_U1_Z_9, U69_U1_Z_10, U69_U1_Z_11,
         U69_U1_Z_12, U69_U1_Z_13, U69_U1_Z_14, U69_U1_Z_15, U69_U2_Z_0,
         U69_U2_Z_1, U69_U2_Z_2, U69_U2_Z_3, U69_U2_Z_4, U69_U2_Z_5,
         U69_U2_Z_6, U69_U2_Z_7, U69_U2_Z_8, U69_U2_Z_9, U69_U2_Z_10,
         U69_U2_Z_11, U69_U2_Z_12, U69_U2_Z_13, U69_U2_Z_14, U69_U2_Z_15,
         U69_U3_Z_0, U69_U3_Z_1, U69_U3_Z_2, U69_U3_Z_3, U69_U3_Z_4,
         U69_U3_Z_5, U69_U3_Z_6, U69_U3_Z_7, U69_U3_Z_8, U69_U3_Z_9,
         U69_U3_Z_10, U69_U3_Z_11, U69_U3_Z_12, U69_U3_Z_13, U69_U3_Z_14,
         U69_U3_Z_15, U69_U4_Z_0, U69_U4_Z_1, U69_U4_Z_2, U69_U4_Z_3,
         U69_U4_Z_4, U69_U4_Z_5, U69_U4_Z_6, U69_U4_Z_7, U69_U4_Z_8,
         U69_U4_Z_9, U69_U4_Z_10, U69_U4_Z_11, U69_U4_Z_12, U69_U4_Z_13,
         U69_U4_Z_14, U69_U4_Z_15, U69_U5_Z_0, U69_U5_Z_1, U69_U5_Z_2,
         U69_U5_Z_3, U69_U5_Z_4, U69_U5_Z_5, U69_U5_Z_6, U69_U5_Z_7,
         U69_U6_Z_0, U69_U6_Z_1, U69_U6_Z_2, U69_U6_Z_3, U69_U6_Z_4,
         U69_U6_Z_5, U69_U6_Z_6, U69_U6_Z_7, U69_U7_Z_0, U69_U7_Z_1,
         U69_U7_Z_2, U69_U7_Z_3, U69_U7_Z_4, U69_U7_Z_5, U69_U7_Z_6,
         U69_U7_Z_7, U69_U7_Z_8, U69_U7_Z_9, U69_U7_Z_10, U69_U7_Z_11,
         U69_U7_Z_12, U69_U7_Z_13, U69_U7_Z_14, U69_U7_Z_15, U69_U8_Z_0,
         U69_U8_Z_1, U69_U8_Z_2, U69_U8_Z_3, U69_U8_Z_4, U69_U8_Z_5,
         U69_U8_Z_6, U69_U8_Z_7, U69_U8_Z_8, U69_U8_Z_9, U69_U8_Z_10,
         U69_U8_Z_11, U69_U8_Z_12, U69_U8_Z_13, U69_U8_Z_14, U69_U8_Z_15,
         U69_U9_Z_0, U69_U9_Z_1, U69_U9_Z_2, U69_U9_Z_3, U69_U9_Z_4,
         U69_U9_Z_5, U69_U9_Z_6, U69_U9_Z_7, U69_U9_Z_8, U69_U9_Z_9,
         U69_U9_Z_10, U69_U9_Z_11, U69_U9_Z_12, U69_U9_Z_13, U69_U9_Z_14,
         U69_U9_Z_15, U69_U10_Z_0, U69_U10_Z_1, U69_U10_Z_2, U69_U10_Z_3,
         U69_U10_Z_4, U69_U10_Z_5, U69_U10_Z_6, U69_U10_Z_7, U69_U10_Z_8,
         U69_U10_Z_9, U69_U10_Z_10, U69_U10_Z_11, U69_U10_Z_12, U69_U10_Z_13,
         U69_U10_Z_14, U69_U10_Z_15, U69_U11_Z_0, U69_U11_Z_1, U69_U11_Z_2,
         U69_U11_Z_3, U69_U11_Z_4, U69_U11_Z_5, U69_U11_Z_6, U69_U11_Z_7,
         U69_U12_Z_0, U69_U12_Z_1, U69_U12_Z_2, U69_U12_Z_3, U69_U12_Z_4,
         U69_U12_Z_5, U69_U12_Z_6, U69_U12_Z_7, U69_U13_Z_0, U69_U13_Z_1,
         U69_U13_Z_2, U69_U13_Z_3, U69_U13_Z_4, U69_U13_Z_5, U69_U13_Z_6,
         U69_U13_Z_7, U69_U14_Z_0, U69_U14_Z_1, U69_U14_Z_2, U69_U14_Z_3,
         U69_U14_Z_4, U69_U14_Z_5, U69_U14_Z_6, U69_U14_Z_7, U69_U15_Z_0,
         U69_U15_Z_1, U69_U15_Z_2, U69_U15_Z_3, U69_U15_Z_4, U69_U15_Z_5,
         U69_U15_Z_6, U69_U15_Z_7, U69_U16_Z_0, U69_U16_Z_1, U69_U16_Z_2,
         U69_U16_Z_3, U69_U16_Z_4, U69_U16_Z_5, U69_U16_Z_6, U69_U16_Z_7,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279;

  alu_DW_mult_uns_8 r119 ( .a({U69_U1_Z_15, U69_U1_Z_14, U69_U1_Z_13, 
        U69_U1_Z_12, U69_U1_Z_11, U69_U1_Z_10, U69_U1_Z_9, U69_U1_Z_8, 
        U69_U1_Z_7, U69_U1_Z_6, U69_U1_Z_5, U69_U1_Z_4, U69_U1_Z_3, U69_U1_Z_2, 
        U69_U1_Z_1, U69_U1_Z_0}), .b({U69_U2_Z_15, U69_U2_Z_14, U69_U2_Z_13, 
        U69_U2_Z_12, U69_U2_Z_11, U69_U2_Z_10, U69_U2_Z_9, U69_U2_Z_8, 
        U69_U2_Z_7, U69_U2_Z_6, U69_U2_Z_5, U69_U2_Z_4, U69_U2_Z_3, U69_U2_Z_2, 
        U69_U2_Z_1, U69_U2_Z_0}), .product({n213_1_, n213_2_, n213_3_, 
        slice396_4_, slice396_5_, n213_6_, slice396_7_, slice396_8_, 
        slice396_9_, slice396_10_, slice396_11_, slice396_12_, slice396_13_, 
        slice396_14_, slice396_15_, slice396_16_, slice396_17_, slice396_18_, 
        slice396_19_, slice396_20_, slice396_21_, slice396_22_, slice396_23_, 
        slice396_24_, slice396_25_, slice396_26_, slice396_27_, slice396_28_, 
        slice396_29_, slice396_30_, slice396_31_, slice396_32_}) );
  alu_DW_mult_uns_7 r435 ( .a({U69_U3_Z_15, U69_U3_Z_14, U69_U3_Z_13, 
        U69_U3_Z_12, U69_U3_Z_11, U69_U3_Z_10, U69_U3_Z_9, U69_U3_Z_8, 
        U69_U3_Z_7, U69_U3_Z_6, U69_U3_Z_5, U69_U3_Z_4, U69_U3_Z_3, U69_U3_Z_2, 
        U69_U3_Z_1, U69_U3_Z_0}), .b({U69_U4_Z_15, U69_U4_Z_14, U69_U4_Z_13, 
        U69_U4_Z_12, U69_U4_Z_11, U69_U4_Z_10, U69_U4_Z_9, U69_U4_Z_8, 
        U69_U4_Z_7, U69_U4_Z_6, U69_U4_Z_5, U69_U4_Z_4, U69_U4_Z_3, U69_U4_Z_2, 
        U69_U4_Z_1, U69_U4_Z_0}), .product({n208_1_, n208_2_, n208_3_, 
        slice376_4_, slice376_5_, n208_6_, slice376_7_, slice376_8_, 
        slice376_9_, slice376_10_, slice376_11_, slice376_12_, slice376_13_, 
        slice376_14_, slice376_15_, slice376_16_, slice376_17_, slice376_18_, 
        slice376_19_, slice376_20_, slice376_21_, slice376_22_, slice376_23_, 
        slice376_24_, slice376_25_, slice376_26_, slice376_27_, slice376_28_, 
        slice376_29_, slice376_30_, slice376_31_, slice376_32_}) );
  alu_DW_mult_uns_6 r436 ( .a({U69_U5_Z_7, U69_U5_Z_6, U69_U5_Z_5, U69_U5_Z_4, 
        U69_U5_Z_3, U69_U5_Z_2, U69_U5_Z_1, U69_U5_Z_0}), .b({U69_U6_Z_7, 
        U69_U6_Z_6, U69_U6_Z_5, U69_U6_Z_4, U69_U6_Z_3, U69_U6_Z_2, U69_U6_Z_1, 
        U69_U6_Z_0}), .product({n328_1_, n328_2_, n328_3_, slice753_4_, 
        slice753_5_, n328_6_, slice753_7_, slice753_8_, slice753_9_, 
        slice753_10_, slice753_11_, slice753_12_, slice753_13_, slice753_14_, 
        slice753_15_, slice753_16_}) );
  alu_DW_mult_uns_5 r437 ( .a({U69_U7_Z_15, U69_U7_Z_14, U69_U7_Z_13, 
        U69_U7_Z_12, U69_U7_Z_11, U69_U7_Z_10, U69_U7_Z_9, U69_U7_Z_8, 
        U69_U7_Z_7, U69_U7_Z_6, U69_U7_Z_5, U69_U7_Z_4, U69_U7_Z_3, U69_U7_Z_2, 
        U69_U7_Z_1, U69_U7_Z_0}), .b({U69_U8_Z_15, U69_U8_Z_14, U69_U8_Z_13, 
        U69_U8_Z_12, U69_U8_Z_11, U69_U8_Z_10, U69_U8_Z_9, U69_U8_Z_8, 
        U69_U8_Z_7, U69_U8_Z_6, U69_U8_Z_5, U69_U8_Z_4, U69_U8_Z_3, U69_U8_Z_2, 
        U69_U8_Z_1, U69_U8_Z_0}), .product({n218_1_, n218_2_, n218_3_, 
        slice416_4_, slice416_5_, n218_6_, slice416_7_, slice416_8_, 
        slice416_9_, slice416_10_, slice416_11_, slice416_12_, slice416_13_, 
        slice416_14_, slice416_15_, slice416_16_, n313_1_, n313_2_, n313_3_, 
        slice693_4_, slice693_5_, n313_6_, slice693_7_, slice693_8_, 
        slice693_9_, slice693_10_, slice693_11_, slice693_12_, slice693_13_, 
        slice693_14_, slice693_15_, slice693_16_}) );
  alu_DW_mult_uns_4 r438 ( .a({U69_U9_Z_15, U69_U9_Z_14, U69_U9_Z_13, 
        U69_U9_Z_12, U69_U9_Z_11, U69_U9_Z_10, U69_U9_Z_9, U69_U9_Z_8, 
        U69_U9_Z_7, U69_U9_Z_6, U69_U9_Z_5, U69_U9_Z_4, U69_U9_Z_3, U69_U9_Z_2, 
        U69_U9_Z_1, U69_U9_Z_0}), .b({U69_U10_Z_15, U69_U10_Z_14, U69_U10_Z_13, 
        U69_U10_Z_12, U69_U10_Z_11, U69_U10_Z_10, U69_U10_Z_9, U69_U10_Z_8, 
        U69_U10_Z_7, U69_U10_Z_6, U69_U10_Z_5, U69_U10_Z_4, U69_U10_Z_3, 
        U69_U10_Z_2, U69_U10_Z_1, U69_U10_Z_0}), .product({n203_1_, 
        slice356_2_, slice356_3_, n203_4_, slice356_5_, slice356_6_, 
        slice356_7_, slice356_8_, slice356_9_, slice356_10_, slice356_11_, 
        slice356_12_, slice356_13_, slice356_14_, slice356_15_, slice356_16_, 
        n228_1_, n228_2_, n228_3_, slice455_4_, slice455_5_, n228_6_, 
        slice455_7_, slice455_8_, slice455_9_, slice455_10_, slice455_11_, 
        slice455_12_, slice455_13_, slice455_14_, slice455_15_, slice455_16_})
         );
  alu_DW_mult_uns_3 r439 ( .a({U69_U11_Z_7, U69_U11_Z_6, U69_U11_Z_5, 
        U69_U11_Z_4, U69_U11_Z_3, U69_U11_Z_2, U69_U11_Z_1, U69_U11_Z_0}), .b(
        {U69_U12_Z_7, U69_U12_Z_6, U69_U12_Z_5, U69_U12_Z_4, U69_U12_Z_3, 
        U69_U12_Z_2, U69_U12_Z_1, U69_U12_Z_0}), .product({n333_1_, n333_2_, 
        n333_3_, slice773_4_, slice773_5_, n333_6_, slice773_7_, slice773_8_, 
        slice773_9_, slice773_10_, slice773_11_, slice773_12_, slice773_13_, 
        slice773_14_, slice773_15_, slice773_16_}) );
  alu_DW_mult_uns_2 r440 ( .a({U69_U13_Z_7, U69_U13_Z_6, U69_U13_Z_5, 
        U69_U13_Z_4, U69_U13_Z_3, U69_U13_Z_2, U69_U13_Z_1, U69_U13_Z_0}), .b(
        {U69_U14_Z_7, U69_U14_Z_6, U69_U14_Z_5, U69_U14_Z_4, U69_U14_Z_3, 
        U69_U14_Z_2, U69_U14_Z_1, U69_U14_Z_0}), .product({slice673_1_, 
        slice673_2_, slice673_3_, slice673_4_, slice673_5_, slice673_6_, 
        slice673_7_, slice673_8_, slice673_9_, slice673_10_, slice673_11_, 
        slice673_12_, slice673_13_, slice673_14_, slice673_15_, slice673_16_})
         );
  alu_DW_mult_uns_1 r441 ( .a({U69_U15_Z_7, U69_U15_Z_6, U69_U15_Z_5, 
        U69_U15_Z_4, U69_U15_Z_3, U69_U15_Z_2, U69_U15_Z_1, U69_U15_Z_0}), .b(
        {U69_U16_Z_7, U69_U16_Z_6, U69_U16_Z_5, U69_U16_Z_4, U69_U16_Z_3, 
        U69_U16_Z_2, U69_U16_Z_1, U69_U16_Z_0}), .product({n338_1_, n338_2_, 
        n338_3_, slice793_4_, slice793_5_, n338_6_, slice793_7_, slice793_8_, 
        slice793_9_, slice793_10_, slice793_11_, slice793_12_, slice793_13_, 
        slice793_14_, slice793_15_, slice793_16_}) );
  BUFX2 U918 ( .A(n1777), .Y(n1764) );
  INVX1 U919 ( .A(n1775), .Y(n1765) );
  BUFX2 U920 ( .A(n2048), .Y(n1766) );
  INVX4 U921 ( .A(n1852), .Y(n1775) );
  INVX4 U922 ( .A(n1891), .Y(n1773) );
  INVX4 U923 ( .A(n1890), .Y(n1774) );
  INVX4 U924 ( .A(n2007), .Y(n1772) );
  INVX4 U925 ( .A(n2160), .Y(n1767) );
  INVX4 U926 ( .A(alu_op[2]), .Y(n2011) );
  INVX4 U927 ( .A(n2158), .Y(n1768) );
  INVX2 U928 ( .A(n2020), .Y(n1769) );
  NAND2X1 U929 ( .A(n1770), .B(n1771), .Y(result[9]) );
  AOI22X1 U930 ( .A(slice376_10_), .B(n1772), .C(slice356_10_), .D(n1773), .Y(
        n1771) );
  AOI22X1 U931 ( .A(slice673_10_), .B(n1774), .C(slice396_26_), .D(n1775), .Y(
        n1770) );
  INVX1 U932 ( .A(n1776), .Y(result[99]) );
  AOI22X1 U933 ( .A(slice416_4_), .B(n1764), .C(slice793_4_), .D(n1778), .Y(
        n1776) );
  INVX1 U934 ( .A(n1779), .Y(result[98]) );
  AOI22X1 U935 ( .A(n218_3_), .B(n1764), .C(n338_3_), .D(n1778), .Y(n1779) );
  INVX1 U936 ( .A(n1780), .Y(result[97]) );
  AOI22X1 U937 ( .A(n218_2_), .B(n1764), .C(n338_2_), .D(n1778), .Y(n1780) );
  INVX1 U938 ( .A(n1781), .Y(result[96]) );
  AOI22X1 U939 ( .A(n218_1_), .B(n1764), .C(n338_1_), .D(n1778), .Y(n1781) );
  NAND2X1 U940 ( .A(n1782), .B(n1783), .Y(result[95]) );
  AOI22X1 U941 ( .A(slice455_16_), .B(n1772), .C(slice396_32_), .D(n1773), .Y(
        n1783) );
  AOI22X1 U942 ( .A(slice773_16_), .B(n1774), .C(slice673_16_), .D(n1775), .Y(
        n1782) );
  NAND2X1 U943 ( .A(n1784), .B(n1785), .Y(result[94]) );
  AOI22X1 U944 ( .A(slice455_15_), .B(n1772), .C(slice396_31_), .D(n1773), .Y(
        n1785) );
  AOI22X1 U945 ( .A(slice773_15_), .B(n1774), .C(slice673_15_), .D(n1775), .Y(
        n1784) );
  NAND2X1 U946 ( .A(n1786), .B(n1787), .Y(result[93]) );
  AOI22X1 U947 ( .A(slice455_14_), .B(n1772), .C(slice396_30_), .D(n1773), .Y(
        n1787) );
  AOI22X1 U948 ( .A(slice773_14_), .B(n1774), .C(slice673_14_), .D(n1775), .Y(
        n1786) );
  NAND2X1 U949 ( .A(n1788), .B(n1789), .Y(result[92]) );
  AOI22X1 U950 ( .A(slice455_13_), .B(n1772), .C(slice396_29_), .D(n1773), .Y(
        n1789) );
  AOI22X1 U951 ( .A(slice773_13_), .B(n1774), .C(slice673_13_), .D(n1775), .Y(
        n1788) );
  NAND2X1 U952 ( .A(n1790), .B(n1791), .Y(result[91]) );
  AOI22X1 U953 ( .A(slice455_12_), .B(n1772), .C(slice396_28_), .D(n1773), .Y(
        n1791) );
  AOI22X1 U954 ( .A(slice773_12_), .B(n1774), .C(slice673_12_), .D(n1775), .Y(
        n1790) );
  NAND2X1 U955 ( .A(n1792), .B(n1793), .Y(result[90]) );
  AOI22X1 U956 ( .A(slice455_11_), .B(n1772), .C(slice396_27_), .D(n1773), .Y(
        n1793) );
  AOI22X1 U957 ( .A(slice773_11_), .B(n1774), .C(slice673_11_), .D(n1775), .Y(
        n1792) );
  NAND2X1 U958 ( .A(n1794), .B(n1795), .Y(result[8]) );
  AOI22X1 U959 ( .A(slice376_9_), .B(n1772), .C(slice356_9_), .D(n1773), .Y(
        n1795) );
  AOI22X1 U960 ( .A(slice673_9_), .B(n1774), .C(slice396_25_), .D(n1775), .Y(
        n1794) );
  NAND2X1 U961 ( .A(n1796), .B(n1797), .Y(result[89]) );
  AOI22X1 U962 ( .A(slice455_10_), .B(n1772), .C(slice396_26_), .D(n1773), .Y(
        n1797) );
  AOI22X1 U963 ( .A(slice773_10_), .B(n1774), .C(n1775), .D(slice673_10_), .Y(
        n1796) );
  NAND2X1 U964 ( .A(n1798), .B(n1799), .Y(result[88]) );
  AOI22X1 U965 ( .A(slice455_9_), .B(n1772), .C(slice396_25_), .D(n1773), .Y(
        n1799) );
  AOI22X1 U966 ( .A(slice773_9_), .B(n1774), .C(slice673_9_), .D(n1775), .Y(
        n1798) );
  NAND2X1 U967 ( .A(n1800), .B(n1801), .Y(result[87]) );
  AOI22X1 U968 ( .A(slice455_8_), .B(n1772), .C(slice396_24_), .D(n1773), .Y(
        n1801) );
  AOI22X1 U969 ( .A(slice773_8_), .B(n1774), .C(slice673_8_), .D(n1775), .Y(
        n1800) );
  NAND2X1 U970 ( .A(n1802), .B(n1803), .Y(result[86]) );
  AOI22X1 U971 ( .A(slice455_7_), .B(n1772), .C(slice396_23_), .D(n1773), .Y(
        n1803) );
  AOI22X1 U972 ( .A(slice773_7_), .B(n1774), .C(slice673_7_), .D(n1775), .Y(
        n1802) );
  NAND2X1 U973 ( .A(n1804), .B(n1805), .Y(result[85]) );
  AOI22X1 U974 ( .A(n228_6_), .B(n1772), .C(slice396_22_), .D(n1773), .Y(n1805) );
  AOI22X1 U975 ( .A(n333_6_), .B(n1774), .C(slice673_6_), .D(n1775), .Y(n1804)
         );
  NAND2X1 U976 ( .A(n1806), .B(n1807), .Y(result[84]) );
  AOI22X1 U977 ( .A(slice455_5_), .B(n1772), .C(slice396_21_), .D(n1773), .Y(
        n1807) );
  AOI22X1 U978 ( .A(slice773_5_), .B(n1774), .C(slice673_5_), .D(n1775), .Y(
        n1806) );
  NAND2X1 U979 ( .A(n1808), .B(n1809), .Y(result[83]) );
  AOI22X1 U980 ( .A(slice455_4_), .B(n1772), .C(slice396_20_), .D(n1773), .Y(
        n1809) );
  AOI22X1 U981 ( .A(slice773_4_), .B(n1774), .C(slice673_4_), .D(n1775), .Y(
        n1808) );
  NAND2X1 U982 ( .A(n1810), .B(n1811), .Y(result[82]) );
  AOI22X1 U983 ( .A(n228_3_), .B(n1772), .C(slice396_19_), .D(n1773), .Y(n1811) );
  AOI22X1 U984 ( .A(n333_3_), .B(n1774), .C(slice673_3_), .D(n1775), .Y(n1810)
         );
  NAND2X1 U985 ( .A(n1812), .B(n1813), .Y(result[81]) );
  AOI22X1 U986 ( .A(n228_2_), .B(n1772), .C(slice396_18_), .D(n1773), .Y(n1813) );
  AOI22X1 U987 ( .A(n333_2_), .B(n1774), .C(slice673_2_), .D(n1775), .Y(n1812)
         );
  NAND2X1 U988 ( .A(n1814), .B(n1815), .Y(result[80]) );
  AOI22X1 U989 ( .A(n228_1_), .B(n1772), .C(slice396_17_), .D(n1773), .Y(n1815) );
  AOI22X1 U990 ( .A(n333_1_), .B(n1774), .C(slice673_1_), .D(n1775), .Y(n1814)
         );
  NAND2X1 U991 ( .A(n1816), .B(n1817), .Y(result[7]) );
  AOI22X1 U992 ( .A(slice376_8_), .B(n1772), .C(slice356_8_), .D(n1773), .Y(
        n1817) );
  AOI22X1 U993 ( .A(slice673_8_), .B(n1774), .C(slice396_24_), .D(n1775), .Y(
        n1816) );
  NAND2X1 U994 ( .A(n1818), .B(n1819), .Y(result[79]) );
  AOI22X1 U995 ( .A(slice356_16_), .B(n1772), .C(slice396_16_), .D(n1773), .Y(
        n1819) );
  AOI22X1 U996 ( .A(slice753_16_), .B(n1774), .C(slice376_32_), .D(n1775), .Y(
        n1818) );
  NAND2X1 U997 ( .A(n1820), .B(n1821), .Y(result[78]) );
  AOI22X1 U998 ( .A(slice356_15_), .B(n1772), .C(slice396_15_), .D(n1773), .Y(
        n1821) );
  AOI22X1 U999 ( .A(slice753_15_), .B(n1774), .C(slice376_31_), .D(n1775), .Y(
        n1820) );
  NAND2X1 U1000 ( .A(n1822), .B(n1823), .Y(result[77]) );
  AOI22X1 U1001 ( .A(slice356_14_), .B(n1772), .C(slice396_14_), .D(n1773), 
        .Y(n1823) );
  AOI22X1 U1002 ( .A(slice753_14_), .B(n1774), .C(slice376_30_), .D(n1775), 
        .Y(n1822) );
  NAND2X1 U1003 ( .A(n1824), .B(n1825), .Y(result[76]) );
  AOI22X1 U1004 ( .A(slice356_13_), .B(n1772), .C(slice396_13_), .D(n1773), 
        .Y(n1825) );
  AOI22X1 U1005 ( .A(slice753_13_), .B(n1774), .C(slice376_29_), .D(n1775), 
        .Y(n1824) );
  NAND2X1 U1006 ( .A(n1826), .B(n1827), .Y(result[75]) );
  AOI22X1 U1007 ( .A(slice356_12_), .B(n1772), .C(slice396_12_), .D(n1773), 
        .Y(n1827) );
  AOI22X1 U1008 ( .A(slice753_12_), .B(n1774), .C(slice376_28_), .D(n1775), 
        .Y(n1826) );
  NAND2X1 U1009 ( .A(n1828), .B(n1829), .Y(result[74]) );
  AOI22X1 U1010 ( .A(slice356_11_), .B(n1772), .C(slice396_11_), .D(n1773), 
        .Y(n1829) );
  AOI22X1 U1011 ( .A(slice753_11_), .B(n1774), .C(slice376_27_), .D(n1775), 
        .Y(n1828) );
  NAND2X1 U1012 ( .A(n1830), .B(n1831), .Y(result[73]) );
  AOI22X1 U1013 ( .A(slice356_10_), .B(n1772), .C(slice396_10_), .D(n1773), 
        .Y(n1831) );
  AOI22X1 U1014 ( .A(slice753_10_), .B(n1774), .C(slice376_26_), .D(n1775), 
        .Y(n1830) );
  NAND2X1 U1015 ( .A(n1832), .B(n1833), .Y(result[72]) );
  AOI22X1 U1016 ( .A(slice356_9_), .B(n1772), .C(slice396_9_), .D(n1773), .Y(
        n1833) );
  AOI22X1 U1017 ( .A(slice753_9_), .B(n1774), .C(slice376_25_), .D(n1775), .Y(
        n1832) );
  NAND2X1 U1018 ( .A(n1834), .B(n1835), .Y(result[71]) );
  AOI22X1 U1019 ( .A(slice356_8_), .B(n1772), .C(slice396_8_), .D(n1773), .Y(
        n1835) );
  AOI22X1 U1020 ( .A(slice753_8_), .B(n1774), .C(slice376_24_), .D(n1775), .Y(
        n1834) );
  NAND2X1 U1021 ( .A(n1836), .B(n1837), .Y(result[70]) );
  AOI22X1 U1022 ( .A(slice356_7_), .B(n1772), .C(slice396_7_), .D(n1773), .Y(
        n1837) );
  AOI22X1 U1023 ( .A(slice753_7_), .B(n1774), .C(slice376_23_), .D(n1775), .Y(
        n1836) );
  NAND2X1 U1024 ( .A(n1838), .B(n1839), .Y(result[6]) );
  AOI22X1 U1025 ( .A(slice376_7_), .B(n1772), .C(slice356_7_), .D(n1773), .Y(
        n1839) );
  AOI22X1 U1026 ( .A(slice673_7_), .B(n1774), .C(slice396_23_), .D(n1775), .Y(
        n1838) );
  NAND2X1 U1027 ( .A(n1840), .B(n1841), .Y(result[69]) );
  AOI22X1 U1028 ( .A(slice356_6_), .B(n1772), .C(n213_6_), .D(n1773), .Y(n1841) );
  AOI22X1 U1029 ( .A(n328_6_), .B(n1774), .C(slice376_22_), .D(n1775), .Y(
        n1840) );
  NAND2X1 U1030 ( .A(n1842), .B(n1843), .Y(result[68]) );
  AOI22X1 U1031 ( .A(slice356_5_), .B(n1772), .C(slice396_5_), .D(n1773), .Y(
        n1843) );
  AOI22X1 U1032 ( .A(slice753_5_), .B(n1774), .C(slice376_21_), .D(n1775), .Y(
        n1842) );
  NAND2X1 U1033 ( .A(n1844), .B(n1845), .Y(result[67]) );
  AOI22X1 U1034 ( .A(n203_4_), .B(n1772), .C(slice396_4_), .D(n1773), .Y(n1845) );
  AOI22X1 U1035 ( .A(slice753_4_), .B(n1774), .C(slice376_20_), .D(n1775), .Y(
        n1844) );
  NAND2X1 U1036 ( .A(n1846), .B(n1847), .Y(result[66]) );
  AOI22X1 U1037 ( .A(slice356_3_), .B(n1772), .C(n213_3_), .D(n1773), .Y(n1847) );
  AOI22X1 U1038 ( .A(n328_3_), .B(n1774), .C(slice376_19_), .D(n1775), .Y(
        n1846) );
  NAND2X1 U1039 ( .A(n1848), .B(n1849), .Y(result[65]) );
  AOI22X1 U1040 ( .A(slice356_2_), .B(n1772), .C(n213_2_), .D(n1773), .Y(n1849) );
  AOI22X1 U1041 ( .A(n328_2_), .B(n1774), .C(slice376_18_), .D(n1775), .Y(
        n1848) );
  NAND2X1 U1042 ( .A(n1850), .B(n1851), .Y(result[64]) );
  AOI22X1 U1043 ( .A(n203_1_), .B(n1772), .C(n213_1_), .D(n1773), .Y(n1851) );
  AOI22X1 U1044 ( .A(n328_1_), .B(n1774), .C(slice376_17_), .D(n1775), .Y(
        n1850) );
  OAI21X1 U1045 ( .A(n1765), .B(n1853), .C(n1854), .Y(result[63]) );
  AOI22X1 U1046 ( .A(slice376_32_), .B(n1855), .C(slice396_32_), .D(n1772), 
        .Y(n1854) );
  OAI21X1 U1047 ( .A(n1765), .B(n1856), .C(n1857), .Y(result[62]) );
  AOI22X1 U1048 ( .A(slice376_31_), .B(n1855), .C(slice396_31_), .D(n1772), 
        .Y(n1857) );
  OAI21X1 U1049 ( .A(n1852), .B(n1858), .C(n1859), .Y(result[61]) );
  AOI22X1 U1050 ( .A(slice376_30_), .B(n1855), .C(slice396_30_), .D(n1772), 
        .Y(n1859) );
  OAI21X1 U1051 ( .A(n1852), .B(n1860), .C(n1861), .Y(result[60]) );
  AOI22X1 U1052 ( .A(slice376_29_), .B(n1855), .C(slice396_29_), .D(n1772), 
        .Y(n1861) );
  NAND2X1 U1053 ( .A(n1862), .B(n1863), .Y(result[5]) );
  AOI22X1 U1054 ( .A(n208_6_), .B(n1772), .C(slice356_6_), .D(n1773), .Y(n1863) );
  AOI22X1 U1055 ( .A(slice673_6_), .B(n1774), .C(slice396_22_), .D(n1775), .Y(
        n1862) );
  OAI21X1 U1056 ( .A(n1852), .B(n1864), .C(n1865), .Y(result[59]) );
  AOI22X1 U1057 ( .A(slice376_28_), .B(n1855), .C(slice396_28_), .D(n1772), 
        .Y(n1865) );
  OAI21X1 U1058 ( .A(n1852), .B(n1866), .C(n1867), .Y(result[58]) );
  AOI22X1 U1059 ( .A(slice376_27_), .B(n1855), .C(slice396_27_), .D(n1772), 
        .Y(n1867) );
  OAI21X1 U1060 ( .A(n1852), .B(n1868), .C(n1869), .Y(result[57]) );
  AOI22X1 U1061 ( .A(slice376_26_), .B(n1855), .C(slice396_26_), .D(n1772), 
        .Y(n1869) );
  OAI21X1 U1062 ( .A(n1852), .B(n1870), .C(n1871), .Y(result[56]) );
  AOI22X1 U1063 ( .A(slice376_25_), .B(n1855), .C(slice396_25_), .D(n1772), 
        .Y(n1871) );
  OAI21X1 U1064 ( .A(n1852), .B(n1872), .C(n1873), .Y(result[55]) );
  AOI22X1 U1065 ( .A(slice376_24_), .B(n1855), .C(slice396_24_), .D(n1772), 
        .Y(n1873) );
  OAI21X1 U1066 ( .A(n1852), .B(n1874), .C(n1875), .Y(result[54]) );
  AOI22X1 U1067 ( .A(slice376_23_), .B(n1855), .C(slice396_23_), .D(n1772), 
        .Y(n1875) );
  OAI21X1 U1068 ( .A(n1852), .B(n1876), .C(n1877), .Y(result[53]) );
  AOI22X1 U1069 ( .A(slice376_22_), .B(n1855), .C(slice396_22_), .D(n1772), 
        .Y(n1877) );
  OAI21X1 U1070 ( .A(n1852), .B(n1878), .C(n1879), .Y(result[52]) );
  AOI22X1 U1071 ( .A(slice376_21_), .B(n1855), .C(slice396_21_), .D(n1772), 
        .Y(n1879) );
  OAI21X1 U1072 ( .A(n1852), .B(n1880), .C(n1881), .Y(result[51]) );
  AOI22X1 U1073 ( .A(slice376_20_), .B(n1855), .C(slice396_20_), .D(n1772), 
        .Y(n1881) );
  OAI21X1 U1074 ( .A(n1852), .B(n1882), .C(n1883), .Y(result[50]) );
  AOI22X1 U1075 ( .A(slice376_19_), .B(n1855), .C(slice396_19_), .D(n1772), 
        .Y(n1883) );
  NAND2X1 U1076 ( .A(n1884), .B(n1885), .Y(result[4]) );
  AOI22X1 U1077 ( .A(slice376_5_), .B(n1772), .C(slice356_5_), .D(n1773), .Y(
        n1885) );
  AOI22X1 U1078 ( .A(slice673_5_), .B(n1774), .C(slice396_21_), .D(n1775), .Y(
        n1884) );
  OAI21X1 U1079 ( .A(n1852), .B(n1886), .C(n1887), .Y(result[49]) );
  AOI22X1 U1080 ( .A(slice376_18_), .B(n1855), .C(slice396_18_), .D(n1772), 
        .Y(n1887) );
  OAI21X1 U1081 ( .A(n1765), .B(n1888), .C(n1889), .Y(result[48]) );
  AOI22X1 U1082 ( .A(slice376_17_), .B(n1855), .C(slice396_17_), .D(n1772), 
        .Y(n1889) );
  NAND2X1 U1083 ( .A(n1890), .B(n1891), .Y(n1855) );
  NAND2X1 U1084 ( .A(n1892), .B(n1893), .Y(result[47]) );
  AOI22X1 U1085 ( .A(slice396_16_), .B(n1772), .C(slice376_16_), .D(n1773), 
        .Y(n1893) );
  AOI22X1 U1086 ( .A(slice455_16_), .B(n1774), .C(slice773_16_), .D(n1775), 
        .Y(n1892) );
  NAND2X1 U1087 ( .A(n1894), .B(n1895), .Y(result[46]) );
  AOI22X1 U1088 ( .A(slice396_15_), .B(n1772), .C(slice376_15_), .D(n1773), 
        .Y(n1895) );
  AOI22X1 U1089 ( .A(slice455_15_), .B(n1774), .C(slice773_15_), .D(n1775), 
        .Y(n1894) );
  NAND2X1 U1090 ( .A(n1896), .B(n1897), .Y(result[45]) );
  AOI22X1 U1091 ( .A(slice396_14_), .B(n1772), .C(slice376_14_), .D(n1773), 
        .Y(n1897) );
  AOI22X1 U1092 ( .A(slice455_14_), .B(n1774), .C(slice773_14_), .D(n1775), 
        .Y(n1896) );
  NAND2X1 U1093 ( .A(n1898), .B(n1899), .Y(result[44]) );
  AOI22X1 U1094 ( .A(slice396_13_), .B(n1772), .C(slice376_13_), .D(n1773), 
        .Y(n1899) );
  AOI22X1 U1095 ( .A(slice455_13_), .B(n1774), .C(slice773_13_), .D(n1775), 
        .Y(n1898) );
  NAND2X1 U1096 ( .A(n1900), .B(n1901), .Y(result[43]) );
  AOI22X1 U1097 ( .A(slice396_12_), .B(n1772), .C(slice376_12_), .D(n1773), 
        .Y(n1901) );
  AOI22X1 U1098 ( .A(slice455_12_), .B(n1774), .C(slice773_12_), .D(n1775), 
        .Y(n1900) );
  NAND2X1 U1099 ( .A(n1902), .B(n1903), .Y(result[42]) );
  AOI22X1 U1100 ( .A(slice396_11_), .B(n1772), .C(slice376_11_), .D(n1773), 
        .Y(n1903) );
  AOI22X1 U1101 ( .A(slice455_11_), .B(n1774), .C(slice773_11_), .D(n1775), 
        .Y(n1902) );
  NAND2X1 U1102 ( .A(n1904), .B(n1905), .Y(result[41]) );
  AOI22X1 U1103 ( .A(slice396_10_), .B(n1772), .C(n1773), .D(slice376_10_), 
        .Y(n1905) );
  AOI22X1 U1104 ( .A(slice455_10_), .B(n1774), .C(slice773_10_), .D(n1775), 
        .Y(n1904) );
  NAND2X1 U1105 ( .A(n1906), .B(n1907), .Y(result[40]) );
  AOI22X1 U1106 ( .A(slice396_9_), .B(n1772), .C(slice376_9_), .D(n1773), .Y(
        n1907) );
  AOI22X1 U1107 ( .A(slice455_9_), .B(n1774), .C(slice773_9_), .D(n1775), .Y(
        n1906) );
  NAND2X1 U1108 ( .A(n1908), .B(n1909), .Y(result[3]) );
  AOI22X1 U1109 ( .A(slice376_4_), .B(n1772), .C(n203_4_), .D(n1773), .Y(n1909) );
  AOI22X1 U1110 ( .A(slice673_4_), .B(n1774), .C(slice396_20_), .D(n1775), .Y(
        n1908) );
  NAND2X1 U1111 ( .A(n1910), .B(n1911), .Y(result[39]) );
  AOI22X1 U1112 ( .A(slice396_8_), .B(n1772), .C(slice376_8_), .D(n1773), .Y(
        n1911) );
  AOI22X1 U1113 ( .A(slice455_8_), .B(n1774), .C(slice773_8_), .D(n1775), .Y(
        n1910) );
  NAND2X1 U1114 ( .A(n1912), .B(n1913), .Y(result[38]) );
  AOI22X1 U1115 ( .A(slice396_7_), .B(n1772), .C(slice376_7_), .D(n1773), .Y(
        n1913) );
  AOI22X1 U1116 ( .A(slice455_7_), .B(n1774), .C(slice773_7_), .D(n1775), .Y(
        n1912) );
  NAND2X1 U1117 ( .A(n1914), .B(n1915), .Y(result[37]) );
  AOI22X1 U1118 ( .A(n213_6_), .B(n1772), .C(n208_6_), .D(n1773), .Y(n1915) );
  AOI22X1 U1119 ( .A(n228_6_), .B(n1774), .C(n333_6_), .D(n1775), .Y(n1914) );
  NAND2X1 U1120 ( .A(n1916), .B(n1917), .Y(result[36]) );
  AOI22X1 U1121 ( .A(slice396_5_), .B(n1772), .C(slice376_5_), .D(n1773), .Y(
        n1917) );
  AOI22X1 U1122 ( .A(slice455_5_), .B(n1774), .C(slice773_5_), .D(n1775), .Y(
        n1916) );
  NAND2X1 U1123 ( .A(n1918), .B(n1919), .Y(result[35]) );
  AOI22X1 U1124 ( .A(slice396_4_), .B(n1772), .C(slice376_4_), .D(n1773), .Y(
        n1919) );
  AOI22X1 U1125 ( .A(slice455_4_), .B(n1774), .C(slice773_4_), .D(n1775), .Y(
        n1918) );
  NAND2X1 U1126 ( .A(n1920), .B(n1921), .Y(result[34]) );
  AOI22X1 U1127 ( .A(n213_3_), .B(n1772), .C(n208_3_), .D(n1773), .Y(n1921) );
  AOI22X1 U1128 ( .A(n228_3_), .B(n1774), .C(n333_3_), .D(n1775), .Y(n1920) );
  NAND2X1 U1129 ( .A(n1922), .B(n1923), .Y(result[33]) );
  AOI22X1 U1130 ( .A(n213_2_), .B(n1772), .C(n208_2_), .D(n1773), .Y(n1923) );
  AOI22X1 U1131 ( .A(n228_2_), .B(n1774), .C(n333_2_), .D(n1775), .Y(n1922) );
  NAND2X1 U1132 ( .A(n1924), .B(n1925), .Y(result[32]) );
  AOI22X1 U1133 ( .A(n213_1_), .B(n1772), .C(n208_1_), .D(n1773), .Y(n1925) );
  AOI22X1 U1134 ( .A(n228_1_), .B(n1774), .C(n333_1_), .D(n1775), .Y(n1924) );
  OAI21X1 U1135 ( .A(n1890), .B(n1853), .C(n1926), .Y(result[31]) );
  AOI22X1 U1136 ( .A(n1927), .B(slice455_16_), .C(slice376_32_), .D(n1772), 
        .Y(n1926) );
  INVX1 U1137 ( .A(slice693_16_), .Y(n1853) );
  OAI21X1 U1138 ( .A(n1890), .B(n1856), .C(n1928), .Y(result[30]) );
  AOI22X1 U1139 ( .A(n1927), .B(slice455_15_), .C(slice376_31_), .D(n1772), 
        .Y(n1928) );
  INVX1 U1140 ( .A(slice693_15_), .Y(n1856) );
  NAND2X1 U1141 ( .A(n1929), .B(n1930), .Y(result[2]) );
  AOI22X1 U1142 ( .A(n208_3_), .B(n1772), .C(slice356_3_), .D(n1773), .Y(n1930) );
  AOI22X1 U1143 ( .A(slice673_3_), .B(n1774), .C(slice396_19_), .D(n1775), .Y(
        n1929) );
  OAI21X1 U1144 ( .A(n1890), .B(n1858), .C(n1931), .Y(result[29]) );
  AOI22X1 U1145 ( .A(n1927), .B(slice455_14_), .C(slice376_30_), .D(n1772), 
        .Y(n1931) );
  INVX1 U1146 ( .A(slice693_14_), .Y(n1858) );
  OAI21X1 U1147 ( .A(n1890), .B(n1860), .C(n1932), .Y(result[28]) );
  AOI22X1 U1148 ( .A(n1927), .B(slice455_13_), .C(slice376_29_), .D(n1772), 
        .Y(n1932) );
  INVX1 U1149 ( .A(slice693_13_), .Y(n1860) );
  OAI21X1 U1150 ( .A(n1890), .B(n1864), .C(n1933), .Y(result[27]) );
  AOI22X1 U1151 ( .A(n1927), .B(slice455_12_), .C(slice376_28_), .D(n1772), 
        .Y(n1933) );
  INVX1 U1152 ( .A(slice693_12_), .Y(n1864) );
  OAI21X1 U1153 ( .A(n1890), .B(n1866), .C(n1934), .Y(result[26]) );
  AOI22X1 U1154 ( .A(n1927), .B(slice455_11_), .C(slice376_27_), .D(n1772), 
        .Y(n1934) );
  INVX1 U1155 ( .A(slice693_11_), .Y(n1866) );
  OAI21X1 U1156 ( .A(n1890), .B(n1868), .C(n1935), .Y(result[25]) );
  AOI22X1 U1157 ( .A(n1927), .B(slice455_10_), .C(slice376_26_), .D(n1772), 
        .Y(n1935) );
  INVX1 U1158 ( .A(slice693_10_), .Y(n1868) );
  OAI21X1 U1159 ( .A(n1890), .B(n1870), .C(n1936), .Y(result[24]) );
  AOI22X1 U1160 ( .A(n1927), .B(slice455_9_), .C(slice376_25_), .D(n1772), .Y(
        n1936) );
  INVX1 U1161 ( .A(slice693_9_), .Y(n1870) );
  OAI21X1 U1162 ( .A(n1890), .B(n1872), .C(n1937), .Y(result[23]) );
  AOI22X1 U1163 ( .A(n1927), .B(slice455_8_), .C(slice376_24_), .D(n1772), .Y(
        n1937) );
  INVX1 U1164 ( .A(slice693_8_), .Y(n1872) );
  OAI21X1 U1165 ( .A(n1890), .B(n1874), .C(n1938), .Y(result[22]) );
  AOI22X1 U1166 ( .A(n1927), .B(slice455_7_), .C(slice376_23_), .D(n1772), .Y(
        n1938) );
  INVX1 U1167 ( .A(slice693_7_), .Y(n1874) );
  OAI21X1 U1168 ( .A(n1890), .B(n1876), .C(n1939), .Y(result[21]) );
  AOI22X1 U1169 ( .A(n1927), .B(n228_6_), .C(slice376_22_), .D(n1772), .Y(
        n1939) );
  INVX1 U1170 ( .A(n313_6_), .Y(n1876) );
  OAI21X1 U1171 ( .A(n1890), .B(n1878), .C(n1940), .Y(result[20]) );
  AOI22X1 U1172 ( .A(n1927), .B(slice455_5_), .C(slice376_21_), .D(n1772), .Y(
        n1940) );
  INVX1 U1173 ( .A(slice693_5_), .Y(n1878) );
  NAND2X1 U1174 ( .A(n1941), .B(n1942), .Y(result[1]) );
  AOI22X1 U1175 ( .A(n208_2_), .B(n1772), .C(slice356_2_), .D(n1773), .Y(n1942) );
  AOI22X1 U1176 ( .A(slice673_2_), .B(n1774), .C(slice396_18_), .D(n1775), .Y(
        n1941) );
  OAI21X1 U1177 ( .A(n1890), .B(n1880), .C(n1943), .Y(result[19]) );
  AOI22X1 U1178 ( .A(n1927), .B(slice455_4_), .C(slice376_20_), .D(n1772), .Y(
        n1943) );
  INVX1 U1179 ( .A(slice693_4_), .Y(n1880) );
  OAI21X1 U1180 ( .A(n1890), .B(n1882), .C(n1944), .Y(result[18]) );
  AOI22X1 U1181 ( .A(n1927), .B(n228_3_), .C(slice376_19_), .D(n1772), .Y(
        n1944) );
  INVX1 U1182 ( .A(n313_3_), .Y(n1882) );
  OAI21X1 U1183 ( .A(n1890), .B(n1886), .C(n1945), .Y(result[17]) );
  AOI22X1 U1184 ( .A(n1927), .B(n228_2_), .C(slice376_18_), .D(n1772), .Y(
        n1945) );
  INVX1 U1185 ( .A(n313_2_), .Y(n1886) );
  OAI21X1 U1186 ( .A(n1890), .B(n1888), .C(n1946), .Y(result[16]) );
  AOI22X1 U1187 ( .A(n1927), .B(n228_1_), .C(slice376_17_), .D(n1772), .Y(
        n1946) );
  INVX1 U1188 ( .A(n1947), .Y(n1927) );
  OAI21X1 U1189 ( .A(n1948), .B(n1949), .C(n1950), .Y(n1947) );
  INVX1 U1190 ( .A(n313_1_), .Y(n1888) );
  NAND2X1 U1191 ( .A(n1951), .B(n1952), .Y(result[15]) );
  AOI22X1 U1192 ( .A(slice376_16_), .B(n1772), .C(slice356_16_), .D(n1773), 
        .Y(n1952) );
  AOI22X1 U1193 ( .A(slice673_16_), .B(n1774), .C(slice396_32_), .D(n1775), 
        .Y(n1951) );
  NAND2X1 U1194 ( .A(n1953), .B(n1954), .Y(result[14]) );
  AOI22X1 U1195 ( .A(slice376_15_), .B(n1772), .C(slice356_15_), .D(n1773), 
        .Y(n1954) );
  AOI22X1 U1196 ( .A(slice673_15_), .B(n1774), .C(slice396_31_), .D(n1775), 
        .Y(n1953) );
  NAND2X1 U1197 ( .A(n1955), .B(n1956), .Y(result[13]) );
  AOI22X1 U1198 ( .A(slice376_14_), .B(n1772), .C(slice356_14_), .D(n1773), 
        .Y(n1956) );
  AOI22X1 U1199 ( .A(slice673_14_), .B(n1774), .C(slice396_30_), .D(n1775), 
        .Y(n1955) );
  NAND2X1 U1200 ( .A(n1957), .B(n1958), .Y(result[12]) );
  AOI22X1 U1201 ( .A(slice376_13_), .B(n1772), .C(slice356_13_), .D(n1773), 
        .Y(n1958) );
  AOI22X1 U1202 ( .A(slice673_13_), .B(n1774), .C(slice396_29_), .D(n1775), 
        .Y(n1957) );
  OAI21X1 U1203 ( .A(n1852), .B(n1959), .C(n1960), .Y(result[127]) );
  AOI22X1 U1204 ( .A(slice693_16_), .B(n1764), .C(slice396_32_), .D(n1774), 
        .Y(n1960) );
  INVX1 U1205 ( .A(slice753_16_), .Y(n1959) );
  OAI21X1 U1206 ( .A(n1852), .B(n1961), .C(n1962), .Y(result[126]) );
  AOI22X1 U1207 ( .A(slice693_15_), .B(n1764), .C(slice396_31_), .D(n1774), 
        .Y(n1962) );
  INVX1 U1208 ( .A(slice753_15_), .Y(n1961) );
  OAI21X1 U1209 ( .A(n1852), .B(n1963), .C(n1964), .Y(result[125]) );
  AOI22X1 U1210 ( .A(slice693_14_), .B(n1764), .C(slice396_30_), .D(n1774), 
        .Y(n1964) );
  INVX1 U1211 ( .A(slice753_14_), .Y(n1963) );
  OAI21X1 U1212 ( .A(n1852), .B(n1965), .C(n1966), .Y(result[124]) );
  AOI22X1 U1213 ( .A(slice693_13_), .B(n1764), .C(slice396_29_), .D(n1774), 
        .Y(n1966) );
  INVX1 U1214 ( .A(slice753_13_), .Y(n1965) );
  OAI21X1 U1215 ( .A(n1852), .B(n1967), .C(n1968), .Y(result[123]) );
  AOI22X1 U1216 ( .A(slice693_12_), .B(n1764), .C(slice396_28_), .D(n1774), 
        .Y(n1968) );
  INVX1 U1217 ( .A(slice753_12_), .Y(n1967) );
  OAI21X1 U1218 ( .A(n1852), .B(n1969), .C(n1970), .Y(result[122]) );
  AOI22X1 U1219 ( .A(slice693_11_), .B(n1764), .C(slice396_27_), .D(n1774), 
        .Y(n1970) );
  INVX1 U1220 ( .A(slice753_11_), .Y(n1969) );
  OAI21X1 U1221 ( .A(n1852), .B(n1971), .C(n1972), .Y(result[121]) );
  AOI22X1 U1222 ( .A(slice693_10_), .B(n1764), .C(slice396_26_), .D(n1774), 
        .Y(n1972) );
  INVX1 U1223 ( .A(slice753_10_), .Y(n1971) );
  OAI21X1 U1224 ( .A(n1852), .B(n1973), .C(n1974), .Y(result[120]) );
  AOI22X1 U1225 ( .A(slice693_9_), .B(n1764), .C(slice396_25_), .D(n1774), .Y(
        n1974) );
  INVX1 U1226 ( .A(slice753_9_), .Y(n1973) );
  NAND2X1 U1227 ( .A(n1975), .B(n1976), .Y(result[11]) );
  AOI22X1 U1228 ( .A(slice376_12_), .B(n1772), .C(slice356_12_), .D(n1773), 
        .Y(n1976) );
  AOI22X1 U1229 ( .A(slice673_12_), .B(n1774), .C(slice396_28_), .D(n1775), 
        .Y(n1975) );
  OAI21X1 U1230 ( .A(n1852), .B(n1977), .C(n1978), .Y(result[119]) );
  AOI22X1 U1231 ( .A(slice693_8_), .B(n1764), .C(slice396_24_), .D(n1774), .Y(
        n1978) );
  INVX1 U1232 ( .A(slice753_8_), .Y(n1977) );
  OAI21X1 U1233 ( .A(n1852), .B(n1979), .C(n1980), .Y(result[118]) );
  AOI22X1 U1234 ( .A(slice693_7_), .B(n1764), .C(slice396_23_), .D(n1774), .Y(
        n1980) );
  INVX1 U1235 ( .A(slice753_7_), .Y(n1979) );
  OAI21X1 U1236 ( .A(n1852), .B(n1981), .C(n1982), .Y(result[117]) );
  AOI22X1 U1237 ( .A(n313_6_), .B(n1764), .C(slice396_22_), .D(n1774), .Y(
        n1982) );
  INVX1 U1238 ( .A(n328_6_), .Y(n1981) );
  OAI21X1 U1239 ( .A(n1852), .B(n1983), .C(n1984), .Y(result[116]) );
  AOI22X1 U1240 ( .A(slice693_5_), .B(n1764), .C(slice396_21_), .D(n1774), .Y(
        n1984) );
  INVX1 U1241 ( .A(slice753_5_), .Y(n1983) );
  OAI21X1 U1242 ( .A(n1765), .B(n1985), .C(n1986), .Y(result[115]) );
  AOI22X1 U1243 ( .A(slice693_4_), .B(n1764), .C(slice396_20_), .D(n1774), .Y(
        n1986) );
  INVX1 U1244 ( .A(slice753_4_), .Y(n1985) );
  OAI21X1 U1245 ( .A(n1765), .B(n1987), .C(n1988), .Y(result[114]) );
  AOI22X1 U1246 ( .A(n313_3_), .B(n1764), .C(slice396_19_), .D(n1774), .Y(
        n1988) );
  INVX1 U1247 ( .A(n328_3_), .Y(n1987) );
  OAI21X1 U1248 ( .A(n1765), .B(n1989), .C(n1990), .Y(result[113]) );
  AOI22X1 U1249 ( .A(n313_2_), .B(n1764), .C(slice396_18_), .D(n1774), .Y(
        n1990) );
  INVX1 U1250 ( .A(n328_2_), .Y(n1989) );
  OAI21X1 U1251 ( .A(n1852), .B(n1991), .C(n1992), .Y(result[112]) );
  AOI22X1 U1252 ( .A(n313_1_), .B(n1764), .C(slice396_17_), .D(n1774), .Y(
        n1992) );
  INVX1 U1253 ( .A(n328_1_), .Y(n1991) );
  INVX1 U1254 ( .A(n1993), .Y(result[111]) );
  AOI22X1 U1255 ( .A(slice416_16_), .B(n1764), .C(slice793_16_), .D(n1778), 
        .Y(n1993) );
  INVX1 U1256 ( .A(n1994), .Y(result[110]) );
  AOI22X1 U1257 ( .A(slice416_15_), .B(n1764), .C(slice793_15_), .D(n1778), 
        .Y(n1994) );
  NAND2X1 U1258 ( .A(n1995), .B(n1996), .Y(result[10]) );
  AOI22X1 U1259 ( .A(slice376_11_), .B(n1772), .C(slice356_11_), .D(n1773), 
        .Y(n1996) );
  AOI22X1 U1260 ( .A(slice673_11_), .B(n1774), .C(slice396_27_), .D(n1775), 
        .Y(n1995) );
  INVX1 U1261 ( .A(n1997), .Y(result[109]) );
  AOI22X1 U1262 ( .A(slice416_14_), .B(n1764), .C(slice793_14_), .D(n1778), 
        .Y(n1997) );
  INVX1 U1263 ( .A(n1998), .Y(result[108]) );
  AOI22X1 U1264 ( .A(slice416_13_), .B(n1764), .C(slice793_13_), .D(n1778), 
        .Y(n1998) );
  INVX1 U1265 ( .A(n1999), .Y(result[107]) );
  AOI22X1 U1266 ( .A(slice416_12_), .B(n1764), .C(slice793_12_), .D(n1778), 
        .Y(n1999) );
  INVX1 U1267 ( .A(n2000), .Y(result[106]) );
  AOI22X1 U1268 ( .A(slice416_11_), .B(n1764), .C(slice793_11_), .D(n1778), 
        .Y(n2000) );
  INVX1 U1269 ( .A(n2001), .Y(result[105]) );
  AOI22X1 U1270 ( .A(slice416_10_), .B(n1764), .C(slice793_10_), .D(n1778), 
        .Y(n2001) );
  INVX1 U1271 ( .A(n2002), .Y(result[104]) );
  AOI22X1 U1272 ( .A(slice416_9_), .B(n1764), .C(slice793_9_), .D(n1778), .Y(
        n2002) );
  INVX1 U1273 ( .A(n2003), .Y(result[103]) );
  AOI22X1 U1274 ( .A(slice416_8_), .B(n1764), .C(slice793_8_), .D(n1778), .Y(
        n2003) );
  INVX1 U1275 ( .A(n2004), .Y(result[102]) );
  AOI22X1 U1276 ( .A(slice416_7_), .B(n1764), .C(slice793_7_), .D(n1778), .Y(
        n2004) );
  INVX1 U1277 ( .A(n2005), .Y(result[101]) );
  AOI22X1 U1278 ( .A(n218_6_), .B(n1764), .C(n338_6_), .D(n1778), .Y(n2005) );
  INVX1 U1279 ( .A(n2006), .Y(result[100]) );
  AOI22X1 U1280 ( .A(slice416_5_), .B(n1764), .C(slice793_5_), .D(n1778), .Y(
        n2006) );
  NAND2X1 U1281 ( .A(n1765), .B(n1890), .Y(n1778) );
  NAND2X1 U1282 ( .A(n1891), .B(n2007), .Y(n1777) );
  NAND2X1 U1283 ( .A(n2008), .B(n2009), .Y(result[0]) );
  AOI22X1 U1284 ( .A(n208_1_), .B(n1772), .C(n203_1_), .D(n1773), .Y(n2009) );
  NAND2X1 U1285 ( .A(n1950), .B(n1948), .Y(n1891) );
  NAND3X1 U1286 ( .A(n2010), .B(n2011), .C(n1948), .Y(n2007) );
  NOR2X1 U1287 ( .A(n2012), .B(ctrl_ww[0]), .Y(n1948) );
  AOI22X1 U1288 ( .A(slice673_1_), .B(n1774), .C(slice396_17_), .D(n1775), .Y(
        n2008) );
  NAND2X1 U1289 ( .A(n1949), .B(n1950), .Y(n1852) );
  NOR2X1 U1290 ( .A(n2011), .B(n2013), .Y(n1950) );
  NAND3X1 U1291 ( .A(n2010), .B(n2011), .C(n1949), .Y(n1890) );
  NOR2X1 U1292 ( .A(ctrl_ww[1]), .B(ctrl_ww[0]), .Y(n1949) );
  INVX1 U1293 ( .A(n2013), .Y(n2010) );
  NAND3X1 U1294 ( .A(alu_op[3]), .B(alu_op[1]), .C(n2014), .Y(n2013) );
  NOR2X1 U1295 ( .A(alu_op[4]), .B(n2015), .Y(n2014) );
  INVX1 U1296 ( .A(alu_op[0]), .Y(n2015) );
  INVX1 U1297 ( .A(n2016), .Y(U69_U9_Z_9) );
  AOI22X1 U1298 ( .A(n1768), .B(reg_A[70]), .C(n2018), .D(reg_A[22]), .Y(n2016) );
  INVX1 U1299 ( .A(n2019), .Y(U69_U9_Z_8) );
  AOI22X1 U1300 ( .A(n1768), .B(reg_A[71]), .C(n1767), .D(reg_A[23]), .Y(n2019) );
  OAI21X1 U1301 ( .A(n2020), .B(n2021), .C(n2022), .Y(U69_U9_Z_7) );
  AOI22X1 U1302 ( .A(reg_A[24]), .B(n2023), .C(reg_A[72]), .D(n1768), .Y(n2022) );
  INVX1 U1303 ( .A(reg_A[32]), .Y(n2021) );
  OAI21X1 U1304 ( .A(n2020), .B(n2024), .C(n2025), .Y(U69_U9_Z_6) );
  AOI22X1 U1305 ( .A(reg_A[25]), .B(n2023), .C(reg_A[73]), .D(n1768), .Y(n2025) );
  INVX1 U1306 ( .A(reg_A[33]), .Y(n2024) );
  OAI21X1 U1307 ( .A(n2020), .B(n2026), .C(n2027), .Y(U69_U9_Z_5) );
  AOI22X1 U1308 ( .A(reg_A[26]), .B(n2023), .C(reg_A[74]), .D(n2017), .Y(n2027) );
  INVX1 U1309 ( .A(reg_A[34]), .Y(n2026) );
  OAI21X1 U1310 ( .A(n2020), .B(n2028), .C(n2029), .Y(U69_U9_Z_4) );
  AOI22X1 U1311 ( .A(reg_A[27]), .B(n2023), .C(reg_A[75]), .D(n1768), .Y(n2029) );
  INVX1 U1312 ( .A(reg_A[35]), .Y(n2028) );
  OAI21X1 U1313 ( .A(n2020), .B(n2030), .C(n2031), .Y(U69_U9_Z_3) );
  AOI22X1 U1314 ( .A(reg_A[28]), .B(n2023), .C(reg_A[76]), .D(n2017), .Y(n2031) );
  INVX1 U1315 ( .A(reg_A[36]), .Y(n2030) );
  OAI21X1 U1316 ( .A(n2020), .B(n2032), .C(n2033), .Y(U69_U9_Z_2) );
  AOI22X1 U1317 ( .A(reg_A[29]), .B(n2023), .C(reg_A[77]), .D(n1768), .Y(n2033) );
  INVX1 U1318 ( .A(reg_A[37]), .Y(n2032) );
  INVX1 U1319 ( .A(n2034), .Y(U69_U9_Z_15) );
  AOI22X1 U1320 ( .A(n1768), .B(reg_A[64]), .C(n1767), .D(reg_A[16]), .Y(n2034) );
  INVX1 U1321 ( .A(n2035), .Y(U69_U9_Z_14) );
  AOI22X1 U1322 ( .A(n1768), .B(reg_A[65]), .C(n1767), .D(reg_A[17]), .Y(n2035) );
  INVX1 U1323 ( .A(n2036), .Y(U69_U9_Z_13) );
  AOI22X1 U1324 ( .A(n1768), .B(reg_A[66]), .C(n2018), .D(reg_A[18]), .Y(n2036) );
  INVX1 U1325 ( .A(n2037), .Y(U69_U9_Z_12) );
  AOI22X1 U1326 ( .A(n1768), .B(reg_A[67]), .C(n2018), .D(reg_A[19]), .Y(n2037) );
  INVX1 U1327 ( .A(n2038), .Y(U69_U9_Z_11) );
  AOI22X1 U1328 ( .A(n1768), .B(reg_A[68]), .C(n1767), .D(reg_A[20]), .Y(n2038) );
  INVX1 U1329 ( .A(n2039), .Y(U69_U9_Z_10) );
  AOI22X1 U1330 ( .A(n1768), .B(reg_A[69]), .C(n1767), .D(reg_A[21]), .Y(n2039) );
  OAI21X1 U1331 ( .A(n2020), .B(n2040), .C(n2041), .Y(U69_U9_Z_1) );
  AOI22X1 U1332 ( .A(reg_A[30]), .B(n2023), .C(reg_A[78]), .D(n1768), .Y(n2041) );
  INVX1 U1333 ( .A(reg_A[38]), .Y(n2040) );
  OAI21X1 U1334 ( .A(n2020), .B(n2042), .C(n2043), .Y(U69_U9_Z_0) );
  AOI22X1 U1335 ( .A(reg_A[31]), .B(n2023), .C(reg_A[79]), .D(n2017), .Y(n2043) );
  INVX1 U1336 ( .A(reg_A[39]), .Y(n2042) );
  INVX1 U1337 ( .A(n2044), .Y(U69_U8_Z_9) );
  AOI22X1 U1338 ( .A(n1768), .B(reg_B[102]), .C(n2018), .D(reg_B[118]), .Y(
        n2044) );
  INVX1 U1339 ( .A(n2045), .Y(U69_U8_Z_8) );
  AOI22X1 U1340 ( .A(n1768), .B(reg_B[103]), .C(n1767), .D(reg_B[119]), .Y(
        n2045) );
  NAND2X1 U1341 ( .A(n2046), .B(n2047), .Y(U69_U8_Z_7) );
  AOI22X1 U1342 ( .A(reg_B[120]), .B(n1767), .C(reg_B[104]), .D(n1768), .Y(
        n2047) );
  AOI22X1 U1343 ( .A(reg_B[56]), .B(n1766), .C(reg_B[16]), .D(n2049), .Y(n2046) );
  NAND2X1 U1344 ( .A(n2050), .B(n2051), .Y(U69_U8_Z_6) );
  AOI22X1 U1345 ( .A(reg_B[121]), .B(n1767), .C(reg_B[105]), .D(n1768), .Y(
        n2051) );
  AOI22X1 U1346 ( .A(reg_B[57]), .B(n1766), .C(reg_B[17]), .D(n2049), .Y(n2050) );
  NAND2X1 U1347 ( .A(n2052), .B(n2053), .Y(U69_U8_Z_5) );
  AOI22X1 U1348 ( .A(reg_B[122]), .B(n1767), .C(reg_B[106]), .D(n1768), .Y(
        n2053) );
  AOI22X1 U1349 ( .A(reg_B[58]), .B(n1766), .C(reg_B[18]), .D(n2049), .Y(n2052) );
  NAND2X1 U1350 ( .A(n2054), .B(n2055), .Y(U69_U8_Z_4) );
  AOI22X1 U1351 ( .A(reg_B[123]), .B(n1767), .C(reg_B[107]), .D(n1768), .Y(
        n2055) );
  AOI22X1 U1352 ( .A(reg_B[59]), .B(n1766), .C(reg_B[19]), .D(n2049), .Y(n2054) );
  NAND2X1 U1353 ( .A(n2056), .B(n2057), .Y(U69_U8_Z_3) );
  AOI22X1 U1354 ( .A(reg_B[124]), .B(n1767), .C(reg_B[108]), .D(n1768), .Y(
        n2057) );
  AOI22X1 U1355 ( .A(reg_B[60]), .B(n1766), .C(reg_B[20]), .D(n2049), .Y(n2056) );
  NAND2X1 U1356 ( .A(n2058), .B(n2059), .Y(U69_U8_Z_2) );
  AOI22X1 U1357 ( .A(reg_B[125]), .B(n1767), .C(reg_B[109]), .D(n1768), .Y(
        n2059) );
  AOI22X1 U1358 ( .A(reg_B[61]), .B(n1766), .C(reg_B[21]), .D(n2049), .Y(n2058) );
  INVX1 U1359 ( .A(n2060), .Y(U69_U8_Z_15) );
  AOI22X1 U1360 ( .A(n1768), .B(reg_B[96]), .C(n1767), .D(reg_B[112]), .Y(
        n2060) );
  INVX1 U1361 ( .A(n2061), .Y(U69_U8_Z_14) );
  AOI22X1 U1362 ( .A(n1768), .B(reg_B[97]), .C(n1767), .D(reg_B[113]), .Y(
        n2061) );
  INVX1 U1363 ( .A(n2062), .Y(U69_U8_Z_13) );
  AOI22X1 U1364 ( .A(n1768), .B(reg_B[98]), .C(n1767), .D(reg_B[114]), .Y(
        n2062) );
  INVX1 U1365 ( .A(n2063), .Y(U69_U8_Z_12) );
  AOI22X1 U1366 ( .A(n1768), .B(reg_B[99]), .C(n2018), .D(reg_B[115]), .Y(
        n2063) );
  INVX1 U1367 ( .A(n2064), .Y(U69_U8_Z_11) );
  AOI22X1 U1368 ( .A(n1768), .B(reg_B[100]), .C(n1767), .D(reg_B[116]), .Y(
        n2064) );
  INVX1 U1369 ( .A(n2065), .Y(U69_U8_Z_10) );
  AOI22X1 U1370 ( .A(n1768), .B(reg_B[101]), .C(n1767), .D(reg_B[117]), .Y(
        n2065) );
  NAND2X1 U1371 ( .A(n2066), .B(n2067), .Y(U69_U8_Z_1) );
  AOI22X1 U1372 ( .A(reg_B[126]), .B(n1767), .C(reg_B[110]), .D(n1768), .Y(
        n2067) );
  AOI22X1 U1373 ( .A(reg_B[62]), .B(n1766), .C(reg_B[22]), .D(n2049), .Y(n2066) );
  NAND2X1 U1374 ( .A(n2068), .B(n2069), .Y(U69_U8_Z_0) );
  AOI22X1 U1375 ( .A(reg_B[127]), .B(n1767), .C(reg_B[111]), .D(n1768), .Y(
        n2069) );
  AOI22X1 U1376 ( .A(reg_B[63]), .B(n1766), .C(reg_B[23]), .D(n2049), .Y(n2068) );
  INVX1 U1377 ( .A(n2070), .Y(U69_U7_Z_9) );
  AOI22X1 U1378 ( .A(n1768), .B(reg_A[102]), .C(n1767), .D(reg_A[118]), .Y(
        n2070) );
  INVX1 U1379 ( .A(n2071), .Y(U69_U7_Z_8) );
  AOI22X1 U1380 ( .A(n1768), .B(reg_A[103]), .C(n2018), .D(reg_A[119]), .Y(
        n2071) );
  NAND2X1 U1381 ( .A(n2072), .B(n2073), .Y(U69_U7_Z_7) );
  AOI22X1 U1382 ( .A(reg_A[120]), .B(n1767), .C(reg_A[104]), .D(n1768), .Y(
        n2073) );
  AOI22X1 U1383 ( .A(reg_A[56]), .B(n1766), .C(reg_A[16]), .D(n2049), .Y(n2072) );
  NAND2X1 U1384 ( .A(n2074), .B(n2075), .Y(U69_U7_Z_6) );
  AOI22X1 U1385 ( .A(reg_A[121]), .B(n1767), .C(reg_A[105]), .D(n2017), .Y(
        n2075) );
  AOI22X1 U1386 ( .A(reg_A[57]), .B(n1766), .C(reg_A[17]), .D(n2049), .Y(n2074) );
  NAND2X1 U1387 ( .A(n2076), .B(n2077), .Y(U69_U7_Z_5) );
  AOI22X1 U1388 ( .A(reg_A[122]), .B(n1767), .C(reg_A[106]), .D(n1768), .Y(
        n2077) );
  AOI22X1 U1389 ( .A(reg_A[58]), .B(n1766), .C(reg_A[18]), .D(n2049), .Y(n2076) );
  NAND2X1 U1390 ( .A(n2078), .B(n2079), .Y(U69_U7_Z_4) );
  AOI22X1 U1391 ( .A(reg_A[123]), .B(n1767), .C(reg_A[107]), .D(n1768), .Y(
        n2079) );
  AOI22X1 U1392 ( .A(reg_A[59]), .B(n1766), .C(reg_A[19]), .D(n1769), .Y(n2078) );
  NAND2X1 U1393 ( .A(n2080), .B(n2081), .Y(U69_U7_Z_3) );
  AOI22X1 U1394 ( .A(reg_A[124]), .B(n1767), .C(reg_A[108]), .D(n1768), .Y(
        n2081) );
  AOI22X1 U1395 ( .A(reg_A[60]), .B(n1766), .C(reg_A[20]), .D(n2049), .Y(n2080) );
  NAND2X1 U1396 ( .A(n2082), .B(n2083), .Y(U69_U7_Z_2) );
  AOI22X1 U1397 ( .A(reg_A[125]), .B(n1767), .C(reg_A[109]), .D(n1768), .Y(
        n2083) );
  AOI22X1 U1398 ( .A(reg_A[61]), .B(n1766), .C(reg_A[21]), .D(n2049), .Y(n2082) );
  INVX1 U1399 ( .A(n2084), .Y(U69_U7_Z_15) );
  AOI22X1 U1400 ( .A(n1768), .B(reg_A[96]), .C(n1767), .D(reg_A[112]), .Y(
        n2084) );
  INVX1 U1401 ( .A(n2085), .Y(U69_U7_Z_14) );
  AOI22X1 U1402 ( .A(n1768), .B(reg_A[97]), .C(n1767), .D(reg_A[113]), .Y(
        n2085) );
  INVX1 U1403 ( .A(n2086), .Y(U69_U7_Z_13) );
  AOI22X1 U1404 ( .A(n1768), .B(reg_A[98]), .C(n2018), .D(reg_A[114]), .Y(
        n2086) );
  INVX1 U1405 ( .A(n2087), .Y(U69_U7_Z_12) );
  AOI22X1 U1406 ( .A(n1768), .B(reg_A[99]), .C(n2018), .D(reg_A[115]), .Y(
        n2087) );
  INVX1 U1407 ( .A(n2088), .Y(U69_U7_Z_11) );
  AOI22X1 U1408 ( .A(n1768), .B(reg_A[100]), .C(n1767), .D(reg_A[116]), .Y(
        n2088) );
  INVX1 U1409 ( .A(n2089), .Y(U69_U7_Z_10) );
  AOI22X1 U1410 ( .A(n1768), .B(reg_A[101]), .C(n1767), .D(reg_A[117]), .Y(
        n2089) );
  NAND2X1 U1411 ( .A(n2090), .B(n2091), .Y(U69_U7_Z_1) );
  AOI22X1 U1412 ( .A(reg_A[126]), .B(n1767), .C(reg_A[110]), .D(n1768), .Y(
        n2091) );
  AOI22X1 U1413 ( .A(reg_A[62]), .B(n1766), .C(n1769), .D(reg_A[22]), .Y(n2090) );
  NAND2X1 U1414 ( .A(n2092), .B(n2093), .Y(U69_U7_Z_0) );
  AOI22X1 U1415 ( .A(reg_A[127]), .B(n1767), .C(reg_A[111]), .D(n1768), .Y(
        n2093) );
  AOI22X1 U1416 ( .A(reg_A[63]), .B(n1766), .C(n1769), .D(reg_A[23]), .Y(n2092) );
  INVX1 U1417 ( .A(n2094), .Y(U69_U6_Z_7) );
  MUX2X1 U1418 ( .B(reg_B[120]), .A(reg_B[64]), .S(n2011), .Y(n2094) );
  INVX1 U1419 ( .A(n2095), .Y(U69_U6_Z_6) );
  MUX2X1 U1420 ( .B(reg_B[121]), .A(reg_B[65]), .S(n2011), .Y(n2095) );
  INVX1 U1421 ( .A(n2096), .Y(U69_U6_Z_5) );
  MUX2X1 U1422 ( .B(reg_B[122]), .A(reg_B[66]), .S(n2011), .Y(n2096) );
  INVX1 U1423 ( .A(n2097), .Y(U69_U6_Z_4) );
  MUX2X1 U1424 ( .B(reg_B[123]), .A(reg_B[67]), .S(n2011), .Y(n2097) );
  INVX1 U1425 ( .A(n2098), .Y(U69_U6_Z_3) );
  MUX2X1 U1426 ( .B(reg_B[124]), .A(reg_B[68]), .S(n2011), .Y(n2098) );
  INVX1 U1427 ( .A(n2099), .Y(U69_U6_Z_2) );
  MUX2X1 U1428 ( .B(reg_B[125]), .A(reg_B[69]), .S(n2011), .Y(n2099) );
  INVX1 U1429 ( .A(n2100), .Y(U69_U6_Z_1) );
  MUX2X1 U1430 ( .B(reg_B[126]), .A(reg_B[70]), .S(n2011), .Y(n2100) );
  INVX1 U1431 ( .A(n2101), .Y(U69_U6_Z_0) );
  MUX2X1 U1432 ( .B(reg_B[127]), .A(reg_B[71]), .S(n2011), .Y(n2101) );
  INVX1 U1433 ( .A(n2102), .Y(U69_U5_Z_7) );
  MUX2X1 U1434 ( .B(reg_A[120]), .A(reg_A[64]), .S(n2011), .Y(n2102) );
  INVX1 U1435 ( .A(n2103), .Y(U69_U5_Z_6) );
  MUX2X1 U1436 ( .B(reg_A[121]), .A(reg_A[65]), .S(n2011), .Y(n2103) );
  INVX1 U1437 ( .A(n2104), .Y(U69_U5_Z_5) );
  MUX2X1 U1438 ( .B(reg_A[122]), .A(reg_A[66]), .S(n2011), .Y(n2104) );
  INVX1 U1439 ( .A(n2105), .Y(U69_U5_Z_4) );
  MUX2X1 U1440 ( .B(reg_A[123]), .A(reg_A[67]), .S(n2011), .Y(n2105) );
  INVX1 U1441 ( .A(n2106), .Y(U69_U5_Z_3) );
  MUX2X1 U1442 ( .B(reg_A[124]), .A(reg_A[68]), .S(n2011), .Y(n2106) );
  INVX1 U1443 ( .A(n2107), .Y(U69_U5_Z_2) );
  MUX2X1 U1444 ( .B(reg_A[125]), .A(reg_A[69]), .S(n2011), .Y(n2107) );
  INVX1 U1445 ( .A(n2108), .Y(U69_U5_Z_1) );
  MUX2X1 U1446 ( .B(reg_A[126]), .A(reg_A[70]), .S(n2011), .Y(n2108) );
  INVX1 U1447 ( .A(n2109), .Y(U69_U5_Z_0) );
  MUX2X1 U1448 ( .B(reg_A[127]), .A(reg_A[71]), .S(n2011), .Y(n2109) );
  INVX1 U1449 ( .A(n2110), .Y(U69_U4_Z_9) );
  AOI22X1 U1450 ( .A(n1768), .B(reg_B[6]), .C(n1767), .D(reg_B[54]), .Y(n2110)
         );
  INVX1 U1451 ( .A(n2111), .Y(U69_U4_Z_8) );
  AOI22X1 U1452 ( .A(n1768), .B(reg_B[7]), .C(n1767), .D(reg_B[55]), .Y(n2111)
         );
  NAND2X1 U1453 ( .A(n2112), .B(n2113), .Y(U69_U4_Z_7) );
  AOI22X1 U1454 ( .A(reg_B[56]), .B(n1767), .C(reg_B[8]), .D(n2017), .Y(n2113)
         );
  AOI22X1 U1455 ( .A(reg_B[72]), .B(n1766), .C(reg_B[48]), .D(n2049), .Y(n2112) );
  NAND2X1 U1456 ( .A(n2114), .B(n2115), .Y(U69_U4_Z_6) );
  AOI22X1 U1457 ( .A(reg_B[57]), .B(n1767), .C(reg_B[9]), .D(n2017), .Y(n2115)
         );
  AOI22X1 U1458 ( .A(reg_B[73]), .B(n1766), .C(reg_B[49]), .D(n2049), .Y(n2114) );
  NAND2X1 U1459 ( .A(n2116), .B(n2117), .Y(U69_U4_Z_5) );
  AOI22X1 U1460 ( .A(reg_B[58]), .B(n1767), .C(reg_B[10]), .D(n2017), .Y(n2117) );
  AOI22X1 U1461 ( .A(reg_B[74]), .B(n1766), .C(reg_B[50]), .D(n2049), .Y(n2116) );
  NAND2X1 U1462 ( .A(n2118), .B(n2119), .Y(U69_U4_Z_4) );
  AOI22X1 U1463 ( .A(reg_B[59]), .B(n1767), .C(reg_B[11]), .D(n1768), .Y(n2119) );
  AOI22X1 U1464 ( .A(reg_B[75]), .B(n1766), .C(reg_B[51]), .D(n2049), .Y(n2118) );
  NAND2X1 U1465 ( .A(n2120), .B(n2121), .Y(U69_U4_Z_3) );
  AOI22X1 U1466 ( .A(reg_B[60]), .B(n1767), .C(reg_B[12]), .D(n1768), .Y(n2121) );
  AOI22X1 U1467 ( .A(reg_B[76]), .B(n1766), .C(reg_B[52]), .D(n2049), .Y(n2120) );
  NAND2X1 U1468 ( .A(n2122), .B(n2123), .Y(U69_U4_Z_2) );
  AOI22X1 U1469 ( .A(reg_B[61]), .B(n1767), .C(reg_B[13]), .D(n2017), .Y(n2123) );
  AOI22X1 U1470 ( .A(reg_B[77]), .B(n1766), .C(reg_B[53]), .D(n2049), .Y(n2122) );
  INVX1 U1471 ( .A(n2124), .Y(U69_U4_Z_15) );
  AOI22X1 U1472 ( .A(n1768), .B(reg_B[0]), .C(n1767), .D(reg_B[48]), .Y(n2124)
         );
  INVX1 U1473 ( .A(n2125), .Y(U69_U4_Z_14) );
  AOI22X1 U1474 ( .A(n1768), .B(reg_B[1]), .C(n1767), .D(reg_B[49]), .Y(n2125)
         );
  INVX1 U1475 ( .A(n2126), .Y(U69_U4_Z_13) );
  AOI22X1 U1476 ( .A(n1768), .B(reg_B[2]), .C(n1767), .D(reg_B[50]), .Y(n2126)
         );
  INVX1 U1477 ( .A(n2127), .Y(U69_U4_Z_12) );
  AOI22X1 U1478 ( .A(n1768), .B(reg_B[3]), .C(n2018), .D(reg_B[51]), .Y(n2127)
         );
  INVX1 U1479 ( .A(n2128), .Y(U69_U4_Z_11) );
  AOI22X1 U1480 ( .A(n1768), .B(reg_B[4]), .C(n1767), .D(reg_B[52]), .Y(n2128)
         );
  INVX1 U1481 ( .A(n2129), .Y(U69_U4_Z_10) );
  AOI22X1 U1482 ( .A(n1768), .B(reg_B[5]), .C(n1767), .D(reg_B[53]), .Y(n2129)
         );
  NAND2X1 U1483 ( .A(n2130), .B(n2131), .Y(U69_U4_Z_1) );
  AOI22X1 U1484 ( .A(reg_B[62]), .B(n1767), .C(reg_B[14]), .D(n1768), .Y(n2131) );
  AOI22X1 U1485 ( .A(reg_B[78]), .B(n1766), .C(reg_B[54]), .D(n1769), .Y(n2130) );
  NAND2X1 U1486 ( .A(n2132), .B(n2133), .Y(U69_U4_Z_0) );
  AOI22X1 U1487 ( .A(reg_B[63]), .B(n1767), .C(reg_B[15]), .D(n1768), .Y(n2133) );
  AOI22X1 U1488 ( .A(reg_B[79]), .B(n1766), .C(reg_B[55]), .D(n2049), .Y(n2132) );
  INVX1 U1489 ( .A(n2134), .Y(U69_U3_Z_9) );
  AOI22X1 U1490 ( .A(n1768), .B(reg_A[6]), .C(n1767), .D(reg_A[54]), .Y(n2134)
         );
  INVX1 U1491 ( .A(n2135), .Y(U69_U3_Z_8) );
  AOI22X1 U1492 ( .A(n1768), .B(reg_A[7]), .C(n2018), .D(reg_A[55]), .Y(n2135)
         );
  NAND2X1 U1493 ( .A(n2136), .B(n2137), .Y(U69_U3_Z_7) );
  AOI22X1 U1494 ( .A(reg_A[56]), .B(n1767), .C(reg_A[8]), .D(n2017), .Y(n2137)
         );
  AOI22X1 U1495 ( .A(n1766), .B(reg_A[72]), .C(reg_A[48]), .D(n1769), .Y(n2136) );
  NAND2X1 U1496 ( .A(n2138), .B(n2139), .Y(U69_U3_Z_6) );
  AOI22X1 U1497 ( .A(reg_A[57]), .B(n1767), .C(reg_A[9]), .D(n2017), .Y(n2139)
         );
  AOI22X1 U1498 ( .A(n1766), .B(reg_A[73]), .C(reg_A[49]), .D(n1769), .Y(n2138) );
  NAND2X1 U1499 ( .A(n2140), .B(n2141), .Y(U69_U3_Z_5) );
  AOI22X1 U1500 ( .A(reg_A[58]), .B(n1767), .C(reg_A[10]), .D(n1768), .Y(n2141) );
  AOI22X1 U1501 ( .A(n1766), .B(reg_A[74]), .C(reg_A[50]), .D(n1769), .Y(n2140) );
  NAND2X1 U1502 ( .A(n2142), .B(n2143), .Y(U69_U3_Z_4) );
  AOI22X1 U1503 ( .A(reg_A[59]), .B(n1767), .C(reg_A[11]), .D(n1768), .Y(n2143) );
  AOI22X1 U1504 ( .A(n1766), .B(reg_A[75]), .C(reg_A[51]), .D(n1769), .Y(n2142) );
  NAND2X1 U1505 ( .A(n2144), .B(n2145), .Y(U69_U3_Z_3) );
  AOI22X1 U1506 ( .A(reg_A[60]), .B(n1767), .C(reg_A[12]), .D(n1768), .Y(n2145) );
  AOI22X1 U1507 ( .A(n1766), .B(reg_A[76]), .C(reg_A[52]), .D(n1769), .Y(n2144) );
  NAND2X1 U1508 ( .A(n2146), .B(n2147), .Y(U69_U3_Z_2) );
  AOI22X1 U1509 ( .A(reg_A[61]), .B(n1767), .C(reg_A[13]), .D(n1768), .Y(n2147) );
  AOI22X1 U1510 ( .A(n1766), .B(reg_A[77]), .C(reg_A[53]), .D(n1769), .Y(n2146) );
  INVX1 U1511 ( .A(n2148), .Y(U69_U3_Z_15) );
  AOI22X1 U1512 ( .A(n1768), .B(reg_A[0]), .C(n1767), .D(reg_A[48]), .Y(n2148)
         );
  INVX1 U1513 ( .A(n2149), .Y(U69_U3_Z_14) );
  AOI22X1 U1514 ( .A(n1768), .B(reg_A[1]), .C(n2018), .D(reg_A[49]), .Y(n2149)
         );
  INVX1 U1515 ( .A(n2150), .Y(U69_U3_Z_13) );
  AOI22X1 U1516 ( .A(n1768), .B(reg_A[2]), .C(n2018), .D(reg_A[50]), .Y(n2150)
         );
  INVX1 U1517 ( .A(n2151), .Y(U69_U3_Z_12) );
  AOI22X1 U1518 ( .A(n1768), .B(reg_A[3]), .C(n1767), .D(reg_A[51]), .Y(n2151)
         );
  INVX1 U1519 ( .A(n2152), .Y(U69_U3_Z_11) );
  AOI22X1 U1520 ( .A(n1768), .B(reg_A[4]), .C(n2018), .D(reg_A[52]), .Y(n2152)
         );
  INVX1 U1521 ( .A(n2153), .Y(U69_U3_Z_10) );
  AOI22X1 U1522 ( .A(n1768), .B(reg_A[5]), .C(n1767), .D(reg_A[53]), .Y(n2153)
         );
  NAND2X1 U1523 ( .A(n2154), .B(n2155), .Y(U69_U3_Z_1) );
  AOI22X1 U1524 ( .A(reg_A[62]), .B(n1767), .C(reg_A[14]), .D(n1768), .Y(n2155) );
  AOI22X1 U1525 ( .A(n1766), .B(reg_A[78]), .C(reg_A[54]), .D(n1769), .Y(n2154) );
  NAND2X1 U1526 ( .A(n2156), .B(n2157), .Y(U69_U3_Z_0) );
  AOI22X1 U1527 ( .A(reg_A[63]), .B(n1767), .C(reg_A[15]), .D(n2017), .Y(n2157) );
  AOI22X1 U1528 ( .A(n1766), .B(reg_A[79]), .C(reg_A[55]), .D(n1769), .Y(n2156) );
  OAI22X1 U1529 ( .A(n2158), .B(n2159), .C(n2160), .D(n2161), .Y(U69_U2_Z_9)
         );
  INVX1 U1530 ( .A(reg_B[86]), .Y(n2161) );
  OAI22X1 U1531 ( .A(n2158), .B(n2162), .C(n2160), .D(n2163), .Y(U69_U2_Z_8)
         );
  INVX1 U1532 ( .A(reg_B[87]), .Y(n2163) );
  NAND2X1 U1533 ( .A(n2164), .B(n2165), .Y(U69_U2_Z_7) );
  AOI22X1 U1534 ( .A(reg_B[88]), .B(n1767), .C(reg_B[40]), .D(n2017), .Y(n2165) );
  AOI22X1 U1535 ( .A(reg_B[8]), .B(n1766), .C(reg_B[112]), .D(n1769), .Y(n2164) );
  NAND2X1 U1536 ( .A(n2166), .B(n2167), .Y(U69_U2_Z_6) );
  AOI22X1 U1537 ( .A(reg_B[89]), .B(n1767), .C(reg_B[41]), .D(n1768), .Y(n2167) );
  AOI22X1 U1538 ( .A(reg_B[9]), .B(n1766), .C(reg_B[113]), .D(n1769), .Y(n2166) );
  NAND2X1 U1539 ( .A(n2168), .B(n2169), .Y(U69_U2_Z_5) );
  AOI22X1 U1540 ( .A(reg_B[90]), .B(n1767), .C(reg_B[42]), .D(n1768), .Y(n2169) );
  AOI22X1 U1541 ( .A(reg_B[10]), .B(n1766), .C(reg_B[114]), .D(n1769), .Y(
        n2168) );
  NAND2X1 U1542 ( .A(n2170), .B(n2171), .Y(U69_U2_Z_4) );
  AOI22X1 U1543 ( .A(reg_B[91]), .B(n1767), .C(reg_B[43]), .D(n1768), .Y(n2171) );
  AOI22X1 U1544 ( .A(reg_B[11]), .B(n1766), .C(reg_B[115]), .D(n1769), .Y(
        n2170) );
  NAND2X1 U1545 ( .A(n2172), .B(n2173), .Y(U69_U2_Z_3) );
  AOI22X1 U1546 ( .A(reg_B[92]), .B(n1767), .C(reg_B[44]), .D(n2017), .Y(n2173) );
  AOI22X1 U1547 ( .A(reg_B[12]), .B(n1766), .C(reg_B[116]), .D(n1769), .Y(
        n2172) );
  NAND2X1 U1548 ( .A(n2174), .B(n2175), .Y(U69_U2_Z_2) );
  AOI22X1 U1549 ( .A(reg_B[93]), .B(n1767), .C(reg_B[45]), .D(n1768), .Y(n2175) );
  AOI22X1 U1550 ( .A(reg_B[13]), .B(n1766), .C(reg_B[117]), .D(n1769), .Y(
        n2174) );
  OAI22X1 U1551 ( .A(n2158), .B(n2176), .C(n2160), .D(n2177), .Y(U69_U2_Z_15)
         );
  INVX1 U1552 ( .A(reg_B[80]), .Y(n2177) );
  OAI22X1 U1553 ( .A(n2158), .B(n2178), .C(n2160), .D(n2179), .Y(U69_U2_Z_14)
         );
  INVX1 U1554 ( .A(reg_B[81]), .Y(n2179) );
  OAI22X1 U1555 ( .A(n2158), .B(n2180), .C(n2160), .D(n2181), .Y(U69_U2_Z_13)
         );
  INVX1 U1556 ( .A(reg_B[82]), .Y(n2181) );
  OAI22X1 U1557 ( .A(n2158), .B(n2182), .C(n2160), .D(n2183), .Y(U69_U2_Z_12)
         );
  INVX1 U1558 ( .A(reg_B[83]), .Y(n2183) );
  OAI22X1 U1559 ( .A(n2158), .B(n2184), .C(n2160), .D(n2185), .Y(U69_U2_Z_11)
         );
  INVX1 U1560 ( .A(reg_B[84]), .Y(n2185) );
  OAI22X1 U1561 ( .A(n2158), .B(n2186), .C(n2160), .D(n2187), .Y(U69_U2_Z_10)
         );
  INVX1 U1562 ( .A(reg_B[85]), .Y(n2187) );
  INVX1 U1563 ( .A(n2018), .Y(n2160) );
  INVX1 U1564 ( .A(n2017), .Y(n2158) );
  NAND2X1 U1565 ( .A(n2188), .B(n2189), .Y(U69_U2_Z_1) );
  AOI22X1 U1566 ( .A(reg_B[94]), .B(n1767), .C(reg_B[46]), .D(n1768), .Y(n2189) );
  AOI22X1 U1567 ( .A(reg_B[14]), .B(n1766), .C(reg_B[118]), .D(n1769), .Y(
        n2188) );
  NAND2X1 U1568 ( .A(n2190), .B(n2191), .Y(U69_U2_Z_0) );
  AOI22X1 U1569 ( .A(reg_B[95]), .B(n1767), .C(reg_B[47]), .D(n1768), .Y(n2191) );
  AOI22X1 U1570 ( .A(reg_B[15]), .B(n1766), .C(reg_B[119]), .D(n1769), .Y(
        n2190) );
  INVX1 U1571 ( .A(n2192), .Y(U69_U16_Z_7) );
  MUX2X1 U1572 ( .B(reg_B[104]), .A(reg_B[96]), .S(n2011), .Y(n2192) );
  INVX1 U1573 ( .A(n2193), .Y(U69_U16_Z_6) );
  MUX2X1 U1574 ( .B(reg_B[105]), .A(reg_B[97]), .S(n2011), .Y(n2193) );
  INVX1 U1575 ( .A(n2194), .Y(U69_U16_Z_5) );
  MUX2X1 U1576 ( .B(reg_B[106]), .A(reg_B[98]), .S(n2011), .Y(n2194) );
  INVX1 U1577 ( .A(n2195), .Y(U69_U16_Z_4) );
  MUX2X1 U1578 ( .B(reg_B[107]), .A(reg_B[99]), .S(n2011), .Y(n2195) );
  INVX1 U1579 ( .A(n2196), .Y(U69_U16_Z_3) );
  MUX2X1 U1580 ( .B(reg_B[108]), .A(reg_B[100]), .S(n2011), .Y(n2196) );
  INVX1 U1581 ( .A(n2197), .Y(U69_U16_Z_2) );
  MUX2X1 U1582 ( .B(reg_B[109]), .A(reg_B[101]), .S(n2011), .Y(n2197) );
  INVX1 U1583 ( .A(n2198), .Y(U69_U16_Z_1) );
  MUX2X1 U1584 ( .B(reg_B[110]), .A(reg_B[102]), .S(n2011), .Y(n2198) );
  INVX1 U1585 ( .A(n2199), .Y(U69_U16_Z_0) );
  MUX2X1 U1586 ( .B(reg_B[111]), .A(reg_B[103]), .S(n2011), .Y(n2199) );
  INVX1 U1587 ( .A(n2200), .Y(U69_U15_Z_7) );
  MUX2X1 U1588 ( .B(reg_A[104]), .A(reg_A[96]), .S(n2011), .Y(n2200) );
  INVX1 U1589 ( .A(n2201), .Y(U69_U15_Z_6) );
  MUX2X1 U1590 ( .B(reg_A[105]), .A(reg_A[97]), .S(n2011), .Y(n2201) );
  INVX1 U1591 ( .A(n2202), .Y(U69_U15_Z_5) );
  MUX2X1 U1592 ( .B(reg_A[106]), .A(reg_A[98]), .S(n2011), .Y(n2202) );
  INVX1 U1593 ( .A(n2203), .Y(U69_U15_Z_4) );
  MUX2X1 U1594 ( .B(reg_A[107]), .A(reg_A[99]), .S(n2011), .Y(n2203) );
  INVX1 U1595 ( .A(n2204), .Y(U69_U15_Z_3) );
  MUX2X1 U1596 ( .B(reg_A[108]), .A(reg_A[100]), .S(n2011), .Y(n2204) );
  INVX1 U1597 ( .A(n2205), .Y(U69_U15_Z_2) );
  MUX2X1 U1598 ( .B(reg_A[109]), .A(reg_A[101]), .S(n2011), .Y(n2205) );
  INVX1 U1599 ( .A(n2206), .Y(U69_U15_Z_1) );
  MUX2X1 U1600 ( .B(reg_A[110]), .A(reg_A[102]), .S(n2011), .Y(n2206) );
  INVX1 U1601 ( .A(n2207), .Y(U69_U15_Z_0) );
  MUX2X1 U1602 ( .B(reg_A[111]), .A(reg_A[103]), .S(n2011), .Y(n2207) );
  INVX1 U1603 ( .A(n2208), .Y(U69_U14_Z_7) );
  MUX2X1 U1604 ( .B(reg_B[88]), .A(reg_B[0]), .S(n2011), .Y(n2208) );
  INVX1 U1605 ( .A(n2209), .Y(U69_U14_Z_6) );
  MUX2X1 U1606 ( .B(reg_B[89]), .A(reg_B[1]), .S(n2011), .Y(n2209) );
  INVX1 U1607 ( .A(n2210), .Y(U69_U14_Z_5) );
  MUX2X1 U1608 ( .B(reg_B[90]), .A(reg_B[2]), .S(n2011), .Y(n2210) );
  INVX1 U1609 ( .A(n2211), .Y(U69_U14_Z_4) );
  MUX2X1 U1610 ( .B(reg_B[91]), .A(reg_B[3]), .S(n2011), .Y(n2211) );
  INVX1 U1611 ( .A(n2212), .Y(U69_U14_Z_3) );
  MUX2X1 U1612 ( .B(reg_B[92]), .A(reg_B[4]), .S(n2011), .Y(n2212) );
  INVX1 U1613 ( .A(n2213), .Y(U69_U14_Z_2) );
  MUX2X1 U1614 ( .B(reg_B[93]), .A(reg_B[5]), .S(n2011), .Y(n2213) );
  INVX1 U1615 ( .A(n2214), .Y(U69_U14_Z_1) );
  MUX2X1 U1616 ( .B(reg_B[94]), .A(reg_B[6]), .S(n2011), .Y(n2214) );
  INVX1 U1617 ( .A(n2215), .Y(U69_U14_Z_0) );
  MUX2X1 U1618 ( .B(reg_B[95]), .A(reg_B[7]), .S(n2011), .Y(n2215) );
  INVX1 U1619 ( .A(n2216), .Y(U69_U13_Z_7) );
  MUX2X1 U1620 ( .B(reg_A[88]), .A(reg_A[0]), .S(n2011), .Y(n2216) );
  INVX1 U1621 ( .A(n2217), .Y(U69_U13_Z_6) );
  MUX2X1 U1622 ( .B(reg_A[89]), .A(reg_A[1]), .S(n2011), .Y(n2217) );
  INVX1 U1623 ( .A(n2218), .Y(U69_U13_Z_5) );
  MUX2X1 U1624 ( .B(reg_A[90]), .A(reg_A[2]), .S(n2011), .Y(n2218) );
  INVX1 U1625 ( .A(n2219), .Y(U69_U13_Z_4) );
  MUX2X1 U1626 ( .B(reg_A[91]), .A(reg_A[3]), .S(n2011), .Y(n2219) );
  INVX1 U1627 ( .A(n2220), .Y(U69_U13_Z_3) );
  MUX2X1 U1628 ( .B(reg_A[92]), .A(reg_A[4]), .S(n2011), .Y(n2220) );
  INVX1 U1629 ( .A(n2221), .Y(U69_U13_Z_2) );
  MUX2X1 U1630 ( .B(reg_A[93]), .A(reg_A[5]), .S(n2011), .Y(n2221) );
  INVX1 U1631 ( .A(n2222), .Y(U69_U13_Z_1) );
  MUX2X1 U1632 ( .B(reg_A[94]), .A(reg_A[6]), .S(n2011), .Y(n2222) );
  INVX1 U1633 ( .A(n2223), .Y(U69_U13_Z_0) );
  MUX2X1 U1634 ( .B(reg_A[95]), .A(reg_A[7]), .S(n2011), .Y(n2223) );
  INVX1 U1635 ( .A(n2224), .Y(U69_U12_Z_7) );
  MUX2X1 U1636 ( .B(reg_B[40]), .A(reg_B[80]), .S(n2011), .Y(n2224) );
  INVX1 U1637 ( .A(n2225), .Y(U69_U12_Z_6) );
  MUX2X1 U1638 ( .B(reg_B[41]), .A(reg_B[81]), .S(n2011), .Y(n2225) );
  INVX1 U1639 ( .A(n2226), .Y(U69_U12_Z_5) );
  MUX2X1 U1640 ( .B(reg_B[42]), .A(reg_B[82]), .S(n2011), .Y(n2226) );
  INVX1 U1641 ( .A(n2227), .Y(U69_U12_Z_4) );
  MUX2X1 U1642 ( .B(reg_B[43]), .A(reg_B[83]), .S(n2011), .Y(n2227) );
  INVX1 U1643 ( .A(n2228), .Y(U69_U12_Z_3) );
  MUX2X1 U1644 ( .B(reg_B[44]), .A(reg_B[84]), .S(n2011), .Y(n2228) );
  INVX1 U1645 ( .A(n2229), .Y(U69_U12_Z_2) );
  MUX2X1 U1646 ( .B(reg_B[45]), .A(reg_B[85]), .S(n2011), .Y(n2229) );
  INVX1 U1647 ( .A(n2230), .Y(U69_U12_Z_1) );
  MUX2X1 U1648 ( .B(reg_B[46]), .A(reg_B[86]), .S(n2011), .Y(n2230) );
  INVX1 U1649 ( .A(n2231), .Y(U69_U12_Z_0) );
  MUX2X1 U1650 ( .B(reg_B[47]), .A(reg_B[87]), .S(n2011), .Y(n2231) );
  INVX1 U1651 ( .A(n2232), .Y(U69_U11_Z_7) );
  MUX2X1 U1652 ( .B(reg_A[40]), .A(reg_A[80]), .S(n2011), .Y(n2232) );
  INVX1 U1653 ( .A(n2233), .Y(U69_U11_Z_6) );
  MUX2X1 U1654 ( .B(reg_A[41]), .A(reg_A[81]), .S(n2011), .Y(n2233) );
  INVX1 U1655 ( .A(n2234), .Y(U69_U11_Z_5) );
  MUX2X1 U1656 ( .B(reg_A[42]), .A(reg_A[82]), .S(n2011), .Y(n2234) );
  INVX1 U1657 ( .A(n2235), .Y(U69_U11_Z_4) );
  MUX2X1 U1658 ( .B(reg_A[43]), .A(reg_A[83]), .S(n2011), .Y(n2235) );
  INVX1 U1659 ( .A(n2236), .Y(U69_U11_Z_3) );
  MUX2X1 U1660 ( .B(reg_A[44]), .A(reg_A[84]), .S(n2011), .Y(n2236) );
  INVX1 U1661 ( .A(n2237), .Y(U69_U11_Z_2) );
  MUX2X1 U1662 ( .B(reg_A[45]), .A(reg_A[85]), .S(n2011), .Y(n2237) );
  INVX1 U1663 ( .A(n2238), .Y(U69_U11_Z_1) );
  MUX2X1 U1664 ( .B(reg_A[46]), .A(reg_A[86]), .S(n2011), .Y(n2238) );
  INVX1 U1665 ( .A(n2239), .Y(U69_U11_Z_0) );
  MUX2X1 U1666 ( .B(reg_A[47]), .A(reg_A[87]), .S(n2011), .Y(n2239) );
  INVX1 U1667 ( .A(n2240), .Y(U69_U10_Z_9) );
  AOI22X1 U1668 ( .A(n1768), .B(reg_B[70]), .C(n2018), .D(reg_B[22]), .Y(n2240) );
  INVX1 U1669 ( .A(n2241), .Y(U69_U10_Z_8) );
  AOI22X1 U1670 ( .A(n1768), .B(reg_B[71]), .C(n2018), .D(reg_B[23]), .Y(n2241) );
  OAI21X1 U1671 ( .A(n2020), .B(n2176), .C(n2242), .Y(U69_U10_Z_7) );
  AOI22X1 U1672 ( .A(reg_B[24]), .B(n2023), .C(reg_B[72]), .D(n1768), .Y(n2242) );
  INVX1 U1673 ( .A(reg_B[32]), .Y(n2176) );
  OAI21X1 U1674 ( .A(n2020), .B(n2178), .C(n2243), .Y(U69_U10_Z_6) );
  AOI22X1 U1675 ( .A(reg_B[25]), .B(n2023), .C(reg_B[73]), .D(n2017), .Y(n2243) );
  INVX1 U1676 ( .A(reg_B[33]), .Y(n2178) );
  OAI21X1 U1677 ( .A(n2020), .B(n2180), .C(n2244), .Y(U69_U10_Z_5) );
  AOI22X1 U1678 ( .A(reg_B[26]), .B(n2023), .C(reg_B[74]), .D(n2017), .Y(n2244) );
  INVX1 U1679 ( .A(reg_B[34]), .Y(n2180) );
  OAI21X1 U1680 ( .A(n2020), .B(n2182), .C(n2245), .Y(U69_U10_Z_4) );
  AOI22X1 U1681 ( .A(reg_B[27]), .B(n2023), .C(reg_B[75]), .D(n2017), .Y(n2245) );
  INVX1 U1682 ( .A(reg_B[35]), .Y(n2182) );
  OAI21X1 U1683 ( .A(n2020), .B(n2184), .C(n2246), .Y(U69_U10_Z_3) );
  AOI22X1 U1684 ( .A(reg_B[28]), .B(n2023), .C(reg_B[76]), .D(n1768), .Y(n2246) );
  INVX1 U1685 ( .A(reg_B[36]), .Y(n2184) );
  OAI21X1 U1686 ( .A(n2020), .B(n2186), .C(n2247), .Y(U69_U10_Z_2) );
  AOI22X1 U1687 ( .A(reg_B[29]), .B(n2023), .C(reg_B[77]), .D(n2017), .Y(n2247) );
  INVX1 U1688 ( .A(reg_B[37]), .Y(n2186) );
  INVX1 U1689 ( .A(n2248), .Y(U69_U10_Z_15) );
  AOI22X1 U1690 ( .A(n1768), .B(reg_B[64]), .C(n1767), .D(reg_B[16]), .Y(n2248) );
  INVX1 U1691 ( .A(n2249), .Y(U69_U10_Z_14) );
  AOI22X1 U1692 ( .A(n1768), .B(reg_B[65]), .C(n1767), .D(reg_B[17]), .Y(n2249) );
  INVX1 U1693 ( .A(n2250), .Y(U69_U10_Z_13) );
  AOI22X1 U1694 ( .A(n1768), .B(reg_B[66]), .C(n1767), .D(reg_B[18]), .Y(n2250) );
  INVX1 U1695 ( .A(n2251), .Y(U69_U10_Z_12) );
  AOI22X1 U1696 ( .A(n1768), .B(reg_B[67]), .C(n1767), .D(reg_B[19]), .Y(n2251) );
  INVX1 U1697 ( .A(n2252), .Y(U69_U10_Z_11) );
  AOI22X1 U1698 ( .A(n1768), .B(reg_B[68]), .C(n1767), .D(reg_B[20]), .Y(n2252) );
  INVX1 U1699 ( .A(n2253), .Y(U69_U10_Z_10) );
  AOI22X1 U1700 ( .A(n1768), .B(reg_B[69]), .C(n2018), .D(reg_B[21]), .Y(n2253) );
  OAI21X1 U1701 ( .A(n2020), .B(n2159), .C(n2254), .Y(U69_U10_Z_1) );
  AOI22X1 U1702 ( .A(reg_B[30]), .B(n2023), .C(reg_B[78]), .D(n2017), .Y(n2254) );
  INVX1 U1703 ( .A(reg_B[38]), .Y(n2159) );
  OAI21X1 U1704 ( .A(n2020), .B(n2162), .C(n2255), .Y(U69_U10_Z_0) );
  AOI22X1 U1705 ( .A(reg_B[31]), .B(n2023), .C(reg_B[79]), .D(n1768), .Y(n2255) );
  OR2X1 U1706 ( .A(n1766), .B(n1767), .Y(n2023) );
  INVX1 U1707 ( .A(reg_B[39]), .Y(n2162) );
  INVX1 U1708 ( .A(n2049), .Y(n2020) );
  INVX1 U1709 ( .A(n2256), .Y(U69_U1_Z_9) );
  AOI22X1 U1710 ( .A(n1768), .B(reg_A[38]), .C(n1767), .D(reg_A[86]), .Y(n2256) );
  INVX1 U1711 ( .A(n2257), .Y(U69_U1_Z_8) );
  AOI22X1 U1712 ( .A(n1768), .B(reg_A[39]), .C(n2018), .D(reg_A[87]), .Y(n2257) );
  NAND2X1 U1713 ( .A(n2258), .B(n2259), .Y(U69_U1_Z_7) );
  AOI22X1 U1714 ( .A(reg_A[88]), .B(n1767), .C(reg_A[40]), .D(n2017), .Y(n2259) );
  AOI22X1 U1715 ( .A(reg_A[8]), .B(n1766), .C(reg_A[112]), .D(n1769), .Y(n2258) );
  NAND2X1 U1716 ( .A(n2260), .B(n2261), .Y(U69_U1_Z_6) );
  AOI22X1 U1717 ( .A(reg_A[89]), .B(n1767), .C(reg_A[41]), .D(n1768), .Y(n2261) );
  AOI22X1 U1718 ( .A(reg_A[9]), .B(n1766), .C(reg_A[113]), .D(n1769), .Y(n2260) );
  NAND2X1 U1719 ( .A(n2262), .B(n2263), .Y(U69_U1_Z_5) );
  AOI22X1 U1720 ( .A(reg_A[90]), .B(n1767), .C(reg_A[42]), .D(n1768), .Y(n2263) );
  AOI22X1 U1721 ( .A(reg_A[10]), .B(n1766), .C(reg_A[114]), .D(n1769), .Y(
        n2262) );
  NAND2X1 U1722 ( .A(n2264), .B(n2265), .Y(U69_U1_Z_4) );
  AOI22X1 U1723 ( .A(reg_A[91]), .B(n1767), .C(reg_A[43]), .D(n2017), .Y(n2265) );
  AOI22X1 U1724 ( .A(reg_A[11]), .B(n1766), .C(reg_A[115]), .D(n1769), .Y(
        n2264) );
  NAND2X1 U1725 ( .A(n2266), .B(n2267), .Y(U69_U1_Z_3) );
  AOI22X1 U1726 ( .A(reg_A[92]), .B(n1767), .C(reg_A[44]), .D(n1768), .Y(n2267) );
  AOI22X1 U1727 ( .A(reg_A[12]), .B(n1766), .C(reg_A[116]), .D(n1769), .Y(
        n2266) );
  NAND2X1 U1728 ( .A(n2268), .B(n2269), .Y(U69_U1_Z_2) );
  AOI22X1 U1729 ( .A(reg_A[93]), .B(n1767), .C(reg_A[45]), .D(n1768), .Y(n2269) );
  AOI22X1 U1730 ( .A(reg_A[13]), .B(n1766), .C(reg_A[117]), .D(n1769), .Y(
        n2268) );
  INVX1 U1731 ( .A(n2270), .Y(U69_U1_Z_15) );
  AOI22X1 U1732 ( .A(n1768), .B(reg_A[32]), .C(n1767), .D(reg_A[80]), .Y(n2270) );
  INVX1 U1733 ( .A(n2271), .Y(U69_U1_Z_14) );
  AOI22X1 U1734 ( .A(n1768), .B(reg_A[33]), .C(n1767), .D(reg_A[81]), .Y(n2271) );
  INVX1 U1735 ( .A(n2272), .Y(U69_U1_Z_13) );
  AOI22X1 U1736 ( .A(n1768), .B(reg_A[34]), .C(n2018), .D(reg_A[82]), .Y(n2272) );
  INVX1 U1737 ( .A(n2273), .Y(U69_U1_Z_12) );
  AOI22X1 U1738 ( .A(n1768), .B(reg_A[35]), .C(n1767), .D(reg_A[83]), .Y(n2273) );
  INVX1 U1739 ( .A(n2274), .Y(U69_U1_Z_11) );
  AOI22X1 U1740 ( .A(n1768), .B(reg_A[36]), .C(n1767), .D(reg_A[84]), .Y(n2274) );
  INVX1 U1741 ( .A(n2275), .Y(U69_U1_Z_10) );
  AOI22X1 U1742 ( .A(n1768), .B(reg_A[37]), .C(n1767), .D(reg_A[85]), .Y(n2275) );
  NAND2X1 U1743 ( .A(n2276), .B(n2277), .Y(U69_U1_Z_1) );
  AOI22X1 U1744 ( .A(reg_A[94]), .B(n1767), .C(reg_A[46]), .D(n2017), .Y(n2277) );
  AOI22X1 U1745 ( .A(reg_A[14]), .B(n1766), .C(reg_A[118]), .D(n1769), .Y(
        n2276) );
  NAND2X1 U1746 ( .A(n2278), .B(n2279), .Y(U69_U1_Z_0) );
  AOI22X1 U1747 ( .A(reg_A[95]), .B(n1767), .C(reg_A[47]), .D(n1768), .Y(n2279) );
  NOR2X1 U1748 ( .A(n2012), .B(alu_op[2]), .Y(n2017) );
  NOR2X1 U1749 ( .A(n2011), .B(n2012), .Y(n2018) );
  INVX1 U1750 ( .A(ctrl_ww[1]), .Y(n2012) );
  AOI22X1 U1751 ( .A(reg_A[15]), .B(n1766), .C(reg_A[119]), .D(n2049), .Y(
        n2278) );
  NOR2X1 U1752 ( .A(ctrl_ww[1]), .B(alu_op[2]), .Y(n2049) );
  NOR2X1 U1753 ( .A(n2011), .B(ctrl_ww[1]), .Y(n2048) );
endmodule

