
module regfile ( data_out, data_in, wraddr, rdaddr, wren, clk );
  output [7:0] data_out;
  input [7:0] data_in;
  input [7:0] wraddr;
  input [7:0] rdaddr;
  input wren, clk;
  wire   n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657;
  wire   [63:0] reg_file;

  DFFPOSX1 reg_file_reg_0__0_ ( .D(n508), .CLK(clk), .Q(reg_file[0]) );
  DFFPOSX1 reg_file_reg_0__1_ ( .D(n507), .CLK(clk), .Q(reg_file[1]) );
  DFFPOSX1 reg_file_reg_0__2_ ( .D(n506), .CLK(clk), .Q(reg_file[2]) );
  DFFPOSX1 reg_file_reg_0__3_ ( .D(n505), .CLK(clk), .Q(reg_file[3]) );
  DFFPOSX1 reg_file_reg_0__4_ ( .D(n504), .CLK(clk), .Q(reg_file[4]) );
  DFFPOSX1 reg_file_reg_0__5_ ( .D(n503), .CLK(clk), .Q(reg_file[5]) );
  DFFPOSX1 reg_file_reg_0__6_ ( .D(n502), .CLK(clk), .Q(reg_file[6]) );
  DFFPOSX1 reg_file_reg_0__7_ ( .D(n501), .CLK(clk), .Q(reg_file[7]) );
  DFFPOSX1 reg_file_reg_1__0_ ( .D(n500), .CLK(clk), .Q(reg_file[8]) );
  DFFPOSX1 reg_file_reg_1__1_ ( .D(n499), .CLK(clk), .Q(reg_file[9]) );
  DFFPOSX1 reg_file_reg_1__2_ ( .D(n498), .CLK(clk), .Q(reg_file[10]) );
  DFFPOSX1 reg_file_reg_1__3_ ( .D(n497), .CLK(clk), .Q(reg_file[11]) );
  DFFPOSX1 reg_file_reg_1__4_ ( .D(n496), .CLK(clk), .Q(reg_file[12]) );
  DFFPOSX1 reg_file_reg_1__5_ ( .D(n495), .CLK(clk), .Q(reg_file[13]) );
  DFFPOSX1 reg_file_reg_1__6_ ( .D(n494), .CLK(clk), .Q(reg_file[14]) );
  DFFPOSX1 reg_file_reg_1__7_ ( .D(n493), .CLK(clk), .Q(reg_file[15]) );
  DFFPOSX1 reg_file_reg_2__0_ ( .D(n492), .CLK(clk), .Q(reg_file[16]) );
  DFFPOSX1 reg_file_reg_2__1_ ( .D(n491), .CLK(clk), .Q(reg_file[17]) );
  DFFPOSX1 reg_file_reg_2__2_ ( .D(n490), .CLK(clk), .Q(reg_file[18]) );
  DFFPOSX1 reg_file_reg_2__3_ ( .D(n489), .CLK(clk), .Q(reg_file[19]) );
  DFFPOSX1 reg_file_reg_2__4_ ( .D(n488), .CLK(clk), .Q(reg_file[20]) );
  DFFPOSX1 reg_file_reg_2__5_ ( .D(n487), .CLK(clk), .Q(reg_file[21]) );
  DFFPOSX1 reg_file_reg_2__6_ ( .D(n486), .CLK(clk), .Q(reg_file[22]) );
  DFFPOSX1 reg_file_reg_2__7_ ( .D(n485), .CLK(clk), .Q(reg_file[23]) );
  DFFPOSX1 reg_file_reg_3__0_ ( .D(n484), .CLK(clk), .Q(reg_file[24]) );
  DFFPOSX1 reg_file_reg_3__1_ ( .D(n483), .CLK(clk), .Q(reg_file[25]) );
  DFFPOSX1 reg_file_reg_3__2_ ( .D(n482), .CLK(clk), .Q(reg_file[26]) );
  DFFPOSX1 reg_file_reg_3__3_ ( .D(n481), .CLK(clk), .Q(reg_file[27]) );
  DFFPOSX1 reg_file_reg_3__4_ ( .D(n480), .CLK(clk), .Q(reg_file[28]) );
  DFFPOSX1 reg_file_reg_3__5_ ( .D(n479), .CLK(clk), .Q(reg_file[29]) );
  DFFPOSX1 reg_file_reg_3__6_ ( .D(n478), .CLK(clk), .Q(reg_file[30]) );
  DFFPOSX1 reg_file_reg_3__7_ ( .D(n477), .CLK(clk), .Q(reg_file[31]) );
  DFFPOSX1 reg_file_reg_4__0_ ( .D(n476), .CLK(clk), .Q(reg_file[32]) );
  DFFPOSX1 reg_file_reg_4__1_ ( .D(n475), .CLK(clk), .Q(reg_file[33]) );
  DFFPOSX1 reg_file_reg_4__2_ ( .D(n474), .CLK(clk), .Q(reg_file[34]) );
  DFFPOSX1 reg_file_reg_4__3_ ( .D(n473), .CLK(clk), .Q(reg_file[35]) );
  DFFPOSX1 reg_file_reg_4__4_ ( .D(n472), .CLK(clk), .Q(reg_file[36]) );
  DFFPOSX1 reg_file_reg_4__5_ ( .D(n471), .CLK(clk), .Q(reg_file[37]) );
  DFFPOSX1 reg_file_reg_4__6_ ( .D(n470), .CLK(clk), .Q(reg_file[38]) );
  DFFPOSX1 reg_file_reg_4__7_ ( .D(n469), .CLK(clk), .Q(reg_file[39]) );
  DFFPOSX1 reg_file_reg_5__0_ ( .D(n468), .CLK(clk), .Q(reg_file[40]) );
  DFFPOSX1 reg_file_reg_5__1_ ( .D(n467), .CLK(clk), .Q(reg_file[41]) );
  DFFPOSX1 reg_file_reg_5__2_ ( .D(n466), .CLK(clk), .Q(reg_file[42]) );
  DFFPOSX1 reg_file_reg_5__3_ ( .D(n465), .CLK(clk), .Q(reg_file[43]) );
  DFFPOSX1 reg_file_reg_5__4_ ( .D(n464), .CLK(clk), .Q(reg_file[44]) );
  DFFPOSX1 reg_file_reg_5__5_ ( .D(n463), .CLK(clk), .Q(reg_file[45]) );
  DFFPOSX1 reg_file_reg_5__6_ ( .D(n462), .CLK(clk), .Q(reg_file[46]) );
  DFFPOSX1 reg_file_reg_5__7_ ( .D(n461), .CLK(clk), .Q(reg_file[47]) );
  DFFPOSX1 reg_file_reg_6__0_ ( .D(n460), .CLK(clk), .Q(reg_file[48]) );
  DFFPOSX1 reg_file_reg_6__1_ ( .D(n459), .CLK(clk), .Q(reg_file[49]) );
  DFFPOSX1 reg_file_reg_6__2_ ( .D(n458), .CLK(clk), .Q(reg_file[50]) );
  DFFPOSX1 reg_file_reg_6__3_ ( .D(n457), .CLK(clk), .Q(reg_file[51]) );
  DFFPOSX1 reg_file_reg_6__4_ ( .D(n456), .CLK(clk), .Q(reg_file[52]) );
  DFFPOSX1 reg_file_reg_6__5_ ( .D(n455), .CLK(clk), .Q(reg_file[53]) );
  DFFPOSX1 reg_file_reg_6__6_ ( .D(n454), .CLK(clk), .Q(reg_file[54]) );
  DFFPOSX1 reg_file_reg_6__7_ ( .D(n453), .CLK(clk), .Q(reg_file[55]) );
  DFFPOSX1 reg_file_reg_7__0_ ( .D(n452), .CLK(clk), .Q(reg_file[56]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n451), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 reg_file_reg_7__1_ ( .D(n450), .CLK(clk), .Q(reg_file[57]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n449), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 reg_file_reg_7__2_ ( .D(n448), .CLK(clk), .Q(reg_file[58]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n447), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 reg_file_reg_7__3_ ( .D(n446), .CLK(clk), .Q(reg_file[59]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n445), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 reg_file_reg_7__4_ ( .D(n444), .CLK(clk), .Q(reg_file[60]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n443), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 reg_file_reg_7__5_ ( .D(n442), .CLK(clk), .Q(reg_file[61]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n441), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 reg_file_reg_7__6_ ( .D(n440), .CLK(clk), .Q(reg_file[62]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n439), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 reg_file_reg_7__7_ ( .D(n438), .CLK(clk), .Q(reg_file[63]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n437), .CLK(clk), .Q(data_out[7]) );
  MUX2X1 U266 ( .B(n509), .A(n510), .S(n511), .Y(n508) );
  MUX2X1 U267 ( .B(n512), .A(n513), .S(n511), .Y(n507) );
  MUX2X1 U268 ( .B(n514), .A(n515), .S(n511), .Y(n506) );
  MUX2X1 U269 ( .B(n516), .A(n517), .S(n511), .Y(n505) );
  MUX2X1 U270 ( .B(n518), .A(n519), .S(n511), .Y(n504) );
  MUX2X1 U271 ( .B(n520), .A(n521), .S(n511), .Y(n503) );
  MUX2X1 U272 ( .B(n522), .A(n523), .S(n511), .Y(n502) );
  MUX2X1 U273 ( .B(n524), .A(n525), .S(n511), .Y(n501) );
  NAND3X1 U274 ( .A(n526), .B(n527), .C(n528), .Y(n511) );
  MUX2X1 U275 ( .B(n509), .A(n529), .S(n530), .Y(n500) );
  MUX2X1 U276 ( .B(n512), .A(n531), .S(n530), .Y(n499) );
  MUX2X1 U277 ( .B(n514), .A(n532), .S(n530), .Y(n498) );
  MUX2X1 U278 ( .B(n516), .A(n533), .S(n530), .Y(n497) );
  MUX2X1 U279 ( .B(n518), .A(n534), .S(n530), .Y(n496) );
  MUX2X1 U280 ( .B(n520), .A(n535), .S(n530), .Y(n495) );
  MUX2X1 U281 ( .B(n522), .A(n536), .S(n530), .Y(n494) );
  MUX2X1 U282 ( .B(n524), .A(n537), .S(n530), .Y(n493) );
  NAND3X1 U283 ( .A(n528), .B(n527), .C(wraddr[0]), .Y(n530) );
  MUX2X1 U284 ( .B(n509), .A(n538), .S(n539), .Y(n492) );
  MUX2X1 U285 ( .B(n512), .A(n540), .S(n539), .Y(n491) );
  MUX2X1 U286 ( .B(n514), .A(n541), .S(n539), .Y(n490) );
  MUX2X1 U287 ( .B(n516), .A(n542), .S(n539), .Y(n489) );
  MUX2X1 U288 ( .B(n518), .A(n543), .S(n539), .Y(n488) );
  MUX2X1 U289 ( .B(n520), .A(n544), .S(n539), .Y(n487) );
  MUX2X1 U290 ( .B(n522), .A(n545), .S(n539), .Y(n486) );
  MUX2X1 U291 ( .B(n524), .A(n546), .S(n539), .Y(n485) );
  NAND3X1 U292 ( .A(n528), .B(n526), .C(wraddr[1]), .Y(n539) );
  MUX2X1 U293 ( .B(n509), .A(n547), .S(n548), .Y(n484) );
  MUX2X1 U294 ( .B(n512), .A(n549), .S(n548), .Y(n483) );
  MUX2X1 U295 ( .B(n514), .A(n550), .S(n548), .Y(n482) );
  MUX2X1 U296 ( .B(n516), .A(n551), .S(n548), .Y(n481) );
  MUX2X1 U297 ( .B(n518), .A(n552), .S(n548), .Y(n480) );
  MUX2X1 U298 ( .B(n520), .A(n553), .S(n548), .Y(n479) );
  MUX2X1 U299 ( .B(n522), .A(n554), .S(n548), .Y(n478) );
  MUX2X1 U300 ( .B(n524), .A(n555), .S(n548), .Y(n477) );
  NAND3X1 U301 ( .A(wraddr[0]), .B(n528), .C(wraddr[1]), .Y(n548) );
  NOR2X1 U302 ( .A(n556), .B(wraddr[2]), .Y(n528) );
  MUX2X1 U303 ( .B(n509), .A(n557), .S(n558), .Y(n476) );
  MUX2X1 U304 ( .B(n512), .A(n559), .S(n558), .Y(n475) );
  MUX2X1 U305 ( .B(n514), .A(n560), .S(n558), .Y(n474) );
  MUX2X1 U306 ( .B(n516), .A(n561), .S(n558), .Y(n473) );
  MUX2X1 U307 ( .B(n518), .A(n562), .S(n558), .Y(n472) );
  MUX2X1 U308 ( .B(n520), .A(n563), .S(n558), .Y(n471) );
  MUX2X1 U309 ( .B(n522), .A(n564), .S(n558), .Y(n470) );
  MUX2X1 U310 ( .B(n524), .A(n565), .S(n558), .Y(n469) );
  NAND3X1 U311 ( .A(n526), .B(n527), .C(n566), .Y(n558) );
  MUX2X1 U312 ( .B(n509), .A(n567), .S(n568), .Y(n468) );
  MUX2X1 U313 ( .B(n512), .A(n569), .S(n568), .Y(n467) );
  MUX2X1 U314 ( .B(n514), .A(n570), .S(n568), .Y(n466) );
  MUX2X1 U315 ( .B(n516), .A(n571), .S(n568), .Y(n465) );
  MUX2X1 U316 ( .B(n518), .A(n572), .S(n568), .Y(n464) );
  MUX2X1 U317 ( .B(n520), .A(n573), .S(n568), .Y(n463) );
  MUX2X1 U318 ( .B(n522), .A(n574), .S(n568), .Y(n462) );
  MUX2X1 U319 ( .B(n524), .A(n575), .S(n568), .Y(n461) );
  NAND3X1 U320 ( .A(wraddr[0]), .B(n527), .C(n566), .Y(n568) );
  INVX1 U321 ( .A(wraddr[1]), .Y(n527) );
  MUX2X1 U322 ( .B(n509), .A(n576), .S(n577), .Y(n460) );
  MUX2X1 U323 ( .B(n512), .A(n578), .S(n577), .Y(n459) );
  MUX2X1 U324 ( .B(n514), .A(n579), .S(n577), .Y(n458) );
  MUX2X1 U325 ( .B(n516), .A(n580), .S(n577), .Y(n457) );
  MUX2X1 U326 ( .B(n518), .A(n581), .S(n577), .Y(n456) );
  MUX2X1 U327 ( .B(n520), .A(n582), .S(n577), .Y(n455) );
  MUX2X1 U328 ( .B(n522), .A(n583), .S(n577), .Y(n454) );
  MUX2X1 U329 ( .B(n524), .A(n584), .S(n577), .Y(n453) );
  NAND3X1 U330 ( .A(wraddr[1]), .B(n526), .C(n566), .Y(n577) );
  INVX1 U331 ( .A(wraddr[0]), .Y(n526) );
  MUX2X1 U332 ( .B(n509), .A(n585), .S(n586), .Y(n452) );
  INVX1 U333 ( .A(data_in[0]), .Y(n509) );
  NAND3X1 U334 ( .A(n587), .B(n588), .C(n589), .Y(n451) );
  NAND2X1 U335 ( .A(data_out[0]), .B(wren), .Y(n589) );
  OAI21X1 U336 ( .A(n590), .B(n591), .C(n592), .Y(n588) );
  OAI22X1 U337 ( .A(n529), .B(n593), .C(n510), .D(n594), .Y(n591) );
  INVX1 U338 ( .A(reg_file[0]), .Y(n510) );
  INVX1 U339 ( .A(reg_file[8]), .Y(n529) );
  OAI22X1 U340 ( .A(n547), .B(n595), .C(n538), .D(n596), .Y(n590) );
  INVX1 U341 ( .A(reg_file[16]), .Y(n538) );
  INVX1 U342 ( .A(reg_file[24]), .Y(n547) );
  OAI21X1 U343 ( .A(n597), .B(n598), .C(n599), .Y(n587) );
  OAI22X1 U344 ( .A(n567), .B(n593), .C(n557), .D(n594), .Y(n598) );
  INVX1 U345 ( .A(reg_file[32]), .Y(n557) );
  INVX1 U346 ( .A(reg_file[40]), .Y(n567) );
  OAI22X1 U347 ( .A(n585), .B(n595), .C(n576), .D(n596), .Y(n597) );
  INVX1 U348 ( .A(reg_file[48]), .Y(n576) );
  INVX1 U349 ( .A(reg_file[56]), .Y(n585) );
  MUX2X1 U350 ( .B(n512), .A(n600), .S(n586), .Y(n450) );
  INVX1 U351 ( .A(data_in[1]), .Y(n512) );
  NAND3X1 U352 ( .A(n601), .B(n602), .C(n603), .Y(n449) );
  NAND2X1 U353 ( .A(data_out[1]), .B(wren), .Y(n603) );
  OAI21X1 U354 ( .A(n604), .B(n605), .C(n592), .Y(n602) );
  OAI22X1 U355 ( .A(n531), .B(n593), .C(n513), .D(n594), .Y(n605) );
  INVX1 U356 ( .A(reg_file[1]), .Y(n513) );
  INVX1 U357 ( .A(reg_file[9]), .Y(n531) );
  OAI22X1 U358 ( .A(n549), .B(n595), .C(n540), .D(n596), .Y(n604) );
  INVX1 U359 ( .A(reg_file[17]), .Y(n540) );
  INVX1 U360 ( .A(reg_file[25]), .Y(n549) );
  OAI21X1 U361 ( .A(n606), .B(n607), .C(n599), .Y(n601) );
  OAI22X1 U362 ( .A(n569), .B(n593), .C(n559), .D(n594), .Y(n607) );
  INVX1 U363 ( .A(reg_file[33]), .Y(n559) );
  INVX1 U364 ( .A(reg_file[41]), .Y(n569) );
  OAI22X1 U365 ( .A(n595), .B(n600), .C(n578), .D(n596), .Y(n606) );
  INVX1 U366 ( .A(reg_file[49]), .Y(n578) );
  INVX1 U367 ( .A(reg_file[57]), .Y(n600) );
  MUX2X1 U368 ( .B(n514), .A(n608), .S(n586), .Y(n448) );
  INVX1 U369 ( .A(data_in[2]), .Y(n514) );
  NAND3X1 U370 ( .A(n609), .B(n610), .C(n611), .Y(n447) );
  NAND2X1 U371 ( .A(data_out[2]), .B(wren), .Y(n611) );
  OAI21X1 U372 ( .A(n612), .B(n613), .C(n592), .Y(n610) );
  OAI22X1 U373 ( .A(n532), .B(n593), .C(n515), .D(n594), .Y(n613) );
  INVX1 U374 ( .A(reg_file[2]), .Y(n515) );
  INVX1 U375 ( .A(reg_file[10]), .Y(n532) );
  OAI22X1 U376 ( .A(n550), .B(n595), .C(n541), .D(n596), .Y(n612) );
  INVX1 U377 ( .A(reg_file[18]), .Y(n541) );
  INVX1 U378 ( .A(reg_file[26]), .Y(n550) );
  OAI21X1 U379 ( .A(n614), .B(n615), .C(n599), .Y(n609) );
  OAI22X1 U380 ( .A(n570), .B(n593), .C(n560), .D(n594), .Y(n615) );
  INVX1 U381 ( .A(reg_file[34]), .Y(n560) );
  INVX1 U382 ( .A(reg_file[42]), .Y(n570) );
  OAI22X1 U383 ( .A(n595), .B(n608), .C(n579), .D(n596), .Y(n614) );
  INVX1 U384 ( .A(reg_file[50]), .Y(n579) );
  INVX1 U385 ( .A(reg_file[58]), .Y(n608) );
  MUX2X1 U386 ( .B(n516), .A(n616), .S(n586), .Y(n446) );
  INVX1 U387 ( .A(data_in[3]), .Y(n516) );
  NAND3X1 U388 ( .A(n617), .B(n618), .C(n619), .Y(n445) );
  NAND2X1 U389 ( .A(data_out[3]), .B(wren), .Y(n619) );
  OAI21X1 U390 ( .A(n620), .B(n621), .C(n592), .Y(n618) );
  OAI22X1 U391 ( .A(n533), .B(n593), .C(n517), .D(n594), .Y(n621) );
  INVX1 U392 ( .A(reg_file[3]), .Y(n517) );
  INVX1 U393 ( .A(reg_file[11]), .Y(n533) );
  OAI22X1 U394 ( .A(n551), .B(n595), .C(n542), .D(n596), .Y(n620) );
  INVX1 U395 ( .A(reg_file[19]), .Y(n542) );
  INVX1 U396 ( .A(reg_file[27]), .Y(n551) );
  OAI21X1 U397 ( .A(n622), .B(n623), .C(n599), .Y(n617) );
  OAI22X1 U398 ( .A(n571), .B(n593), .C(n561), .D(n594), .Y(n623) );
  INVX1 U399 ( .A(reg_file[35]), .Y(n561) );
  INVX1 U400 ( .A(reg_file[43]), .Y(n571) );
  OAI22X1 U401 ( .A(n595), .B(n616), .C(n580), .D(n596), .Y(n622) );
  INVX1 U402 ( .A(reg_file[51]), .Y(n580) );
  INVX1 U403 ( .A(reg_file[59]), .Y(n616) );
  MUX2X1 U404 ( .B(n518), .A(n624), .S(n586), .Y(n444) );
  INVX1 U405 ( .A(data_in[4]), .Y(n518) );
  NAND3X1 U406 ( .A(n625), .B(n626), .C(n627), .Y(n443) );
  NAND2X1 U407 ( .A(data_out[4]), .B(wren), .Y(n627) );
  OAI21X1 U408 ( .A(n628), .B(n629), .C(n592), .Y(n626) );
  OAI22X1 U409 ( .A(n534), .B(n593), .C(n519), .D(n594), .Y(n629) );
  INVX1 U410 ( .A(reg_file[4]), .Y(n519) );
  INVX1 U411 ( .A(reg_file[12]), .Y(n534) );
  OAI22X1 U412 ( .A(n552), .B(n595), .C(n543), .D(n596), .Y(n628) );
  INVX1 U413 ( .A(reg_file[20]), .Y(n543) );
  INVX1 U414 ( .A(reg_file[28]), .Y(n552) );
  OAI21X1 U415 ( .A(n630), .B(n631), .C(n599), .Y(n625) );
  OAI22X1 U416 ( .A(n572), .B(n593), .C(n562), .D(n594), .Y(n631) );
  INVX1 U417 ( .A(reg_file[36]), .Y(n562) );
  INVX1 U418 ( .A(reg_file[44]), .Y(n572) );
  OAI22X1 U419 ( .A(n595), .B(n624), .C(n581), .D(n596), .Y(n630) );
  INVX1 U420 ( .A(reg_file[52]), .Y(n581) );
  INVX1 U421 ( .A(reg_file[60]), .Y(n624) );
  MUX2X1 U422 ( .B(n520), .A(n632), .S(n586), .Y(n442) );
  INVX1 U423 ( .A(data_in[5]), .Y(n520) );
  NAND3X1 U424 ( .A(n633), .B(n634), .C(n635), .Y(n441) );
  NAND2X1 U425 ( .A(data_out[5]), .B(wren), .Y(n635) );
  OAI21X1 U426 ( .A(n636), .B(n637), .C(n592), .Y(n634) );
  OAI22X1 U427 ( .A(n535), .B(n593), .C(n521), .D(n594), .Y(n637) );
  INVX1 U428 ( .A(reg_file[5]), .Y(n521) );
  INVX1 U429 ( .A(reg_file[13]), .Y(n535) );
  OAI22X1 U430 ( .A(n553), .B(n595), .C(n544), .D(n596), .Y(n636) );
  INVX1 U431 ( .A(reg_file[21]), .Y(n544) );
  INVX1 U432 ( .A(reg_file[29]), .Y(n553) );
  OAI21X1 U433 ( .A(n638), .B(n639), .C(n599), .Y(n633) );
  OAI22X1 U434 ( .A(n573), .B(n593), .C(n563), .D(n594), .Y(n639) );
  INVX1 U435 ( .A(reg_file[37]), .Y(n563) );
  INVX1 U436 ( .A(reg_file[45]), .Y(n573) );
  OAI22X1 U437 ( .A(n595), .B(n632), .C(n582), .D(n596), .Y(n638) );
  INVX1 U438 ( .A(reg_file[53]), .Y(n582) );
  INVX1 U439 ( .A(reg_file[61]), .Y(n632) );
  MUX2X1 U440 ( .B(n522), .A(n640), .S(n586), .Y(n440) );
  INVX1 U441 ( .A(data_in[6]), .Y(n522) );
  NAND3X1 U442 ( .A(n641), .B(n642), .C(n643), .Y(n439) );
  NAND2X1 U443 ( .A(data_out[6]), .B(wren), .Y(n643) );
  OAI21X1 U444 ( .A(n644), .B(n645), .C(n592), .Y(n642) );
  OAI22X1 U445 ( .A(n536), .B(n593), .C(n523), .D(n594), .Y(n645) );
  INVX1 U446 ( .A(reg_file[6]), .Y(n523) );
  INVX1 U447 ( .A(reg_file[14]), .Y(n536) );
  OAI22X1 U448 ( .A(n554), .B(n595), .C(n545), .D(n596), .Y(n644) );
  INVX1 U449 ( .A(reg_file[22]), .Y(n545) );
  INVX1 U450 ( .A(reg_file[30]), .Y(n554) );
  OAI21X1 U451 ( .A(n646), .B(n647), .C(n599), .Y(n641) );
  OAI22X1 U452 ( .A(n574), .B(n593), .C(n564), .D(n594), .Y(n647) );
  INVX1 U453 ( .A(reg_file[38]), .Y(n564) );
  INVX1 U454 ( .A(reg_file[46]), .Y(n574) );
  OAI22X1 U455 ( .A(n595), .B(n640), .C(n583), .D(n596), .Y(n646) );
  INVX1 U456 ( .A(reg_file[54]), .Y(n583) );
  INVX1 U457 ( .A(reg_file[62]), .Y(n640) );
  MUX2X1 U458 ( .B(n524), .A(n648), .S(n586), .Y(n438) );
  NAND3X1 U459 ( .A(wraddr[1]), .B(wraddr[0]), .C(n566), .Y(n586) );
  AND2X1 U460 ( .A(wraddr[2]), .B(wren), .Y(n566) );
  INVX1 U461 ( .A(data_in[7]), .Y(n524) );
  NAND3X1 U462 ( .A(n649), .B(n650), .C(n651), .Y(n437) );
  NAND2X1 U463 ( .A(data_out[7]), .B(wren), .Y(n651) );
  OAI21X1 U464 ( .A(n652), .B(n653), .C(n592), .Y(n650) );
  NOR2X1 U465 ( .A(wren), .B(rdaddr[2]), .Y(n592) );
  OAI22X1 U466 ( .A(n537), .B(n593), .C(n525), .D(n594), .Y(n653) );
  INVX1 U467 ( .A(reg_file[7]), .Y(n525) );
  INVX1 U468 ( .A(reg_file[15]), .Y(n537) );
  OAI22X1 U469 ( .A(n555), .B(n595), .C(n546), .D(n596), .Y(n652) );
  INVX1 U470 ( .A(reg_file[23]), .Y(n546) );
  INVX1 U471 ( .A(reg_file[31]), .Y(n555) );
  OAI21X1 U472 ( .A(n654), .B(n655), .C(n599), .Y(n649) );
  AND2X1 U473 ( .A(rdaddr[2]), .B(n556), .Y(n599) );
  INVX1 U474 ( .A(wren), .Y(n556) );
  OAI22X1 U475 ( .A(n575), .B(n593), .C(n565), .D(n594), .Y(n655) );
  NAND2X1 U476 ( .A(n656), .B(n657), .Y(n594) );
  INVX1 U477 ( .A(reg_file[39]), .Y(n565) );
  NAND2X1 U478 ( .A(rdaddr[0]), .B(n656), .Y(n593) );
  INVX1 U479 ( .A(rdaddr[1]), .Y(n656) );
  INVX1 U480 ( .A(reg_file[47]), .Y(n575) );
  OAI22X1 U481 ( .A(n595), .B(n648), .C(n584), .D(n596), .Y(n654) );
  NAND2X1 U482 ( .A(rdaddr[1]), .B(n657), .Y(n596) );
  INVX1 U483 ( .A(rdaddr[0]), .Y(n657) );
  INVX1 U484 ( .A(reg_file[55]), .Y(n584) );
  INVX1 U485 ( .A(reg_file[63]), .Y(n648) );
  NAND2X1 U486 ( .A(rdaddr[0]), .B(rdaddr[1]), .Y(n595) );
endmodule

