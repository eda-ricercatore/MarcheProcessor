
module regfile ( data_out, data_in, wraddr, rdaddr, wren, clk );
  output [7:0] data_out;
  input [7:0] data_in;
  input [7:0] wraddr;
  input [7:0] rdaddr;
  input wren, clk;
  wire   n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048;
  wire   [63:0] reg_file;

  DFFPOSX1 reg_file_reg_0__0_ ( .D(n508), .CLK(clk), .Q(reg_file[0]) );
  DFFPOSX1 reg_file_reg_0__1_ ( .D(n507), .CLK(clk), .Q(reg_file[1]) );
  DFFPOSX1 reg_file_reg_0__2_ ( .D(n506), .CLK(clk), .Q(reg_file[2]) );
  DFFPOSX1 reg_file_reg_0__3_ ( .D(n505), .CLK(clk), .Q(reg_file[3]) );
  DFFPOSX1 reg_file_reg_0__4_ ( .D(n504), .CLK(clk), .Q(reg_file[4]) );
  DFFPOSX1 reg_file_reg_0__5_ ( .D(n503), .CLK(clk), .Q(reg_file[5]) );
  DFFPOSX1 reg_file_reg_0__6_ ( .D(n502), .CLK(clk), .Q(reg_file[6]) );
  DFFPOSX1 reg_file_reg_0__7_ ( .D(n501), .CLK(clk), .Q(reg_file[7]) );
  DFFPOSX1 reg_file_reg_1__0_ ( .D(n500), .CLK(clk), .Q(reg_file[8]) );
  DFFPOSX1 reg_file_reg_1__1_ ( .D(n499), .CLK(clk), .Q(reg_file[9]) );
  DFFPOSX1 reg_file_reg_1__2_ ( .D(n498), .CLK(clk), .Q(reg_file[10]) );
  DFFPOSX1 reg_file_reg_1__3_ ( .D(n497), .CLK(clk), .Q(reg_file[11]) );
  DFFPOSX1 reg_file_reg_1__4_ ( .D(n496), .CLK(clk), .Q(reg_file[12]) );
  DFFPOSX1 reg_file_reg_1__5_ ( .D(n495), .CLK(clk), .Q(reg_file[13]) );
  DFFPOSX1 reg_file_reg_1__6_ ( .D(n494), .CLK(clk), .Q(reg_file[14]) );
  DFFPOSX1 reg_file_reg_1__7_ ( .D(n493), .CLK(clk), .Q(reg_file[15]) );
  DFFPOSX1 reg_file_reg_2__0_ ( .D(n492), .CLK(clk), .Q(reg_file[16]) );
  DFFPOSX1 reg_file_reg_2__1_ ( .D(n491), .CLK(clk), .Q(reg_file[17]) );
  DFFPOSX1 reg_file_reg_2__2_ ( .D(n490), .CLK(clk), .Q(reg_file[18]) );
  DFFPOSX1 reg_file_reg_2__3_ ( .D(n489), .CLK(clk), .Q(reg_file[19]) );
  DFFPOSX1 reg_file_reg_2__4_ ( .D(n488), .CLK(clk), .Q(reg_file[20]) );
  DFFPOSX1 reg_file_reg_2__5_ ( .D(n487), .CLK(clk), .Q(reg_file[21]) );
  DFFPOSX1 reg_file_reg_2__6_ ( .D(n486), .CLK(clk), .Q(reg_file[22]) );
  DFFPOSX1 reg_file_reg_2__7_ ( .D(n485), .CLK(clk), .Q(reg_file[23]) );
  DFFPOSX1 reg_file_reg_3__0_ ( .D(n484), .CLK(clk), .Q(reg_file[24]) );
  DFFPOSX1 reg_file_reg_3__1_ ( .D(n483), .CLK(clk), .Q(reg_file[25]) );
  DFFPOSX1 reg_file_reg_3__2_ ( .D(n482), .CLK(clk), .Q(reg_file[26]) );
  DFFPOSX1 reg_file_reg_3__3_ ( .D(n481), .CLK(clk), .Q(reg_file[27]) );
  DFFPOSX1 reg_file_reg_3__4_ ( .D(n480), .CLK(clk), .Q(reg_file[28]) );
  DFFPOSX1 reg_file_reg_3__5_ ( .D(n479), .CLK(clk), .Q(reg_file[29]) );
  DFFPOSX1 reg_file_reg_3__6_ ( .D(n478), .CLK(clk), .Q(reg_file[30]) );
  DFFPOSX1 reg_file_reg_3__7_ ( .D(n477), .CLK(clk), .Q(reg_file[31]) );
  DFFPOSX1 reg_file_reg_4__0_ ( .D(n476), .CLK(clk), .Q(reg_file[32]) );
  DFFPOSX1 reg_file_reg_4__1_ ( .D(n475), .CLK(clk), .Q(reg_file[33]) );
  DFFPOSX1 reg_file_reg_4__2_ ( .D(n474), .CLK(clk), .Q(reg_file[34]) );
  DFFPOSX1 reg_file_reg_4__3_ ( .D(n473), .CLK(clk), .Q(reg_file[35]) );
  DFFPOSX1 reg_file_reg_4__4_ ( .D(n472), .CLK(clk), .Q(reg_file[36]) );
  DFFPOSX1 reg_file_reg_4__5_ ( .D(n471), .CLK(clk), .Q(reg_file[37]) );
  DFFPOSX1 reg_file_reg_4__6_ ( .D(n470), .CLK(clk), .Q(reg_file[38]) );
  DFFPOSX1 reg_file_reg_4__7_ ( .D(n469), .CLK(clk), .Q(reg_file[39]) );
  DFFPOSX1 reg_file_reg_5__0_ ( .D(n468), .CLK(clk), .Q(reg_file[40]) );
  DFFPOSX1 reg_file_reg_5__1_ ( .D(n467), .CLK(clk), .Q(reg_file[41]) );
  DFFPOSX1 reg_file_reg_5__2_ ( .D(n466), .CLK(clk), .Q(reg_file[42]) );
  DFFPOSX1 reg_file_reg_5__3_ ( .D(n465), .CLK(clk), .Q(reg_file[43]) );
  DFFPOSX1 reg_file_reg_5__4_ ( .D(n464), .CLK(clk), .Q(reg_file[44]) );
  DFFPOSX1 reg_file_reg_5__5_ ( .D(n463), .CLK(clk), .Q(reg_file[45]) );
  DFFPOSX1 reg_file_reg_5__6_ ( .D(n462), .CLK(clk), .Q(reg_file[46]) );
  DFFPOSX1 reg_file_reg_5__7_ ( .D(n461), .CLK(clk), .Q(reg_file[47]) );
  DFFPOSX1 reg_file_reg_6__0_ ( .D(n460), .CLK(clk), .Q(reg_file[48]) );
  DFFPOSX1 reg_file_reg_6__1_ ( .D(n459), .CLK(clk), .Q(reg_file[49]) );
  DFFPOSX1 reg_file_reg_6__2_ ( .D(n458), .CLK(clk), .Q(reg_file[50]) );
  DFFPOSX1 reg_file_reg_6__3_ ( .D(n457), .CLK(clk), .Q(reg_file[51]) );
  DFFPOSX1 reg_file_reg_6__4_ ( .D(n456), .CLK(clk), .Q(reg_file[52]) );
  DFFPOSX1 reg_file_reg_6__5_ ( .D(n455), .CLK(clk), .Q(reg_file[53]) );
  DFFPOSX1 reg_file_reg_6__6_ ( .D(n454), .CLK(clk), .Q(reg_file[54]) );
  DFFPOSX1 reg_file_reg_6__7_ ( .D(n453), .CLK(clk), .Q(reg_file[55]) );
  DFFPOSX1 reg_file_reg_7__0_ ( .D(n452), .CLK(clk), .Q(reg_file[56]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n451), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 reg_file_reg_7__1_ ( .D(n450), .CLK(clk), .Q(reg_file[57]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n449), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 reg_file_reg_7__2_ ( .D(n448), .CLK(clk), .Q(reg_file[58]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n447), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 reg_file_reg_7__3_ ( .D(n446), .CLK(clk), .Q(reg_file[59]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n445), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 reg_file_reg_7__4_ ( .D(n444), .CLK(clk), .Q(reg_file[60]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n443), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 reg_file_reg_7__5_ ( .D(n442), .CLK(clk), .Q(reg_file[61]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n441), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 reg_file_reg_7__6_ ( .D(n440), .CLK(clk), .Q(reg_file[62]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n439), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 reg_file_reg_7__7_ ( .D(n438), .CLK(clk), .Q(reg_file[63]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n437), .CLK(clk), .Q(data_out[7]) );
  MUX2X1 U495 ( .B(n900), .A(n901), .S(n902), .Y(n508) );
  MUX2X1 U496 ( .B(n903), .A(n904), .S(n902), .Y(n507) );
  MUX2X1 U497 ( .B(n905), .A(n906), .S(n902), .Y(n506) );
  MUX2X1 U498 ( .B(n907), .A(n908), .S(n902), .Y(n505) );
  MUX2X1 U499 ( .B(n909), .A(n910), .S(n902), .Y(n504) );
  MUX2X1 U500 ( .B(n911), .A(n912), .S(n902), .Y(n503) );
  MUX2X1 U501 ( .B(n913), .A(n914), .S(n902), .Y(n502) );
  MUX2X1 U502 ( .B(n915), .A(n916), .S(n902), .Y(n501) );
  NAND3X1 U503 ( .A(n917), .B(n918), .C(n919), .Y(n902) );
  MUX2X1 U504 ( .B(n900), .A(n920), .S(n921), .Y(n500) );
  MUX2X1 U505 ( .B(n903), .A(n922), .S(n921), .Y(n499) );
  MUX2X1 U506 ( .B(n905), .A(n923), .S(n921), .Y(n498) );
  MUX2X1 U507 ( .B(n907), .A(n924), .S(n921), .Y(n497) );
  MUX2X1 U508 ( .B(n909), .A(n925), .S(n921), .Y(n496) );
  MUX2X1 U509 ( .B(n911), .A(n926), .S(n921), .Y(n495) );
  MUX2X1 U510 ( .B(n913), .A(n927), .S(n921), .Y(n494) );
  MUX2X1 U511 ( .B(n915), .A(n928), .S(n921), .Y(n493) );
  NAND3X1 U512 ( .A(n919), .B(n918), .C(wraddr[0]), .Y(n921) );
  MUX2X1 U513 ( .B(n900), .A(n929), .S(n930), .Y(n492) );
  MUX2X1 U514 ( .B(n903), .A(n931), .S(n930), .Y(n491) );
  MUX2X1 U515 ( .B(n905), .A(n932), .S(n930), .Y(n490) );
  MUX2X1 U516 ( .B(n907), .A(n933), .S(n930), .Y(n489) );
  MUX2X1 U517 ( .B(n909), .A(n934), .S(n930), .Y(n488) );
  MUX2X1 U518 ( .B(n911), .A(n935), .S(n930), .Y(n487) );
  MUX2X1 U519 ( .B(n913), .A(n936), .S(n930), .Y(n486) );
  MUX2X1 U520 ( .B(n915), .A(n937), .S(n930), .Y(n485) );
  NAND3X1 U521 ( .A(n919), .B(n917), .C(wraddr[1]), .Y(n930) );
  MUX2X1 U522 ( .B(n900), .A(n938), .S(n939), .Y(n484) );
  MUX2X1 U523 ( .B(n903), .A(n940), .S(n939), .Y(n483) );
  MUX2X1 U524 ( .B(n905), .A(n941), .S(n939), .Y(n482) );
  MUX2X1 U525 ( .B(n907), .A(n942), .S(n939), .Y(n481) );
  MUX2X1 U526 ( .B(n909), .A(n943), .S(n939), .Y(n480) );
  MUX2X1 U527 ( .B(n911), .A(n944), .S(n939), .Y(n479) );
  MUX2X1 U528 ( .B(n913), .A(n945), .S(n939), .Y(n478) );
  MUX2X1 U529 ( .B(n915), .A(n946), .S(n939), .Y(n477) );
  NAND3X1 U530 ( .A(wraddr[0]), .B(n919), .C(wraddr[1]), .Y(n939) );
  NOR2X1 U531 ( .A(n947), .B(wraddr[2]), .Y(n919) );
  MUX2X1 U532 ( .B(n900), .A(n948), .S(n949), .Y(n476) );
  MUX2X1 U533 ( .B(n903), .A(n950), .S(n949), .Y(n475) );
  MUX2X1 U534 ( .B(n905), .A(n951), .S(n949), .Y(n474) );
  MUX2X1 U535 ( .B(n907), .A(n952), .S(n949), .Y(n473) );
  MUX2X1 U536 ( .B(n909), .A(n953), .S(n949), .Y(n472) );
  MUX2X1 U537 ( .B(n911), .A(n954), .S(n949), .Y(n471) );
  MUX2X1 U538 ( .B(n913), .A(n955), .S(n949), .Y(n470) );
  MUX2X1 U539 ( .B(n915), .A(n956), .S(n949), .Y(n469) );
  NAND3X1 U540 ( .A(n917), .B(n918), .C(n957), .Y(n949) );
  MUX2X1 U541 ( .B(n900), .A(n958), .S(n959), .Y(n468) );
  MUX2X1 U542 ( .B(n903), .A(n960), .S(n959), .Y(n467) );
  MUX2X1 U543 ( .B(n905), .A(n961), .S(n959), .Y(n466) );
  MUX2X1 U544 ( .B(n907), .A(n962), .S(n959), .Y(n465) );
  MUX2X1 U545 ( .B(n909), .A(n963), .S(n959), .Y(n464) );
  MUX2X1 U546 ( .B(n911), .A(n964), .S(n959), .Y(n463) );
  MUX2X1 U547 ( .B(n913), .A(n965), .S(n959), .Y(n462) );
  MUX2X1 U548 ( .B(n915), .A(n966), .S(n959), .Y(n461) );
  NAND3X1 U549 ( .A(wraddr[0]), .B(n918), .C(n957), .Y(n959) );
  INVX1 U550 ( .A(wraddr[1]), .Y(n918) );
  MUX2X1 U551 ( .B(n900), .A(n967), .S(n968), .Y(n460) );
  MUX2X1 U552 ( .B(n903), .A(n969), .S(n968), .Y(n459) );
  MUX2X1 U553 ( .B(n905), .A(n970), .S(n968), .Y(n458) );
  MUX2X1 U554 ( .B(n907), .A(n971), .S(n968), .Y(n457) );
  MUX2X1 U555 ( .B(n909), .A(n972), .S(n968), .Y(n456) );
  MUX2X1 U556 ( .B(n911), .A(n973), .S(n968), .Y(n455) );
  MUX2X1 U557 ( .B(n913), .A(n974), .S(n968), .Y(n454) );
  MUX2X1 U558 ( .B(n915), .A(n975), .S(n968), .Y(n453) );
  NAND3X1 U559 ( .A(wraddr[1]), .B(n917), .C(n957), .Y(n968) );
  INVX1 U560 ( .A(wraddr[0]), .Y(n917) );
  MUX2X1 U561 ( .B(n900), .A(n976), .S(n977), .Y(n452) );
  INVX1 U562 ( .A(data_in[0]), .Y(n900) );
  NAND3X1 U563 ( .A(n978), .B(n979), .C(n980), .Y(n451) );
  NAND2X1 U564 ( .A(data_out[0]), .B(wren), .Y(n980) );
  OAI21X1 U565 ( .A(n981), .B(n982), .C(n983), .Y(n979) );
  OAI22X1 U566 ( .A(n920), .B(n984), .C(n901), .D(n985), .Y(n982) );
  INVX1 U567 ( .A(reg_file[0]), .Y(n901) );
  INVX1 U568 ( .A(reg_file[8]), .Y(n920) );
  OAI22X1 U569 ( .A(n938), .B(n986), .C(n929), .D(n987), .Y(n981) );
  INVX1 U570 ( .A(reg_file[16]), .Y(n929) );
  INVX1 U571 ( .A(reg_file[24]), .Y(n938) );
  OAI21X1 U572 ( .A(n988), .B(n989), .C(n990), .Y(n978) );
  OAI22X1 U573 ( .A(n958), .B(n984), .C(n948), .D(n985), .Y(n989) );
  INVX1 U574 ( .A(reg_file[32]), .Y(n948) );
  INVX1 U575 ( .A(reg_file[40]), .Y(n958) );
  OAI22X1 U576 ( .A(n976), .B(n986), .C(n967), .D(n987), .Y(n988) );
  INVX1 U577 ( .A(reg_file[48]), .Y(n967) );
  INVX1 U578 ( .A(reg_file[56]), .Y(n976) );
  MUX2X1 U579 ( .B(n903), .A(n991), .S(n977), .Y(n450) );
  INVX1 U580 ( .A(data_in[1]), .Y(n903) );
  NAND3X1 U581 ( .A(n992), .B(n993), .C(n994), .Y(n449) );
  NAND2X1 U582 ( .A(data_out[1]), .B(wren), .Y(n994) );
  OAI21X1 U583 ( .A(n995), .B(n996), .C(n983), .Y(n993) );
  OAI22X1 U584 ( .A(n922), .B(n984), .C(n904), .D(n985), .Y(n996) );
  INVX1 U585 ( .A(reg_file[1]), .Y(n904) );
  INVX1 U586 ( .A(reg_file[9]), .Y(n922) );
  OAI22X1 U587 ( .A(n940), .B(n986), .C(n931), .D(n987), .Y(n995) );
  INVX1 U588 ( .A(reg_file[17]), .Y(n931) );
  INVX1 U589 ( .A(reg_file[25]), .Y(n940) );
  OAI21X1 U590 ( .A(n997), .B(n998), .C(n990), .Y(n992) );
  OAI22X1 U591 ( .A(n960), .B(n984), .C(n950), .D(n985), .Y(n998) );
  INVX1 U592 ( .A(reg_file[33]), .Y(n950) );
  INVX1 U593 ( .A(reg_file[41]), .Y(n960) );
  OAI22X1 U594 ( .A(n986), .B(n991), .C(n969), .D(n987), .Y(n997) );
  INVX1 U595 ( .A(reg_file[49]), .Y(n969) );
  INVX1 U596 ( .A(reg_file[57]), .Y(n991) );
  MUX2X1 U597 ( .B(n905), .A(n999), .S(n977), .Y(n448) );
  INVX1 U598 ( .A(data_in[2]), .Y(n905) );
  NAND3X1 U599 ( .A(n1000), .B(n1001), .C(n1002), .Y(n447) );
  NAND2X1 U600 ( .A(data_out[2]), .B(wren), .Y(n1002) );
  OAI21X1 U601 ( .A(n1003), .B(n1004), .C(n983), .Y(n1001) );
  OAI22X1 U602 ( .A(n923), .B(n984), .C(n906), .D(n985), .Y(n1004) );
  INVX1 U603 ( .A(reg_file[2]), .Y(n906) );
  INVX1 U604 ( .A(reg_file[10]), .Y(n923) );
  OAI22X1 U605 ( .A(n941), .B(n986), .C(n932), .D(n987), .Y(n1003) );
  INVX1 U606 ( .A(reg_file[18]), .Y(n932) );
  INVX1 U607 ( .A(reg_file[26]), .Y(n941) );
  OAI21X1 U608 ( .A(n1005), .B(n1006), .C(n990), .Y(n1000) );
  OAI22X1 U609 ( .A(n961), .B(n984), .C(n951), .D(n985), .Y(n1006) );
  INVX1 U610 ( .A(reg_file[34]), .Y(n951) );
  INVX1 U611 ( .A(reg_file[42]), .Y(n961) );
  OAI22X1 U612 ( .A(n986), .B(n999), .C(n970), .D(n987), .Y(n1005) );
  INVX1 U613 ( .A(reg_file[50]), .Y(n970) );
  INVX1 U614 ( .A(reg_file[58]), .Y(n999) );
  MUX2X1 U615 ( .B(n907), .A(n1007), .S(n977), .Y(n446) );
  INVX1 U616 ( .A(data_in[3]), .Y(n907) );
  NAND3X1 U617 ( .A(n1008), .B(n1009), .C(n1010), .Y(n445) );
  NAND2X1 U618 ( .A(data_out[3]), .B(wren), .Y(n1010) );
  OAI21X1 U619 ( .A(n1011), .B(n1012), .C(n983), .Y(n1009) );
  OAI22X1 U620 ( .A(n924), .B(n984), .C(n908), .D(n985), .Y(n1012) );
  INVX1 U621 ( .A(reg_file[3]), .Y(n908) );
  INVX1 U622 ( .A(reg_file[11]), .Y(n924) );
  OAI22X1 U623 ( .A(n942), .B(n986), .C(n933), .D(n987), .Y(n1011) );
  INVX1 U624 ( .A(reg_file[19]), .Y(n933) );
  INVX1 U625 ( .A(reg_file[27]), .Y(n942) );
  OAI21X1 U626 ( .A(n1013), .B(n1014), .C(n990), .Y(n1008) );
  OAI22X1 U627 ( .A(n962), .B(n984), .C(n952), .D(n985), .Y(n1014) );
  INVX1 U628 ( .A(reg_file[35]), .Y(n952) );
  INVX1 U629 ( .A(reg_file[43]), .Y(n962) );
  OAI22X1 U630 ( .A(n986), .B(n1007), .C(n971), .D(n987), .Y(n1013) );
  INVX1 U631 ( .A(reg_file[51]), .Y(n971) );
  INVX1 U632 ( .A(reg_file[59]), .Y(n1007) );
  MUX2X1 U633 ( .B(n909), .A(n1015), .S(n977), .Y(n444) );
  INVX1 U634 ( .A(data_in[4]), .Y(n909) );
  NAND3X1 U635 ( .A(n1016), .B(n1017), .C(n1018), .Y(n443) );
  NAND2X1 U636 ( .A(data_out[4]), .B(wren), .Y(n1018) );
  OAI21X1 U637 ( .A(n1019), .B(n1020), .C(n983), .Y(n1017) );
  OAI22X1 U638 ( .A(n925), .B(n984), .C(n910), .D(n985), .Y(n1020) );
  INVX1 U639 ( .A(reg_file[4]), .Y(n910) );
  INVX1 U640 ( .A(reg_file[12]), .Y(n925) );
  OAI22X1 U641 ( .A(n943), .B(n986), .C(n934), .D(n987), .Y(n1019) );
  INVX1 U642 ( .A(reg_file[20]), .Y(n934) );
  INVX1 U643 ( .A(reg_file[28]), .Y(n943) );
  OAI21X1 U644 ( .A(n1021), .B(n1022), .C(n990), .Y(n1016) );
  OAI22X1 U645 ( .A(n963), .B(n984), .C(n953), .D(n985), .Y(n1022) );
  INVX1 U646 ( .A(reg_file[36]), .Y(n953) );
  INVX1 U647 ( .A(reg_file[44]), .Y(n963) );
  OAI22X1 U648 ( .A(n986), .B(n1015), .C(n972), .D(n987), .Y(n1021) );
  INVX1 U649 ( .A(reg_file[52]), .Y(n972) );
  INVX1 U650 ( .A(reg_file[60]), .Y(n1015) );
  MUX2X1 U651 ( .B(n911), .A(n1023), .S(n977), .Y(n442) );
  INVX1 U652 ( .A(data_in[5]), .Y(n911) );
  NAND3X1 U653 ( .A(n1024), .B(n1025), .C(n1026), .Y(n441) );
  NAND2X1 U654 ( .A(data_out[5]), .B(wren), .Y(n1026) );
  OAI21X1 U655 ( .A(n1027), .B(n1028), .C(n983), .Y(n1025) );
  OAI22X1 U656 ( .A(n926), .B(n984), .C(n912), .D(n985), .Y(n1028) );
  INVX1 U657 ( .A(reg_file[5]), .Y(n912) );
  INVX1 U658 ( .A(reg_file[13]), .Y(n926) );
  OAI22X1 U659 ( .A(n944), .B(n986), .C(n935), .D(n987), .Y(n1027) );
  INVX1 U660 ( .A(reg_file[21]), .Y(n935) );
  INVX1 U661 ( .A(reg_file[29]), .Y(n944) );
  OAI21X1 U662 ( .A(n1029), .B(n1030), .C(n990), .Y(n1024) );
  OAI22X1 U663 ( .A(n964), .B(n984), .C(n954), .D(n985), .Y(n1030) );
  INVX1 U664 ( .A(reg_file[37]), .Y(n954) );
  INVX1 U665 ( .A(reg_file[45]), .Y(n964) );
  OAI22X1 U666 ( .A(n986), .B(n1023), .C(n973), .D(n987), .Y(n1029) );
  INVX1 U667 ( .A(reg_file[53]), .Y(n973) );
  INVX1 U668 ( .A(reg_file[61]), .Y(n1023) );
  MUX2X1 U669 ( .B(n913), .A(n1031), .S(n977), .Y(n440) );
  INVX1 U670 ( .A(data_in[6]), .Y(n913) );
  NAND3X1 U671 ( .A(n1032), .B(n1033), .C(n1034), .Y(n439) );
  NAND2X1 U672 ( .A(data_out[6]), .B(wren), .Y(n1034) );
  OAI21X1 U673 ( .A(n1035), .B(n1036), .C(n983), .Y(n1033) );
  OAI22X1 U674 ( .A(n927), .B(n984), .C(n914), .D(n985), .Y(n1036) );
  INVX1 U675 ( .A(reg_file[6]), .Y(n914) );
  INVX1 U676 ( .A(reg_file[14]), .Y(n927) );
  OAI22X1 U677 ( .A(n945), .B(n986), .C(n936), .D(n987), .Y(n1035) );
  INVX1 U678 ( .A(reg_file[22]), .Y(n936) );
  INVX1 U679 ( .A(reg_file[30]), .Y(n945) );
  OAI21X1 U680 ( .A(n1037), .B(n1038), .C(n990), .Y(n1032) );
  OAI22X1 U681 ( .A(n965), .B(n984), .C(n955), .D(n985), .Y(n1038) );
  INVX1 U682 ( .A(reg_file[38]), .Y(n955) );
  INVX1 U683 ( .A(reg_file[46]), .Y(n965) );
  OAI22X1 U684 ( .A(n986), .B(n1031), .C(n974), .D(n987), .Y(n1037) );
  INVX1 U685 ( .A(reg_file[54]), .Y(n974) );
  INVX1 U686 ( .A(reg_file[62]), .Y(n1031) );
  MUX2X1 U687 ( .B(n915), .A(n1039), .S(n977), .Y(n438) );
  NAND3X1 U688 ( .A(wraddr[1]), .B(wraddr[0]), .C(n957), .Y(n977) );
  AND2X1 U689 ( .A(wraddr[2]), .B(wren), .Y(n957) );
  INVX1 U690 ( .A(data_in[7]), .Y(n915) );
  NAND3X1 U691 ( .A(n1040), .B(n1041), .C(n1042), .Y(n437) );
  NAND2X1 U692 ( .A(data_out[7]), .B(wren), .Y(n1042) );
  OAI21X1 U693 ( .A(n1043), .B(n1044), .C(n983), .Y(n1041) );
  NOR2X1 U694 ( .A(rdaddr[2]), .B(wren), .Y(n983) );
  OAI22X1 U695 ( .A(n928), .B(n984), .C(n916), .D(n985), .Y(n1044) );
  INVX1 U696 ( .A(reg_file[7]), .Y(n916) );
  INVX1 U697 ( .A(reg_file[15]), .Y(n928) );
  OAI22X1 U698 ( .A(n946), .B(n986), .C(n937), .D(n987), .Y(n1043) );
  INVX1 U699 ( .A(reg_file[23]), .Y(n937) );
  INVX1 U700 ( .A(reg_file[31]), .Y(n946) );
  OAI21X1 U701 ( .A(n1045), .B(n1046), .C(n990), .Y(n1040) );
  AND2X1 U702 ( .A(rdaddr[2]), .B(n947), .Y(n990) );
  INVX1 U703 ( .A(wren), .Y(n947) );
  OAI22X1 U704 ( .A(n966), .B(n984), .C(n956), .D(n985), .Y(n1046) );
  NAND2X1 U705 ( .A(n1047), .B(n1048), .Y(n985) );
  INVX1 U706 ( .A(reg_file[39]), .Y(n956) );
  NAND2X1 U707 ( .A(rdaddr[0]), .B(n1047), .Y(n984) );
  INVX1 U708 ( .A(rdaddr[1]), .Y(n1047) );
  INVX1 U709 ( .A(reg_file[47]), .Y(n966) );
  OAI22X1 U710 ( .A(n986), .B(n1039), .C(n975), .D(n987), .Y(n1045) );
  NAND2X1 U711 ( .A(rdaddr[1]), .B(n1048), .Y(n987) );
  INVX1 U712 ( .A(rdaddr[0]), .Y(n1048) );
  INVX1 U713 ( .A(reg_file[55]), .Y(n975) );
  INVX1 U714 ( .A(reg_file[63]), .Y(n1039) );
  NAND2X1 U715 ( .A(rdaddr[0]), .B(rdaddr[1]), .Y(n986) );
endmodule

