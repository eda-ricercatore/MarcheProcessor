/**
 * This is written by Zhiyang Ong (zhiyango@usc.edu; 6004 9194 12)
 * and Andrew Mattheisen (mattheis@usc.edu; 2134 5147 11)
 * for EE577b Troy WideWord Processor Project
 *
 *
 * @reminder December 1, 2007
 * Remember to remove wrbyteen and ctrl_ppp from the inputs to
 * the ALU and its testbench
 
 */
 
/**
 * Reference:
 * Nestoras Tzartzanis, EE 577B Verilog Example, Jan 25, 1996
 * http://www-scf.usc.edu/~ee577/tutorial/verilog/alu.v
 */

/**
 * Note that all instructions are 32-bits, and that Big-Endian
 * byte and bit labeling is used. Hence, a[0] is the most
 * significant bit, and a[31] is the least significant bit.
 *
 * Use of casex and casez may affect functionality, and produce
 * larger and slower designs that omit the full_case directive
 *
 * Reference:
 * Don Mills and Clifford E. Cummings, "RTL Coding Styles That
 * Yield Simulation and Synthesis Mismatches", SNUG 1999
 *
 * ALU is a combinational logic block without clock signals
 */

`include "control.h"

// Behavioral model for the ALU
module alu (reg_A,reg_B,ctrl_ppp,ctrl_ww,alu_op,result,wrbyteen);

	// Output signals...
	// Result from copmputing an arithmetic or logical operation
	output [0:127] result;
	/**
	 * Overflow fromn arithmetic operations are ignored; use
	 * saturating mode for arithmetic operations - cap the value
	 * at the maximum value.
	 *
	 * Also, an output signal to indicate that an overflow has
	 * occurred will not be provided
	 */
	
	
	
	
	// ===============================================================
	// Input signals
	// Input register A
	input [0:127] reg_A;
	// Input register B
	input [0:127] reg_B;
	// Clock signal
	//input clock;
	// Control signal bits - ppp
	input [0:2] ctrl_ppp;
	// Control signal bits - ww
	input [0:1] ctrl_ww;
	/**
	 * Control signal bits - determine which arithmetic or logic
	 * operation to perform
	 */
	input [0:4] alu_op;
	/**
	 * Byte-write enable signals: one for each byte of the data
	 *
	 * Asserted high when each byte of the address word needs to be
	 * updated during the write operation
	 */
	input [15:0] wrbyteen;
	/**
	 * May also include: branch_offset[n:0], is_branch
	 * Size of branch offset is specified in the Instruction Set
	 * Architecture
	 *
	 * The reset signal for the ALU is ignored
	 */
	
	
	
	
	
	
	
	
	// Defining constants: parameter [name_of_constant] = value;
	parameter max_128_bits = 128'hffffffffffffffffffffffffffffffff;
	//parameter max_128_bits = 128'hfffffffffffffffffffffffffffffffff;
	//parameter max_128_bits = 128'h00112233445566778899aabbccddeeff1;
	//parameter max_128_bits = 128'h123415678901234567890123456789012;
	
	
	
	
	
	
	
	
	// ===============================================================
	// Declare "wire" signals:
	//wire FSM_OUTPUT;
	



	
	// ===============================================================
	// Declare "reg" signals: 
	reg [0:127] result;		// Output signals

	
	
	
	// ===============================================================
	
	always @(reg_A or reg_B or ctrl_ppp or ctrl_ww or alu_op or wrbyteen)
	begin
		/**
		 * Based on the assigned arithmetic or logic instruction,
		 * carry out the appropriate function on the operands
		 */
		case(alu_op)

			/**
			 * In computer science, a logical shift is a shift operator
			 * that shifts all the bits of its operand. Unlike an
			 * arithmetic shift, a logical shift does not preserve
			 * a number's sign bit or distinguish a number's exponent
			 * from its mantissa; every bit in the operand is simply
			 * moved a given number of bit positions, and the vacant
			 * bit-positions are filled in, generally with zeros
			 * (compare with a circular shift).
			 *
			 * SRL,SLL,Srli,sra,srai...
			 */
			// ======================================================

			// ======================================================

			// SRA instruction >> mv to LSB >> bit 127
			`aluwsra:
			begin
				case(ctrl_ww)
					`w8:			// sra AND `w8
					begin
						case(reg_B[5:7])
							0:
							begin
								result[0:7]<=reg_A[0:7]>>0;
								result[8:15]<=reg_A[8:15]>>0;
								result[16:23]<=reg_A[16:23]>>0;
								result[24:31]<=reg_A[24:31]>>0;
								result[32:39]<=reg_A[32:39]>>0;
								result[40:47]<=reg_A[40:47]>>0;
								result[48:55]<=reg_A[48:55]>>0;
								result[56:63]<=reg_A[56:63]>>0;
								result[64:71]<=reg_A[64:71]>>0;
								result[72:79]<=reg_A[72:79]>>0;
								result[80:87]<=reg_A[80:87]>>0;
								result[88:95]<=reg_A[88:95]>>0;
								result[96:103]<=reg_A[96:103]>>0;
								result[104:111]<=reg_A[104:111]>>0;
								result[112:119]<=reg_A[112:119]>>0;
								result[120:127]<=reg_A[120:127]>>0;
							end
							1:
							begin
								result[0:7]<=reg_A[0:7]>>1;
								result[0]<=result[0];
								result[8:15]<=reg_A[8:15]>>1;
								result[8]<=result[8];
								result[16:23]<=reg_A[16:23]>>1;
								result[16]<=result[16];
								result[24:31]<=reg_A[24:31]>>1;
								result[24]<=result[24];
								result[32:39]<=reg_A[32:39]>>1;
								result[32]<=result[32];
								result[40:47]<=reg_A[40:47]>>1;
								result[40]<=result[40];
								result[48:55]<=reg_A[48:55]>>1;
								result[48]<=result[48];
								result[56:63]<=reg_A[56:63]>>1;
								result[56]<=result[56];
								result[64:71]<=reg_A[64:71]>>1;
								result[64]<=result[64];
								result[72:79]<=reg_A[72:79]>>1;
								result[72]<=result[72];
								result[80:87]<=reg_A[80:87]>>1;
								result[80]<=result[80];
								result[88:95]<=reg_A[88:95]>>1;
								result[88]<=result[88];
								result[96:103]<=reg_A[96:103]>>1;
								result[96]<=result[96];
								result[104:111]<=reg_A[104:111]>>1;
								result[104]<=result[104];
								result[112:119]<=reg_A[112:119]>>1;
								result[112]<=result[112];
								result[120:127]<=reg_A[120:127]>>1;
								result[120]<=result[120];
							end
							2:
							begin
								result[0:7]<=reg_A[0:7]>>2;
								result[0]<=result[0];
								result[1]<=result[0];
								result[8:15]<=reg_A[8:15]>>2;
								result[8]<=result[8];
								result[9]<=result[8];
								result[16:23]<=reg_A[16:23]>>2;
								result[16]<=result[16];
								result[17]<=result[16];
								result[24:31]<=reg_A[24:31]>>2;
								result[24]<=result[24];
								result[25]<=result[24];
								result[32:39]<=reg_A[32:39]>>2;
								result[32]<=result[32];
								result[33]<=result[32];
								result[40:47]<=reg_A[40:47]>>2;
								result[40]<=result[40];
								result[41]<=result[40];
								result[48:55]<=reg_A[48:55]>>2;
								result[48]<=result[48];
								result[49]<=result[48];
								result[56:63]<=reg_A[56:63]>>2;
								result[56]<=result[56];
								result[57]<=result[56];
								result[64:71]<=reg_A[64:71]>>2;
								result[64]<=result[64];
								result[65]<=result[64];
								result[72:79]<=reg_A[72:79]>>2;
								result[72]<=result[72];
								result[73]<=result[72];
								result[80:87]<=reg_A[80:87]>>2;
								result[80]<=result[80];
								result[81]<=result[80];
								result[88:95]<=reg_A[88:95]>>2;
								result[88]<=result[88];
								result[89]<=result[88];
								result[96:103]<=reg_A[96:103]>>2;
								result[96]<=result[96];
								result[97]<=result[96];
								result[104:111]<=reg_A[104:111]>>2;
								result[104]<=result[104];
								result[105]<=result[104];
								result[112:119]<=reg_A[112:119]>>2;
								result[112]<=result[112];
								result[113]<=result[112];
								result[120:127]<=reg_A[120:127]>>2;
								result[120]<=result[120];
								result[121]<=result[120];
							end
							3:
							begin
								result[0:7]<=reg_A[0:7]>>3;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[8:15]<=reg_A[8:15]>>3;
								result[8]<=result[8];
								result[9]<=result[8];
								result[10]<=result[8];
								result[16:23]<=reg_A[16:23]>>3;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[24:31]<=reg_A[24:31]>>3;
								result[24]<=result[24];
								result[25]<=result[24];
								result[26]<=result[24];
								result[32:39]<=reg_A[32:39]>>3;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[40:47]<=reg_A[40:47]>>3;
								result[40]<=result[40];
								result[41]<=result[40];
								result[42]<=result[40];
								result[48:55]<=reg_A[48:55]>>3;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[56:63]<=reg_A[56:63]>>3;
								result[56]<=result[56];
								result[57]<=result[56];
								result[58]<=result[56];
								result[64:71]<=reg_A[64:71]>>3;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[72:79]<=reg_A[72:79]>>3;
								result[72]<=result[72];
								result[73]<=result[72];
								result[74]<=result[72];
								result[80:87]<=reg_A[80:87]>>3;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[88:95]<=reg_A[88:95]>>3;
								result[88]<=result[88];
								result[89]<=result[88];
								result[90]<=result[88];
								result[96:103]<=reg_A[96:103]>>3;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[104:111]<=reg_A[104:111]>>3;
								result[104]<=result[104];
								result[105]<=result[104];
								result[106]<=result[104];
								result[112:119]<=reg_A[112:119]>>3;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[120:127]<=reg_A[120:127]>>3;
								result[120]<=result[120];
								result[121]<=result[120];
								result[122]<=result[120];
							end
							4:
							begin
$display("entered 8 - shift 4");
								result[0:7]<=reg_A[0:7]>>4;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[8:15]<=reg_A[8:15]>>4;
								result[8]<=result[8];
								result[9]<=result[8];
								result[10]<=result[8];
								result[11]<=result[8];
								result[16:23]<=reg_A[16:23]>>4;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[24:31]<=reg_A[24:31]>>4;
								result[24]<=result[24];
								result[25]<=result[24];
								result[26]<=result[24];
								result[27]<=result[24];
								result[32:39]<=reg_A[32:39]>>4;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[40:47]<=reg_A[40:47]>>4;
								result[40]<=result[40];
								result[41]<=result[40];
								result[42]<=result[40];
								result[43]<=result[40];
								result[48:55]<=reg_A[48:55]>>4;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[56:63]<=reg_A[56:63]>>4;
								result[56]<=result[56];
								result[57]<=result[56];
								result[58]<=result[56];
								result[59]<=result[56];
								result[64:71]<=reg_A[64:71]>>4;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[72:79]<=reg_A[72:79]>>4;
								result[72]<=result[72];
								result[73]<=result[72];
								result[74]<=result[72];
								result[75]<=result[72];
								result[80:87]<=reg_A[80:87]>>4;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[88:95]<=reg_A[88:95]>>4;
								result[88]<=result[88];
								result[89]<=result[88];
								result[90]<=result[88];
								result[91]<=result[88];
								result[96:103]<=reg_A[96:103]>>4;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[104:111]<=reg_A[104:111]>>4;
								result[104]<=result[104];
								result[105]<=result[104];
								result[106]<=result[104];
								result[107]<=result[104];
								result[112:119]<=reg_A[112:119]>>4;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[120:127]<=reg_A[120:127]>>4;
								result[120]<=result[120];
								result[121]<=result[120];
								result[122]<=result[120];
								result[123]<=result[120];
							end
							5:
							begin
								result[0:7]<=reg_A[0:7]>>5;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[8:15]<=reg_A[8:15]>>5;
								result[8]<=result[8];
								result[9]<=result[8];
								result[10]<=result[8];
								result[11]<=result[8];
								result[12]<=result[8];
								result[16:23]<=reg_A[16:23]>>5;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[24:31]<=reg_A[24:31]>>5;
								result[24]<=result[24];
								result[25]<=result[24];
								result[26]<=result[24];
								result[27]<=result[24];
								result[28]<=result[24];
								result[32:39]<=reg_A[32:39]>>5;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[40:47]<=reg_A[40:47]>>5;
								result[40]<=result[40];
								result[41]<=result[40];
								result[42]<=result[40];
								result[43]<=result[40];
								result[44]<=result[40];
								result[48:55]<=reg_A[48:55]>>5;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[56:63]<=reg_A[56:63]>>5;
								result[56]<=result[56];
								result[57]<=result[56];
								result[58]<=result[56];
								result[59]<=result[56];
								result[60]<=result[56];
								result[64:71]<=reg_A[64:71]>>5;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[72:79]<=reg_A[72:79]>>5;
								result[72]<=result[72];
								result[73]<=result[72];
								result[74]<=result[72];
								result[75]<=result[72];
								result[76]<=result[72];
								result[80:87]<=reg_A[80:87]>>5;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[88:95]<=reg_A[88:95]>>5;
								result[88]<=result[88];
								result[89]<=result[88];
								result[90]<=result[88];
								result[91]<=result[88];
								result[92]<=result[88];
								result[96:103]<=reg_A[96:103]>>5;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[104:111]<=reg_A[104:111]>>5;
								result[104]<=result[104];
								result[105]<=result[104];
								result[106]<=result[104];
								result[107]<=result[104];
								result[108]<=result[104];
								result[112:119]<=reg_A[112:119]>>5;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[120:127]<=reg_A[120:127]>>5;
								result[120]<=result[120];
								result[121]<=result[120];
								result[122]<=result[120];
								result[123]<=result[120];
								result[124]<=result[120];
							end
							6:
							begin
								result[0:7]<=reg_A[0:7]>>6;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[8:15]<=reg_A[8:15]>>6;
								result[8]<=result[8];
								result[9]<=result[8];
								result[10]<=result[8];
								result[11]<=result[8];
								result[12]<=result[8];
								result[13]<=result[8];
								result[16:23]<=reg_A[16:23]>>6;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[24:31]<=reg_A[24:31]>>6;
								result[24]<=result[24];
								result[25]<=result[24];
								result[26]<=result[24];
								result[27]<=result[24];
								result[28]<=result[24];
								result[29]<=result[24];
								result[32:39]<=reg_A[32:39]>>6;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[40:47]<=reg_A[40:47]>>6;
								result[40]<=result[40];
								result[41]<=result[40];
								result[42]<=result[40];
								result[43]<=result[40];
								result[44]<=result[40];
								result[45]<=result[40];
								result[48:55]<=reg_A[48:55]>>6;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[56:63]<=reg_A[56:63]>>6;
								result[56]<=result[56];
								result[57]<=result[56];
								result[58]<=result[56];
								result[59]<=result[56];
								result[60]<=result[56];
								result[61]<=result[56];
								result[64:71]<=reg_A[64:71]>>6;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[72:79]<=reg_A[72:79]>>6;
								result[72]<=result[72];
								result[73]<=result[72];
								result[74]<=result[72];
								result[75]<=result[72];
								result[76]<=result[72];
								result[77]<=result[72];
								result[80:87]<=reg_A[80:87]>>6;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[88:95]<=reg_A[88:95]>>6;
								result[88]<=result[88];
								result[89]<=result[88];
								result[90]<=result[88];
								result[91]<=result[88];
								result[92]<=result[88];
								result[93]<=result[88];
								result[96:103]<=reg_A[96:103]>>6;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[104:111]<=reg_A[104:111]>>6;
								result[104]<=result[104];
								result[105]<=result[104];
								result[106]<=result[104];
								result[107]<=result[104];
								result[108]<=result[104];
								result[109]<=result[104];
								result[112:119]<=reg_A[112:119]>>6;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[120:127]<=reg_A[120:127]>>6;
								result[120]<=result[120];
								result[121]<=result[120];
								result[122]<=result[120];
								result[123]<=result[120];
								result[124]<=result[120];
								result[125]<=result[120];
							end
							default:		//	sra AND `w8 && 7
							begin
								result[0:7]<=reg_A[0:7]>>7;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[8:15]<=reg_A[8:15]>>7;
								result[8]<=result[8];
								result[9]<=result[8];
								result[10]<=result[8];
								result[11]<=result[8];
								result[12]<=result[8];
								result[13]<=result[8];
								result[14]<=result[8];
								result[16:23]<=reg_A[16:23]>>7;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[24:31]<=reg_A[24:31]>>7;
								result[24]<=result[24];
								result[25]<=result[24];
								result[26]<=result[24];
								result[27]<=result[24];
								result[28]<=result[24];
								result[29]<=result[24];
								result[30]<=result[24];
								result[32:39]<=reg_A[32:39]>>7;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[40:47]<=reg_A[40:47]>>7;
								result[40]<=result[40];
								result[41]<=result[40];
								result[42]<=result[40];
								result[43]<=result[40];
								result[44]<=result[40];
								result[45]<=result[40];
								result[46]<=result[40];
								result[48:55]<=reg_A[48:55]>>7;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[56:63]<=reg_A[56:63]>>7;
								result[56]<=result[56];
								result[57]<=result[56];
								result[58]<=result[56];
								result[59]<=result[56];
								result[60]<=result[56];
								result[61]<=result[56];
								result[62]<=result[56];
								result[64:71]<=reg_A[64:71]>>7;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[72:79]<=reg_A[72:79]>>7;
								result[72]<=result[72];
								result[73]<=result[72];
								result[74]<=result[72];
								result[75]<=result[72];
								result[76]<=result[72];
								result[77]<=result[72];
								result[78]<=result[72];
								result[80:87]<=reg_A[80:87]>>7;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[88:95]<=reg_A[88:95]>>7;
								result[88]<=result[88];
								result[89]<=result[88];
								result[90]<=result[88];
								result[91]<=result[88];
								result[92]<=result[88];
								result[93]<=result[88];
								result[94]<=result[88];
								result[96:103]<=reg_A[96:103]>>7;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[104:111]<=reg_A[104:111]>>7;
								result[104]<=result[104];
								result[105]<=result[104];
								result[106]<=result[104];
								result[107]<=result[104];
								result[108]<=result[104];
								result[109]<=result[104];
								result[110]<=result[104];
								result[112:119]<=reg_A[112:119]>>7;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[120:127]<=reg_A[120:127]>>7;
								result[120]<=result[120];
								result[121]<=result[120];
								result[122]<=result[120];
								result[123]<=result[120];
								result[124]<=result[120];
								result[125]<=result[120];
								result[126]<=result[120];
							end
						endcase
					end
					`w16:			// sra AND `w16 
					begin
						case(reg_B[4:7])
							0:
							begin
								result[0:15]<=reg_A[0:15]>>0;
								result[16:31]<=reg_A[16:31]>>0;
								result[32:47]<=reg_A[32:47]>>0;
								result[48:63]<=reg_A[48:63]>>0;
								result[64:79]<=reg_A[64:79]>>0;
								result[80:95]<=reg_A[80:95]>>0;
								result[96:111]<=reg_A[96:111]>>0;
								result[112:127]<=reg_A[112:127]>>0;
							end
							1:
							begin
								result[0:15]<=reg_A[0:15]>>1;
								result[0]<=result[0];
								result[16:31]<=reg_A[16:31]>>1;
								result[16]<=result[16];
								result[32:47]<=reg_A[32:47]>>1;
								result[32]<=result[32];
								result[48:63]<=reg_A[48:63]>>1;
								result[48]<=result[48];
								result[64:79]<=reg_A[64:79]>>1;
								result[64]<=result[64];
								result[80:95]<=reg_A[80:95]>>1;
								result[80]<=result[80];
								result[96:111]<=reg_A[96:111]>>1;
								result[96]<=result[96];
								result[112:127]<=reg_A[112:127]>>1;
								result[112]<=result[112];
							end
							2:
							begin
								result[0:15]<=reg_A[0:15]>>2;
								result[0]<=result[0];
								result[1]<=result[0];
								result[16:31]<=reg_A[16:31]>>2;
								result[16]<=result[16];
								result[17]<=result[16];
								result[32:47]<=reg_A[32:47]>>2;
								result[32]<=result[32];
								result[33]<=result[32];
								result[48:63]<=reg_A[48:63]>>2;
								result[48]<=result[48];
								result[49]<=result[48];
								result[64:79]<=reg_A[64:79]>>2;
								result[64]<=result[64];
								result[65]<=result[64];
								result[80:95]<=reg_A[80:95]>>2;
								result[80]<=result[80];
								result[81]<=result[80];
								result[96:111]<=reg_A[96:111]>>2;
								result[96]<=result[96];
								result[97]<=result[96];
								result[112:127]<=reg_A[112:127]>>2;
								result[112]<=result[112];
								result[113]<=result[112];
							end
							3:
							begin
								result[0:15]<=reg_A[0:15]>>3;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[16:31]<=reg_A[16:31]>>3;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[32:47]<=reg_A[32:47]>>3;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[48:63]<=reg_A[48:63]>>3;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[64:79]<=reg_A[64:79]>>3;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[80:95]<=reg_A[80:95]>>3;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[96:111]<=reg_A[96:111]>>3;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[112:127]<=reg_A[112:127]>>3;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
							end
							4:
							begin
$display("entered 16 - shift 4");
								result[0:15]<=reg_A[0:15]>>4;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[16:31]<=reg_A[16:31]>>4;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[32:47]<=reg_A[32:47]>>4;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[48:63]<=reg_A[48:63]>>4;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[64:79]<=reg_A[64:79]>>4;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[80:95]<=reg_A[80:95]>>4;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[96:111]<=reg_A[96:111]>>4;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[112:127]<=reg_A[112:127]>>4;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
							end
							5:
							begin
								result[0:15]<=reg_A[0:15]>>5;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[16:31]<=reg_A[16:31]>>5;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[32:47]<=reg_A[32:47]>>5;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[48:63]<=reg_A[48:63]>>5;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[64:79]<=reg_A[64:79]>>5;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[80:95]<=reg_A[80:95]>>5;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[96:111]<=reg_A[96:111]>>5;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[112:127]<=reg_A[112:127]>>5;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
							end
							6:
							begin
								result[0:15]<=reg_A[0:15]>>6;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[16:31]<=reg_A[16:31]>>6;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[32:47]<=reg_A[32:47]>>6;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[48:63]<=reg_A[48:63]>>6;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[64:79]<=reg_A[64:79]>>6;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[80:95]<=reg_A[80:95]>>6;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[96:111]<=reg_A[96:111]>>6;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[112:127]<=reg_A[112:127]>>6;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
							end
							7:
							begin
								result[0:15]<=reg_A[0:15]>>7;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[16:31]<=reg_A[16:31]>>7;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[32:47]<=reg_A[32:47]>>7;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[48:63]<=reg_A[48:63]>>7;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[64:79]<=reg_A[64:79]>>7;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[80:95]<=reg_A[80:95]>>7;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[96:111]<=reg_A[96:111]>>7;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[112:127]<=reg_A[112:127]>>7;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
							end
							8:
							begin
$display("entered 16 - shift 8");
								result[0:15]<=reg_A[0:15]>>8;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[16:31]<=reg_A[16:31]>>8;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[32:47]<=reg_A[32:47]>>8;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[48:63]<=reg_A[48:63]>>8;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[64:79]<=reg_A[64:79]>>8;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[80:95]<=reg_A[80:95]>>8;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[96:111]<=reg_A[96:111]>>8;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[112:127]<=reg_A[112:127]>>8;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
							end
							9:
							begin
								result[0:15]<=reg_A[0:15]>>9;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[16:31]<=reg_A[16:31]>>9;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[24]<=result[16];
								result[32:47]<=reg_A[32:47]>>9;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[48:63]<=reg_A[48:63]>>9;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[56]<=result[48];
								result[64:79]<=reg_A[64:79]>>9;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[80:95]<=reg_A[80:95]>>9;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[88]<=result[80];
								result[96:111]<=reg_A[96:111]>>9;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[112:127]<=reg_A[112:127]>>9;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
								result[120]<=result[112];
							end
							10:
							begin
								result[0:15]<=reg_A[0:15]>>10;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[16:31]<=reg_A[16:31]>>10;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[24]<=result[16];
								result[25]<=result[16];
								result[32:47]<=reg_A[32:47]>>10;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[48:63]<=reg_A[48:63]>>10;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[56]<=result[48];
								result[57]<=result[48];
								result[64:79]<=reg_A[64:79]>>10;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[80:95]<=reg_A[80:95]>>10;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[88]<=result[80];
								result[89]<=result[80];
								result[96:111]<=reg_A[96:111]>>10;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[112:127]<=reg_A[112:127]>>10;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
								result[120]<=result[112];
								result[121]<=result[112];
							end
							11:
							begin
								result[0:15]<=reg_A[0:15]>>11;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[16:31]<=reg_A[16:31]>>11;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[24]<=result[16];
								result[25]<=result[16];
								result[26]<=result[16];
								result[32:47]<=reg_A[32:47]>>11;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[48:63]<=reg_A[48:63]>>11;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[56]<=result[48];
								result[57]<=result[48];
								result[58]<=result[48];
								result[64:79]<=reg_A[64:79]>>11;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[80:95]<=reg_A[80:95]>>11;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[88]<=result[80];
								result[89]<=result[80];
								result[90]<=result[80];
								result[96:111]<=reg_A[96:111]>>11;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[112:127]<=reg_A[112:127]>>11;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
								result[120]<=result[112];
								result[121]<=result[112];
								result[122]<=result[112];
							end
							12:
							begin
								result[0:15]<=reg_A[0:15]>>12;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[16:31]<=reg_A[16:31]>>12;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[24]<=result[16];
								result[25]<=result[16];
								result[26]<=result[16];
								result[27]<=result[16];
								result[32:47]<=reg_A[32:47]>>12;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[48:63]<=reg_A[48:63]>>12;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[56]<=result[48];
								result[57]<=result[48];
								result[58]<=result[48];
								result[59]<=result[48];
								result[64:79]<=reg_A[64:79]>>12;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[80:95]<=reg_A[80:95]>>12;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[88]<=result[80];
								result[89]<=result[80];
								result[90]<=result[80];
								result[91]<=result[80];
								result[96:111]<=reg_A[96:111]>>12;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[112:127]<=reg_A[112:127]>>12;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
								result[120]<=result[112];
								result[121]<=result[112];
								result[122]<=result[112];
								result[123]<=result[112];
							end
							13:
							begin
								result[0:15]<=reg_A[0:15]>>13;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[16:31]<=reg_A[16:31]>>13;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[24]<=result[16];
								result[25]<=result[16];
								result[26]<=result[16];
								result[27]<=result[16];
								result[28]<=result[16];
								result[32:47]<=reg_A[32:47]>>13;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[48:63]<=reg_A[48:63]>>13;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[56]<=result[48];
								result[57]<=result[48];
								result[58]<=result[48];
								result[59]<=result[48];
								result[60]<=result[48];
								result[64:79]<=reg_A[64:79]>>13;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[80:95]<=reg_A[80:95]>>13;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[88]<=result[80];
								result[89]<=result[80];
								result[90]<=result[80];
								result[91]<=result[80];
								result[92]<=result[80];
								result[96:111]<=reg_A[96:111]>>13;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[112:127]<=reg_A[112:127]>>13;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
								result[120]<=result[112];
								result[121]<=result[112];
								result[122]<=result[112];
								result[123]<=result[112];
								result[124]<=result[112];
							end
							14:
							begin
$display("entered 16 - shift 14");
								result[0:15]<=reg_A[0:15]>>14;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[16:31]<=reg_A[16:31]>>14;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[24]<=result[16];
								result[25]<=result[16];
								result[26]<=result[16];
								result[27]<=result[16];
								result[28]<=result[16];
								result[29]<=result[16];
								result[32:47]<=reg_A[32:47]>>14;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[48:63]<=reg_A[48:63]>>14;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[56]<=result[48];
								result[57]<=result[48];
								result[58]<=result[48];
								result[59]<=result[48];
								result[60]<=result[48];
								result[61]<=result[48];
								result[64:79]<=reg_A[64:79]>>14;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[80:95]<=reg_A[80:95]>>14;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[88]<=result[80];
								result[89]<=result[80];
								result[90]<=result[80];
								result[91]<=result[80];
								result[92]<=result[80];
								result[93]<=result[80];
								result[96:111]<=reg_A[96:111]>>14;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[112:127]<=reg_A[112:127]>>14;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
								result[120]<=result[112];
								result[121]<=result[112];
								result[122]<=result[112];
								result[123]<=result[112];
								result[124]<=result[112];
								result[125]<=result[112];
							end
							default:			// sra AND `w16 && 15
							begin
								result[0:15]<=reg_A[0:15]>>15;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[16:31]<=reg_A[16:31]>>15;
								result[16]<=result[16];
								result[17]<=result[16];
								result[18]<=result[16];
								result[19]<=result[16];
								result[20]<=result[16];
								result[21]<=result[16];
								result[22]<=result[16];
								result[23]<=result[16];
								result[24]<=result[16];
								result[25]<=result[16];
								result[26]<=result[16];
								result[27]<=result[16];
								result[28]<=result[16];
								result[29]<=result[16];
								result[30]<=result[16];
								result[32:47]<=reg_A[32:47]>>15;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[48:63]<=reg_A[48:63]>>15;
								result[48]<=result[48];
								result[49]<=result[48];
								result[50]<=result[48];
								result[51]<=result[48];
								result[52]<=result[48];
								result[53]<=result[48];
								result[54]<=result[48];
								result[55]<=result[48];
								result[56]<=result[48];
								result[57]<=result[48];
								result[58]<=result[48];
								result[59]<=result[48];
								result[60]<=result[48];
								result[61]<=result[48];
								result[62]<=result[48];
								result[64:79]<=reg_A[64:79]>>15;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[80:95]<=reg_A[80:95]>>15;
								result[80]<=result[80];
								result[81]<=result[80];
								result[82]<=result[80];
								result[83]<=result[80];
								result[84]<=result[80];
								result[85]<=result[80];
								result[86]<=result[80];
								result[87]<=result[80];
								result[88]<=result[80];
								result[89]<=result[80];
								result[90]<=result[80];
								result[91]<=result[80];
								result[92]<=result[80];
								result[93]<=result[80];
								result[94]<=result[80];
								result[96:111]<=reg_A[96:111]>>15;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[112:127]<=reg_A[112:127]>>15;
								result[112]<=result[112];
								result[113]<=result[112];
								result[114]<=result[112];
								result[115]<=result[112];
								result[116]<=result[112];
								result[117]<=result[112];
								result[118]<=result[112];
								result[119]<=result[112];
								result[120]<=result[112];
								result[121]<=result[112];
								result[122]<=result[112];
								result[123]<=result[112];
								result[124]<=result[112];
								result[125]<=result[112];
								result[126]<=result[112];
							end
						endcase
					end
					default:				// sra AND `w32:
					begin
						case(reg_B[5:7])
							0:
							begin
								result[0:31]<=reg_A[0:31]>>0;
								result[32:63]<=reg_A[32:63]>>0;
								result[64:95]<=reg_A[64:95]>>0;
								result[96:127]<=reg_A[96:127]>>0;
							end
							1:
							begin
								result[0:31]<=reg_A[0:31]>>1;
								result[0]<=result[0];
								result[32:63]<=reg_A[32:63]>>1;
								result[32]<=result[32];
								result[64:95]<=reg_A[64:95]>>1;
								result[64]<=result[64];
								result[96:127]<=reg_A[96:127]>>1;
								result[96]<=result[96];
							end
							2:
							begin
								result[0:31]<=reg_A[0:31]>>2;
								result[0]<=result[0];
								result[1]<=result[0];
								result[32:63]<=reg_A[32:63]>>2;
								result[32]<=result[32];
								result[33]<=result[32];
								result[64:95]<=reg_A[64:95]>>2;
								result[64]<=result[64];
								result[65]<=result[64];
								result[96:127]<=reg_A[96:127]>>2;
								result[96]<=result[96];
								result[97]<=result[96];
							end
							3:
							begin
								result[0:31]<=reg_A[0:31]>>3;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[32:63]<=reg_A[32:63]>>3;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[64:95]<=reg_A[64:95]>>3;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[96:127]<=reg_A[96:127]>>3;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
							end
							4:
							begin
								result[0:31]<=reg_A[0:31]>>4;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[32:63]<=reg_A[32:63]>>4;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[64:95]<=reg_A[64:95]>>4;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[96:127]<=reg_A[96:127]>>4;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
							end
							5:
							begin
								result[0:31]<=reg_A[0:31]>>5;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[32:63]<=reg_A[32:63]>>5;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[64:95]<=reg_A[64:95]>>5;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[96:127]<=reg_A[96:127]>>5;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
							end
							6:
							begin
								result[0:31]<=reg_A[0:31]>>6;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[32:63]<=reg_A[32:63]>>6;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[64:95]<=reg_A[64:95]>>6;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[96:127]<=reg_A[96:127]>>6;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
							end
							7:
							begin
								result[0:31]<=reg_A[0:31]>>7;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[32:63]<=reg_A[32:63]>>7;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[64:95]<=reg_A[64:95]>>7;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[96:127]<=reg_A[96:127]>>7;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
							end
							8:
							begin
$display("entered 32 - shift 8");
								result[0:31]<=reg_A[0:31]>>8;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[32:63]<=reg_A[32:63]>>8;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[64:95]<=reg_A[64:95]>>8;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[96:127]<=reg_A[96:127]>>8;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
							end
							9:
							begin
								result[0:31]<=reg_A[0:31]>>9;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[32:63]<=reg_A[32:63]>>9;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[64:95]<=reg_A[64:95]>>9;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[96:127]<=reg_A[96:127]>>9;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
							end
							10:
							begin
								result[0:31]<=reg_A[0:31]>>10;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[32:63]<=reg_A[32:63]>>10;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[64:95]<=reg_A[64:95]>>10;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[96:127]<=reg_A[96:127]>>10;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
							end
							11:
							begin
$display("entered 32 - shift 11");
								result[0:31]<=reg_A[0:31]>>11;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[32:63]<=reg_A[32:63]>>11;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[64:95]<=reg_A[64:95]>>11;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[96:127]<=reg_A[96:127]>>11;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
							end
							12:
							begin
$display("entered 32 - shift 12");
								result[0:31]<=reg_A[0:31]>>12;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[32:63]<=reg_A[32:63]>>12;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[64:95]<=reg_A[64:95]>>12;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[96:127]<=reg_A[96:127]>>12;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
							end
							13:
							begin
								result[0:31]<=reg_A[0:31]>>13;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[32:63]<=reg_A[32:63]>>13;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[64:95]<=reg_A[64:95]>>13;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[96:127]<=reg_A[96:127]>>13;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
							end
							14:
							begin
								result[0:31]<=reg_A[0:31]>>14;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[32:63]<=reg_A[32:63]>>14;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[64:95]<=reg_A[64:95]>>14;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[96:127]<=reg_A[96:127]>>14;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
							end
							15:
							begin
								result[0:31]<=reg_A[0:31]>>15;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[32:63]<=reg_A[32:63]>>15;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[64:95]<=reg_A[64:95]>>15;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[96:127]<=reg_A[96:127]>>15;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
							end
							16:
							begin
$display("entered 32 - shift 16");
								result[0:31]<=reg_A[0:31]>>16;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[32:63]<=reg_A[32:63]>>16;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[64:95]<=reg_A[64:95]>>16;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[96:127]<=reg_A[96:127]>>16;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
							end
							17:
							begin
								result[0:31]<=reg_A[0:31]>>17;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[32:63]<=reg_A[32:63]>>17;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[64:95]<=reg_A[64:95]>>17;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[96:127]<=reg_A[96:127]>>17;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
							end
							18:
							begin
								result[0:31]<=reg_A[0:31]>>18;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[32:63]<=reg_A[32:63]>>18;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[64:95]<=reg_A[64:95]>>18;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[96:127]<=reg_A[96:127]>>18;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
							end
							19:
							begin
								result[0:31]<=reg_A[0:31]>>19;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[32:63]<=reg_A[32:63]>>19;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[64:95]<=reg_A[64:95]>>19;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[96:127]<=reg_A[96:127]>>19;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
							end
							20:
							begin
								result[0:31]<=reg_A[0:31]>>20;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[32:63]<=reg_A[32:63]>>20;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[64:95]<=reg_A[64:95]>>20;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[96:127]<=reg_A[96:127]>>20;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
							end
							21:
							begin
								result[0:31]<=reg_A[0:31]>>21;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[32:63]<=reg_A[32:63]>>21;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[64:95]<=reg_A[64:95]>>21;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[96:127]<=reg_A[96:127]>>21;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
							end
							22:
							begin
								result[0:31]<=reg_A[0:31]>>22;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[32:63]<=reg_A[32:63]>>22;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[64:95]<=reg_A[64:95]>>22;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[96:127]<=reg_A[96:127]>>22;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
							end
							23:
							begin
								result[0:31]<=reg_A[0:31]>>23;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[32:63]<=reg_A[32:63]>>23;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[64:95]<=reg_A[64:95]>>23;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[96:127]<=reg_A[96:127]>>23;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
							end
							24:
							begin
								result[0:31]<=reg_A[0:31]>>24;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[32:63]<=reg_A[32:63]>>24;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[64:95]<=reg_A[64:95]>>24;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[96:127]<=reg_A[96:127]>>24;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
							end
							25:
							begin
								result[0:31]<=reg_A[0:31]>>25;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[24]<=result[0];
								result[32:63]<=reg_A[32:63]>>25;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[56]<=result[32];
								result[64:95]<=reg_A[64:95]>>25;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[88]<=result[64];
								result[96:127]<=reg_A[96:127]>>25;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
								result[120]<=result[96];
							end
							26:
							begin
								result[0:31]<=reg_A[0:31]>>26;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[24]<=result[0];
								result[25]<=result[0];
								result[32:63]<=reg_A[32:63]>>26;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[56]<=result[32];
								result[57]<=result[32];
								result[64:95]<=reg_A[64:95]>>26;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[88]<=result[64];
								result[89]<=result[64];
								result[96:127]<=reg_A[96:127]>>26;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
								result[120]<=result[96];
								result[121]<=result[96];
							end
							27:
							begin
$display("entered 32 - shift 27");
								result[0:31]<=reg_A[0:31]>>27;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[24]<=result[0];
								result[25]<=result[0];
								result[26]<=result[0];
								result[32:63]<=reg_A[32:63]>>27;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[56]<=result[32];
								result[57]<=result[32];
								result[58]<=result[32];
								result[64:95]<=reg_A[64:95]>>27;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[88]<=result[64];
								result[89]<=result[64];
								result[90]<=result[64];
								result[96:127]<=reg_A[96:127]>>27;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
								result[120]<=result[96];
								result[121]<=result[96];
								result[122]<=result[96];
							end
							28:
							begin
								result[0:31]<=reg_A[0:31]>>28;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[24]<=result[0];
								result[25]<=result[0];
								result[26]<=result[0];
								result[27]<=result[0];
								result[32:63]<=reg_A[32:63]>>28;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[56]<=result[32];
								result[57]<=result[32];
								result[58]<=result[32];
								result[59]<=result[32];
								result[64:95]<=reg_A[64:95]>>28;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[88]<=result[64];
								result[89]<=result[64];
								result[90]<=result[64];
								result[91]<=result[64];
								result[96:127]<=reg_A[96:127]>>28;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
								result[120]<=result[96];
								result[121]<=result[96];
								result[122]<=result[96];
								result[123]<=result[96];
							end
							29:
							begin
								result[0:31]<=reg_A[0:31]>>29;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[24]<=result[0];
								result[25]<=result[0];
								result[26]<=result[0];
								result[27]<=result[0];
								result[28]<=result[0];
								result[32:63]<=reg_A[32:63]>>29;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[56]<=result[32];
								result[57]<=result[32];
								result[58]<=result[32];
								result[59]<=result[32];
								result[60]<=result[32];
								result[64:95]<=reg_A[64:95]>>29;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[88]<=result[64];
								result[89]<=result[64];
								result[90]<=result[64];
								result[91]<=result[64];
								result[92]<=result[64];
								result[96:127]<=reg_A[96:127]>>29;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
								result[120]<=result[96];
								result[121]<=result[96];
								result[122]<=result[96];
								result[123]<=result[96];
								result[124]<=result[96];
							end
							30:
							begin
								result[0:31]<=reg_A[0:31]>>30;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[24]<=result[0];
								result[25]<=result[0];
								result[26]<=result[0];
								result[27]<=result[0];
								result[28]<=result[0];
								result[29]<=result[0];
								result[32:63]<=reg_A[32:63]>>30;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[56]<=result[32];
								result[57]<=result[32];
								result[58]<=result[32];
								result[59]<=result[32];
								result[60]<=result[32];
								result[61]<=result[32];
								result[64:95]<=reg_A[64:95]>>30;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[88]<=result[64];
								result[89]<=result[64];
								result[90]<=result[64];
								result[91]<=result[64];
								result[92]<=result[64];
								result[93]<=result[64];
								result[96:127]<=reg_A[96:127]>>30;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
								result[120]<=result[96];
								result[121]<=result[96];
								result[122]<=result[96];
								result[123]<=result[96];
								result[124]<=result[96];
								result[125]<=result[96];
							end
							default:			// sra AND `w32 && 31
							begin
								result[0:31]<=reg_A[0:31]>>31;
								result[0]<=result[0];
								result[1]<=result[0];
								result[2]<=result[0];
								result[3]<=result[0];
								result[4]<=result[0];
								result[5]<=result[0];
								result[6]<=result[0];
								result[7]<=result[0];
								result[8]<=result[0];
								result[9]<=result[0];
								result[10]<=result[0];
								result[11]<=result[0];
								result[12]<=result[0];
								result[13]<=result[0];
								result[14]<=result[0];
								result[15]<=result[0];
								result[16]<=result[0];
								result[17]<=result[0];
								result[18]<=result[0];
								result[19]<=result[0];
								result[20]<=result[0];
								result[21]<=result[0];
								result[22]<=result[0];
								result[23]<=result[0];
								result[24]<=result[0];
								result[25]<=result[0];
								result[26]<=result[0];
								result[27]<=result[0];
								result[28]<=result[0];
								result[29]<=result[0];
								result[30]<=result[0];
								result[32:63]<=reg_A[32:63]>>31;
								result[32]<=result[32];
								result[33]<=result[32];
								result[34]<=result[32];
								result[35]<=result[32];
								result[36]<=result[32];
								result[37]<=result[32];
								result[38]<=result[32];
								result[39]<=result[32];
								result[40]<=result[32];
								result[41]<=result[32];
								result[42]<=result[32];
								result[43]<=result[32];
								result[44]<=result[32];
								result[45]<=result[32];
								result[46]<=result[32];
								result[47]<=result[32];
								result[48]<=result[32];
								result[49]<=result[32];
								result[50]<=result[32];
								result[51]<=result[32];
								result[52]<=result[32];
								result[53]<=result[32];
								result[54]<=result[32];
								result[55]<=result[32];
								result[56]<=result[32];
								result[57]<=result[32];
								result[58]<=result[32];
								result[59]<=result[32];
								result[60]<=result[32];
								result[61]<=result[32];
								result[62]<=result[32];
								result[64:95]<=reg_A[64:95]>>31;
								result[64]<=result[64];
								result[65]<=result[64];
								result[66]<=result[64];
								result[67]<=result[64];
								result[68]<=result[64];
								result[69]<=result[64];
								result[70]<=result[64];
								result[71]<=result[64];
								result[72]<=result[64];
								result[73]<=result[64];
								result[74]<=result[64];
								result[75]<=result[64];
								result[76]<=result[64];
								result[77]<=result[64];
								result[78]<=result[64];
								result[79]<=result[64];
								result[80]<=result[64];
								result[81]<=result[64];
								result[82]<=result[64];
								result[83]<=result[64];
								result[84]<=result[64];
								result[85]<=result[64];
								result[86]<=result[64];
								result[87]<=result[64];
								result[88]<=result[64];
								result[89]<=result[64];
								result[90]<=result[64];
								result[91]<=result[64];
								result[92]<=result[64];
								result[93]<=result[64];
								result[94]<=result[64];
								result[96:127]<=reg_A[96:127]>>31;
								result[96]<=result[96];
								result[97]<=result[96];
								result[98]<=result[96];
								result[99]<=result[96];
								result[100]<=result[96];
								result[101]<=result[96];
								result[102]<=result[96];
								result[103]<=result[96];
								result[104]<=result[96];
								result[105]<=result[96];
								result[106]<=result[96];
								result[107]<=result[96];
								result[108]<=result[96];
								result[109]<=result[96];
								result[110]<=result[96];
								result[111]<=result[96];
								result[112]<=result[96];
								result[113]<=result[96];
								result[114]<=result[96];
								result[115]<=result[96];
								result[116]<=result[96];
								result[117]<=result[96];
								result[118]<=result[96];
								result[119]<=result[96];
								result[120]<=result[96];
								result[121]<=result[96];
								result[122]<=result[96];
								result[123]<=result[96];
								result[124]<=result[96];
								result[125]<=result[96];
								result[126]<=result[96];
							end
						endcase
					end
				endcase
			end


			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			

			
			
			
			// ======================================================
			
			// SLL instruction << mv to LSB << bit 127
			`aluwsll:
			begin
				case(ctrl_ww)
					`w8:	// aluwsll AND `aa AND `w8
					begin
						result[0:7]<=reg_A[0:7]<<reg_B[5:7];
						result[8:15]<=reg_A[8:15]<<reg_B[13:15];
						result[16:23]<=reg_A[16:23]<<reg_B[21:23];
						result[24:31]<=reg_A[24:31]<<reg_B[29:31];
						result[32:39]<=reg_A[32:39]<<reg_B[37:39];
						result[40:47]<=reg_A[40:47]<<reg_B[45:47];
						result[48:55]<=reg_A[48:55]<<reg_B[53:55];
						result[56:63]<=reg_A[56:63]<<reg_B[61:63];
						result[64:71]<=reg_A[64:71]<<reg_B[69:71];
						result[72:79]<=reg_A[72:79]<<reg_B[77:79];
						result[80:87]<=reg_A[80:87]<<reg_B[85:87];
						result[88:95]<=reg_A[88:95]<<reg_B[93:95];
						result[96:103]<=reg_A[96:103]<<reg_B[101:103];
						result[104:111]<=reg_A[104:111]<<reg_B[109:111];
						result[112:119]<=reg_A[112:119]<<reg_B[117:119];
						result[120:127]<=reg_A[120:127]<<reg_B[125:127];
					end
		
					`w16:	// aluwsll AND `aa AND `w16
					begin
						result[0:15]<=reg_A[0:15]<<reg_B[12:15];
						result[16:31]<=reg_A[16:31]<<reg_B[28:31];
						result[32:47]<=reg_A[32:47]<<reg_B[44:47];
						result[48:63]<=reg_A[48:63]<<reg_B[60:63];
						result[64:79]<=reg_A[64:79]<<reg_B[76:79];
						result[80:95]<=reg_A[80:95]<<reg_B[92:95];
						result[96:111]<=reg_A[96:111]<<reg_B[108:111];
						result[112:127]<=reg_A[112:127]<<reg_B[124:127];
					end
		
					`w32:	// aluwsll AND `aa AND `w32
					begin
						result[0:31]<=reg_A[0:31]<<reg_B[27:31];
						result[32:63]<=reg_A[32:63]<<reg_B[59:63];
						result[64:95]<=reg_A[64:95]<<reg_B[91:95];
						result[96:127]<=reg_A[96:127]<<reg_B[123:127];
					end
					
					default:	// aluwsll AND `aa AND Default
					begin
						result<=128'd0;
					end
				endcase
			end

			
			
			/*
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 * ======================================================
			 */
			
			// ======================================================
			
			// SRL instruction >> mv to MSB >> bit 0
			`aluwsrl:
			begin
				case(ctrl_ppp)
					`aa:	// aluwsrl AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwsrl AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]>>reg_B[5:7];
								result[8:15]<=reg_A[8:15]>>reg_B[13:15];
								result[16:23]<=reg_A[16:23]>>reg_B[21:23];
								result[24:31]<=reg_A[24:31]>>reg_B[29:31];
								result[32:39]<=reg_A[32:39]>>reg_B[37:39];
								result[40:47]<=reg_A[40:47]>>reg_B[45:47];
								result[48:55]<=reg_A[48:55]>>reg_B[53:55];
								result[56:63]<=reg_A[56:63]>>reg_B[61:63];
								result[64:71]<=reg_A[64:71]>>reg_B[69:71];
								result[72:79]<=reg_A[72:79]>>reg_B[77:79];
								result[80:87]<=reg_A[80:87]>>reg_B[85:87];
								result[88:95]<=reg_A[88:95]>>reg_B[93:95];
								result[96:103]<=reg_A[96:103]>>reg_B[101:103];
								result[104:111]<=reg_A[104:111]>>reg_B[109:111];
								result[112:119]<=reg_A[112:119]>>reg_B[117:119];
								result[120:127]<=reg_A[120:127]>>reg_B[125:127];
							end
							`w16:	// aluwsrl AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]>>reg_B[12:15];
								result[16:31]<=reg_A[16:31]>>reg_B[28:31];
								result[32:47]<=reg_A[32:47]>>reg_B[44:47];
								result[48:63]<=reg_A[48:63]>>reg_B[60:63];
								result[64:79]<=reg_A[64:79]>>reg_B[76:79];
								result[80:95]<=reg_A[80:95]>>reg_B[92:95];
								result[96:111]<=reg_A[96:111]>>reg_B[108:111];
								result[112:127]<=reg_A[112:127]>>reg_B[124:127];
							end
							`w32:	// aluwsrl AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]>>reg_B[27:31];
								result[32:63]<=reg_A[32:63]>>reg_B[59:63];
								result[64:95]<=reg_A[64:95]>>reg_B[91:95];
								result[96:127]<=reg_A[96:127]>>reg_B[123:127];
							end
							
							default:	// aluwsrl AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwsrl AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwsrl AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]>>reg_B[5:7];
								result[8:15]<=reg_A[8:15]>>reg_B[13:15];
								result[16:23]<=reg_A[16:23]>>reg_B[21:23];
								result[24:31]<=reg_A[24:31]>>reg_B[29:31];
								result[32:39]<=reg_A[32:39]>>reg_B[37:39];
								result[40:47]<=reg_A[40:47]>>reg_B[45:47];
								result[48:55]<=reg_A[48:55]>>reg_B[53:55];
								result[56:63]<=reg_A[56:63]>>reg_B[61:63];
							end
							`w16:	// aluwsrl AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]>>reg_B[12:15];
								result[16:31]<=reg_A[16:31]>>reg_B[28:31];
								result[32:47]<=reg_A[32:47]>>reg_B[44:47];
								result[48:63]<=reg_A[48:63]>>reg_B[60:63];
							end
							`w32:	// aluwsrl AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]>>reg_B[27:31];
								result[32:63]<=reg_A[32:63]>>reg_B[59:63];
							end
							
							default:
							begin
								// aluwsrl AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwsrl AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwsrl AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]>>reg_B[69:71];
								result[72:79]<=reg_A[72:79]>>reg_B[77:79];
								result[80:87]<=reg_A[80:87]>>reg_B[85:87];
								result[88:95]<=reg_A[88:95]>>reg_B[93:95];
								result[96:103]<=reg_A[96:103]>>reg_B[101:103];
								result[104:111]<=reg_A[104:111]>>reg_B[109:111];
								result[112:119]<=reg_A[112:119]>>reg_B[117:119];
								result[120:127]<=reg_A[120:127]>>reg_B[125:127];
							end
							`w16:	// aluwsrl AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]>>reg_B[76:79];
								result[80:95]<=reg_A[80:95]>>reg_B[92:95];
								result[96:111]<=reg_A[96:111]>>reg_B[108:111];
								result[112:127]<=reg_A[112:127]>>reg_B[124:127];
							end
							`w32:	// aluwsrl AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]>>reg_B[91:95];
								result[96:127]<=reg_A[96:127]>>reg_B[123:127];
							end
							
							default:
							begin
									// aluwsrl AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwsrl AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwsrl AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]>>reg_B[5:7];
								result[16:23]<=reg_A[16:23]>>reg_B[21:23];
								result[32:39]<=reg_A[32:39]>>reg_B[37:39];
								result[48:55]<=reg_A[48:55]>>reg_B[53:55];
								result[64:71]<=reg_A[64:71]>>reg_B[69:71];
								result[80:87]<=reg_A[80:87]>>reg_B[85:87];
								result[96:103]<=reg_A[96:103]>>reg_B[101:103];
								result[112:119]<=reg_A[112:119]>>reg_B[117:119];
							end
							`w16:	// aluwsrl AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]>>reg_B[12:15];
								result[32:47]<=reg_A[32:47]>>reg_B[44:47];
								result[64:79]<=reg_A[64:79]>>reg_B[76:79];
								result[96:111]<=reg_A[96:111]>>reg_B[108:111];
							end
							`w32:	// aluwsrl AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]>>reg_B[27:31];
								result[64:95]<=reg_A[64:95]>>reg_B[91:95];
							end
							
							default:
							begin
								// aluwsrl AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwsrl AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwsrl AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]>>reg_B[13:15];
								result[24:31]<=reg_A[24:31]>>reg_B[29:31];
								result[40:47]<=reg_A[40:47]>>reg_B[45:47];
								result[56:63]<=reg_A[56:63]>>reg_B[61:63];
								result[72:79]<=reg_A[72:79]>>reg_B[77:79];
								result[88:95]<=reg_A[88:95]>>reg_B[93:95];
								result[104:111]<=reg_A[104:111]>>reg_B[109:111];
								result[120:127]<=reg_A[120:127]>>reg_B[125:127];
							end
							`w16:	// aluwsrl AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]>>reg_B[28:31];
								result[48:63]<=reg_A[48:63]>>reg_B[60:63];
								result[80:95]<=reg_A[80:95]>>reg_B[92:95];
								result[112:127]<=reg_A[112:127]>>reg_B[124:127];
							end
							`w32:	// aluwsrl AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]>>reg_B[59:63];
								result[96:127]<=reg_A[96:127]>>reg_B[123:127];
							end
							
							default:
							begin
								// aluwsrl AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwsrl AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwsrl AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]>>reg_B[5:7];
							end
							`w16:	// aluwsrl AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]>>reg_B[12:15];
							end
							`w32:	// aluwsrl AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]>>reg_B[27:31];
							end
							
							default:
							begin
								// aluwsrl AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwsrl AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwsrl AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]>>reg_B[125:127];
							end
							`w16:	// aluwsrl AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]>>reg_B[124:127];
							end
							`w32:	// aluwsrl AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]>>reg_B[123:127];
							end
							
							default:
							begin
								// aluwsrl AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwsrl AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end








//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================








			// ================================================
			
			// ADD instruction
			
			`aluwadd:
			begin
				case(ctrl_ppp)
					`aa:	// aluwadd AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
								result[8:15]<=reg_A[8:15]+reg_B[8:15];
								result[16:23]<=reg_A[16:23]+reg_B[16:23];
								result[24:31]<=reg_A[24:31]+reg_B[24:31];
								result[32:39]<=reg_A[32:39]+reg_B[32:39];
								result[40:47]<=reg_A[40:47]+reg_B[40:47];
								result[48:55]<=reg_A[48:55]+reg_B[48:55];
								result[56:63]<=reg_A[56:63]+reg_B[56:63];
								result[64:71]<=reg_A[64:71]+reg_B[64:71];
								result[72:79]<=reg_A[72:79]+reg_B[72:79];
								result[80:87]<=reg_A[80:87]+reg_B[80:87];
								result[88:95]<=reg_A[88:95]+reg_B[88:95];
								result[96:103]<=reg_A[96:103]+reg_B[96:103];
								result[104:111]<=reg_A[104:111]+reg_B[104:111];
								result[112:119]<=reg_A[112:119]+reg_B[112:119];
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
								result[16:31]<=reg_A[16:31]+reg_B[16:31];
								result[32:47]<=reg_A[32:47]+reg_B[32:47];
								result[48:63]<=reg_A[48:63]+reg_B[48:63];
								result[64:79]<=reg_A[64:79]+reg_B[64:79];
								result[80:95]<=reg_A[80:95]+reg_B[80:95];
								result[96:111]<=reg_A[96:111]+reg_B[96:111];
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
								result[32:63]<=reg_A[32:63]+reg_B[32:63];
								result[64:95]<=reg_A[64:95]+reg_B[64:95];
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:	// aluwadd AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwadd AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
								result[8:15]<=reg_A[8:15]+reg_B[8:15];
								result[16:23]<=reg_A[16:23]+reg_B[16:23];
								result[24:31]<=reg_A[24:31]+reg_B[24:31];
								result[32:39]<=reg_A[32:39]+reg_B[32:39];
								result[40:47]<=reg_A[40:47]+reg_B[40:47];
								result[48:55]<=reg_A[48:55]+reg_B[48:55];
								result[56:63]<=reg_A[56:63]+reg_B[56:63];
							end
							`w16:	// aluwadd AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
								result[16:31]<=reg_A[16:31]+reg_B[16:31];
								result[32:47]<=reg_A[32:47]+reg_B[32:47];
								result[48:63]<=reg_A[48:63]+reg_B[48:63];
							end
							`w32:	// aluwadd AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
								result[32:63]<=reg_A[32:63]+reg_B[32:63];
							end
							
							default:
							begin
								// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwadd AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]+reg_B[64:71];
								result[72:79]<=reg_A[72:79]+reg_B[72:79];
								result[80:87]<=reg_A[80:87]+reg_B[80:87];
								result[88:95]<=reg_A[88:95]+reg_B[88:95];
								result[96:103]<=reg_A[96:103]+reg_B[96:103];
								result[104:111]<=reg_A[104:111]+reg_B[104:111];
								result[112:119]<=reg_A[112:119]+reg_B[112:119];
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]+reg_B[64:79];
								result[80:95]<=reg_A[80:95]+reg_B[80:95];
								result[96:111]<=reg_A[96:111]+reg_B[96:111];
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]+reg_B[64:95];
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:
							begin
									// aluwadd AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwadd AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
								result[16:23]<=reg_A[16:23]+reg_B[16:23];
								result[32:39]<=reg_A[32:39]+reg_B[32:39];
								result[48:55]<=reg_A[48:55]+reg_B[48:55];
								result[64:71]<=reg_A[64:71]+reg_B[64:71];
								result[80:87]<=reg_A[80:87]+reg_B[80:87];
								result[96:103]<=reg_A[96:103]+reg_B[96:103];
								result[112:119]<=reg_A[112:119]+reg_B[112:119];
							end
							`w16:	// aluwadd AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
								result[32:47]<=reg_A[32:47]+reg_B[32:47];
								result[64:79]<=reg_A[64:79]+reg_B[64:79];
								result[96:111]<=reg_A[96:111]+reg_B[96:111];
							end
							`w32:	// aluwadd AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
								result[64:95]<=reg_A[64:95]+reg_B[64:95];
							end
							
							default:
							begin
								// aluwadd AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwadd AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]+reg_B[8:15];
								result[24:31]<=reg_A[24:31]+reg_B[24:31];
								result[40:47]<=reg_A[40:47]+reg_B[40:47];
								result[56:63]<=reg_A[56:63]+reg_B[56:63];
								result[72:79]<=reg_A[72:79]+reg_B[72:79];
								result[88:95]<=reg_A[88:95]+reg_B[88:95];
								result[104:111]<=reg_A[104:111]+reg_B[104:111];
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]+reg_B[16:31];
								result[48:63]<=reg_A[48:63]+reg_B[48:63];
								result[80:95]<=reg_A[80:95]+reg_B[80:95];
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]+reg_B[32:63];
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwadd AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]+reg_B[0:7];
							end
							`w16:	// aluwadd AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]+reg_B[0:15];
							end
							`w32:	// aluwadd AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]+reg_B[0:31];
							end
							
							default:
							begin
								// aluwadd AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwadd AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwadd AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]+reg_B[120:127];
							end
							`w16:	// aluwadd AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]+reg_B[112:127];
							end
							`w32:	// aluwadd AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]+reg_B[96:127];
							end
							
							default:
							begin
								// aluwadd AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwadd AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			// ================================================
			
			// AND instruction
			`aluwand:
			begin
				case(ctrl_ppp)
					`aa:	// aluwand AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwand AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
								result[8:15]<=reg_A[8:15]&reg_B[8:15];
								result[16:23]<=reg_A[16:23]&reg_B[16:23];
								result[24:31]<=reg_A[24:31]&reg_B[24:31];
								result[32:39]<=reg_A[32:39]&reg_B[32:39];
								result[40:47]<=reg_A[40:47]&reg_B[40:47];
								result[48:55]<=reg_A[48:55]&reg_B[48:55];
								result[56:63]<=reg_A[56:63]&reg_B[56:63];
								result[64:71]<=reg_A[64:71]&reg_B[64:71];
								result[72:79]<=reg_A[72:79]&reg_B[72:79];
								result[80:87]<=reg_A[80:87]&reg_B[80:87];
								result[88:95]<=reg_A[88:95]&reg_B[88:95];
								result[96:103]<=reg_A[96:103]&reg_B[96:103];
								result[104:111]<=reg_A[104:111]&reg_B[104:111];
								result[112:119]<=reg_A[112:119]&reg_B[112:119];
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwand AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
								result[16:31]<=reg_A[16:31]&reg_B[16:31];
								result[32:47]<=reg_A[32:47]&reg_B[32:47];
								result[48:63]<=reg_A[48:63]&reg_B[48:63];
								result[64:79]<=reg_A[64:79]&reg_B[64:79];
								result[80:95]<=reg_A[80:95]&reg_B[80:95];
								result[96:111]<=reg_A[96:111]&reg_B[96:111];
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwand AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
								result[32:63]<=reg_A[32:63]&reg_B[32:63];
								result[64:95]<=reg_A[64:95]&reg_B[64:95];
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:	// aluwand AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwand AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwand AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
								result[8:15]<=reg_A[8:15]&reg_B[8:15];
								result[16:23]<=reg_A[16:23]&reg_B[16:23];
								result[24:31]<=reg_A[24:31]&reg_B[24:31];
								result[32:39]<=reg_A[32:39]&reg_B[32:39];
								result[40:47]<=reg_A[40:47]&reg_B[40:47];
								result[48:55]<=reg_A[48:55]&reg_B[48:55];
								result[56:63]<=reg_A[56:63]&reg_B[56:63];
							end
							`w16:	// aluwand AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
								result[16:31]<=reg_A[16:31]&reg_B[16:31];
								result[32:47]<=reg_A[32:47]&reg_B[32:47];
								result[48:63]<=reg_A[48:63]&reg_B[48:63];
							end
							`w32:	// aluwand AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
								result[32:63]<=reg_A[32:63]&reg_B[32:63];
							end
							
							default:
							begin
								// aluwand AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwand AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwand AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]&reg_B[64:71];
								result[72:79]<=reg_A[72:79]&reg_B[72:79];
								result[80:87]<=reg_A[80:87]&reg_B[80:87];
								result[88:95]<=reg_A[88:95]&reg_B[88:95];
								result[96:103]<=reg_A[96:103]&reg_B[96:103];
								result[104:111]<=reg_A[104:111]&reg_B[104:111];
								result[112:119]<=reg_A[112:119]&reg_B[112:119];
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwand AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]&reg_B[64:79];
								result[80:95]<=reg_A[80:95]&reg_B[80:95];
								result[96:111]<=reg_A[96:111]&reg_B[96:111];
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwand AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]&reg_B[64:95];
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:
							begin
									// aluwand AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwand AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwand AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
								result[16:23]<=reg_A[16:23]&reg_B[16:23];
								result[32:39]<=reg_A[32:39]&reg_B[32:39];
								result[48:55]<=reg_A[48:55]&reg_B[48:55];
								result[64:71]<=reg_A[64:71]&reg_B[64:71];
								result[80:87]<=reg_A[80:87]&reg_B[80:87];
								result[96:103]<=reg_A[96:103]&reg_B[96:103];
								result[112:119]<=reg_A[112:119]&reg_B[112:119];
							end
							`w16:	// aluwand AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
								result[32:47]<=reg_A[32:47]&reg_B[32:47];
								result[64:79]<=reg_A[64:79]&reg_B[64:79];
								result[96:111]<=reg_A[96:111]&reg_B[96:111];
							end
							`w32:	// aluwand AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
								result[64:95]<=reg_A[64:95]&reg_B[64:95];
							end
							
							default:
							begin
								// aluwand AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwand AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwand AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]&reg_B[8:15];
								result[24:31]<=reg_A[24:31]&reg_B[24:31];
								result[40:47]<=reg_A[40:47]&reg_B[40:47];
								result[56:63]<=reg_A[56:63]&reg_B[56:63];
								result[72:79]<=reg_A[72:79]&reg_B[72:79];
								result[88:95]<=reg_A[88:95]&reg_B[88:95];
								result[104:111]<=reg_A[104:111]&reg_B[104:111];
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwand AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]&reg_B[16:31];
								result[48:63]<=reg_A[48:63]&reg_B[48:63];
								result[80:95]<=reg_A[80:95]&reg_B[80:95];
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwand AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]&reg_B[32:63];
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:
							begin
								// aluwand AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwand AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwand AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]&reg_B[0:7];
							end
							`w16:	// aluwand AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]&reg_B[0:15];
							end
							`w32:	// aluwand AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]&reg_B[0:31];
							end
							
							default:
							begin
								// aluwand AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwand AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwand AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]&reg_B[120:127];
							end
							`w16:	// aluwand AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]&reg_B[112:127];
							end
							`w32:	// aluwand AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]&reg_B[96:127];
							end
							
							default:
							begin
								// aluwand AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwand AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			// ==============================================
			
			
			// ================================================
			
			// NOT instruction
			`aluwnot:
			begin
				case(ctrl_ppp)
					`aa:	// aluwnot AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwnot AND `aa AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
								result[8:15]<=~reg_A[8:15];
								result[16:23]<=~reg_A[16:23];
								result[24:31]<=~reg_A[24:31];
								result[32:39]<=~reg_A[32:39];
								result[40:47]<=~reg_A[40:47];
								result[48:55]<=~reg_A[48:55];
								result[56:63]<=~reg_A[56:63];
								result[64:71]<=~reg_A[64:71];
								result[72:79]<=~reg_A[72:79];
								result[80:87]<=~reg_A[80:87];
								result[88:95]<=~reg_A[88:95];
								result[96:103]<=~reg_A[96:103];
								result[104:111]<=~reg_A[104:111];
								result[112:119]<=~reg_A[112:119];
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwnot AND `aa AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
								result[16:31]<=~reg_A[16:31];
								result[32:47]<=~reg_A[32:47];
								result[48:63]<=~reg_A[48:63];
								result[64:79]<=~reg_A[64:79];
								result[80:95]<=~reg_A[80:95];
								result[96:111]<=~reg_A[96:111];
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwnot AND `aa AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
								result[32:63]<=~reg_A[32:63];
								result[64:95]<=~reg_A[64:95];
								result[96:127]<=~reg_A[96:127];
							end
							
							default:	// aluwnot AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwnot AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwnot AND `uu AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
								result[8:15]<=~reg_A[8:15];
								result[16:23]<=~reg_A[16:23];
								result[24:31]<=~reg_A[24:31];
								result[32:39]<=~reg_A[32:39];
								result[40:47]<=~reg_A[40:47];
								result[48:55]<=~reg_A[48:55];
								result[56:63]<=~reg_A[56:63];
							end
							`w16:	// aluwnot AND `uu AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
								result[16:31]<=~reg_A[16:31];
								result[32:47]<=~reg_A[32:47];
								result[48:63]<=~reg_A[48:63];
							end
							`w32:	// aluwnot AND `uu AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
								result[32:63]<=~reg_A[32:63];
							end
							
							default:
							begin
								// aluwnot AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwnot AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwnot AND `dd AND `w8
							begin
								result[64:71]<=~reg_A[64:71];
								result[72:79]<=~reg_A[72:79];
								result[80:87]<=~reg_A[80:87];
								result[88:95]<=~reg_A[88:95];
								result[96:103]<=~reg_A[96:103];
								result[104:111]<=~reg_A[104:111];
								result[112:119]<=~reg_A[112:119];
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwnot AND `dd AND `w16
							begin
								result[64:79]<=~reg_A[64:79];
								result[80:95]<=~reg_A[80:95];
								result[96:111]<=~reg_A[96:111];
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwnot AND `dd AND `w32
							begin
								result[64:95]<=~reg_A[64:95];
								result[96:127]<=~reg_A[96:127];
							end
							
							default:
							begin
									// aluwnot AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwnot AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwnot AND `ee AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
								result[16:23]<=~reg_A[16:23];
								result[32:39]<=~reg_A[32:39];
								result[48:55]<=~reg_A[48:55];
								result[64:71]<=~reg_A[64:71];
								result[80:87]<=~reg_A[80:87];
								result[96:103]<=~reg_A[96:103];
								result[112:119]<=~reg_A[112:119];
							end
							`w16:	// aluwnot AND `ee AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
								result[32:47]<=~reg_A[32:47];
								result[64:79]<=~reg_A[64:79];
								result[96:111]<=~reg_A[96:111];
							end
							`w32:	// aluwnot AND `ee AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
								result[64:95]<=~reg_A[64:95];
							end
							
							default:
							begin
								// aluwnot AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwnot AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwnot AND `oo AND `w8
							begin
								result[8:15]<=~reg_A[8:15];
								result[24:31]<=~reg_A[24:31];
								result[40:47]<=~reg_A[40:47];
								result[56:63]<=~reg_A[56:63];
								result[72:79]<=~reg_A[72:79];
								result[88:95]<=~reg_A[88:95];
								result[104:111]<=~reg_A[104:111];
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwnot AND `oo AND `w16
							begin
								result[16:31]<=~reg_A[16:31];
								result[48:63]<=~reg_A[48:63];
								result[80:95]<=~reg_A[80:95];
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwnot AND `oo AND `w32
							begin
								result[32:63]<=~reg_A[32:63];
								result[96:127]<=~reg_A[96:127];
							end
							
							default:
							begin
								// aluwnot AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwnot AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwnot AND `mm AND `w8
							begin
								result[0:7]<=~reg_A[0:7];
							end
							`w16:	// aluwnot AND `mm AND `w16
							begin
								result[0:15]<=~reg_A[0:15];
							end
							`w32:	// aluwnot AND `mm AND `w32
							begin
								result[0:31]<=~reg_A[0:31];
							end
							
							default:
							begin
								// aluwnot AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwnot AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwnot AND `ll AND `w8
							begin
								result[120:127]<=~reg_A[120:127];
							end
							`w16:	// aluwnot AND `ll AND `w16
							begin
								result[112:127]<=~reg_A[112:127];
							end
							`w32:	// aluwnot AND `ll AND `w32
							begin
								result[96:127]<=~reg_A[96:127];
							end
							
							default:
							begin
								// aluwnot AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwnot AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			
			
			// ================================================
			
			// OR instruction
			`aluwor:
			begin
				case(ctrl_ppp)
					`aa:	// aluwor AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwor AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
								result[8:15]<=reg_A[8:15]|reg_B[8:15];
								result[16:23]<=reg_A[16:23]|reg_B[16:23];
								result[24:31]<=reg_A[24:31]|reg_B[24:31];
								result[32:39]<=reg_A[32:39]|reg_B[32:39];
								result[40:47]<=reg_A[40:47]|reg_B[40:47];
								result[48:55]<=reg_A[48:55]|reg_B[48:55];
								result[56:63]<=reg_A[56:63]|reg_B[56:63];
								result[64:71]<=reg_A[64:71]|reg_B[64:71];
								result[72:79]<=reg_A[72:79]|reg_B[72:79];
								result[80:87]<=reg_A[80:87]|reg_B[80:87];
								result[88:95]<=reg_A[88:95]|reg_B[88:95];
								result[96:103]<=reg_A[96:103]|reg_B[96:103];
								result[104:111]<=reg_A[104:111]|reg_B[104:111];
								result[112:119]<=reg_A[112:119]|reg_B[112:119];
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwor AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
								result[16:31]<=reg_A[16:31]|reg_B[16:31];
								result[32:47]<=reg_A[32:47]|reg_B[32:47];
								result[48:63]<=reg_A[48:63]|reg_B[48:63];
								result[64:79]<=reg_A[64:79]|reg_B[64:79];
								result[80:95]<=reg_A[80:95]|reg_B[80:95];
								result[96:111]<=reg_A[96:111]|reg_B[96:111];
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwor AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
								result[32:63]<=reg_A[32:63]|reg_B[32:63];
								result[64:95]<=reg_A[64:95]|reg_B[64:95];
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:	// aluwor AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwor AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwor AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
								result[8:15]<=reg_A[8:15]|reg_B[8:15];
								result[16:23]<=reg_A[16:23]|reg_B[16:23];
								result[24:31]<=reg_A[24:31]|reg_B[24:31];
								result[32:39]<=reg_A[32:39]|reg_B[32:39];
								result[40:47]<=reg_A[40:47]|reg_B[40:47];
								result[48:55]<=reg_A[48:55]|reg_B[48:55];
								result[56:63]<=reg_A[56:63]|reg_B[56:63];
							end
							`w16:	// aluwor AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
								result[16:31]<=reg_A[16:31]|reg_B[16:31];
								result[32:47]<=reg_A[32:47]|reg_B[32:47];
								result[48:63]<=reg_A[48:63]|reg_B[48:63];
							end
							`w32:	// aluwor AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
								result[32:63]<=reg_A[32:63]|reg_B[32:63];
							end
							
							default:
							begin
								// aluwor AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwor AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwor AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]|reg_B[64:71];
								result[72:79]<=reg_A[72:79]|reg_B[72:79];
								result[80:87]<=reg_A[80:87]|reg_B[80:87];
								result[88:95]<=reg_A[88:95]|reg_B[88:95];
								result[96:103]<=reg_A[96:103]|reg_B[96:103];
								result[104:111]<=reg_A[104:111]|reg_B[104:111];
								result[112:119]<=reg_A[112:119]|reg_B[112:119];
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwor AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]|reg_B[64:79];
								result[80:95]<=reg_A[80:95]|reg_B[80:95];
								result[96:111]<=reg_A[96:111]|reg_B[96:111];
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwor AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]|reg_B[64:95];
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:
							begin
									// aluwor AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwor AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwor AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
								result[16:23]<=reg_A[16:23]|reg_B[16:23];
								result[32:39]<=reg_A[32:39]|reg_B[32:39];
								result[48:55]<=reg_A[48:55]|reg_B[48:55];
								result[64:71]<=reg_A[64:71]|reg_B[64:71];
								result[80:87]<=reg_A[80:87]|reg_B[80:87];
								result[96:103]<=reg_A[96:103]|reg_B[96:103];
								result[112:119]<=reg_A[112:119]|reg_B[112:119];
							end
							`w16:	// aluwor AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
								result[32:47]<=reg_A[32:47]|reg_B[32:47];
								result[64:79]<=reg_A[64:79]|reg_B[64:79];
								result[96:111]<=reg_A[96:111]|reg_B[96:111];
							end
							`w32:	// aluwor AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
								result[64:95]<=reg_A[64:95]|reg_B[64:95];
							end
							
							default:
							begin
								// aluwor AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwor AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwor AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]|reg_B[8:15];
								result[24:31]<=reg_A[24:31]|reg_B[24:31];
								result[40:47]<=reg_A[40:47]|reg_B[40:47];
								result[56:63]<=reg_A[56:63]|reg_B[56:63];
								result[72:79]<=reg_A[72:79]|reg_B[72:79];
								result[88:95]<=reg_A[88:95]|reg_B[88:95];
								result[104:111]<=reg_A[104:111]|reg_B[104:111];
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwor AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]|reg_B[16:31];
								result[48:63]<=reg_A[48:63]|reg_B[48:63];
								result[80:95]<=reg_A[80:95]|reg_B[80:95];
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwor AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]|reg_B[32:63];
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:
							begin
								// aluwor AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwor AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwor AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]|reg_B[0:7];
							end
							`w16:	// aluwor AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]|reg_B[0:15];
							end
							`w32:	// aluwor AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]|reg_B[0:31];
							end
							
							default:
							begin
								// aluwor AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwor AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwor AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]|reg_B[120:127];
							end
							`w16:	// aluwor AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]|reg_B[112:127];
							end
							`w32:	// aluwor AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]|reg_B[96:127];
							end
							
							default:
							begin
								// aluwor AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwor AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end
			
			
			// ========================================================
			
			// XOR instruction
			`aluwxor:
			begin
				case(ctrl_ppp)
					`aa:	// aluwxor AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwxor AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]^reg_B[0:7];
								result[8:15]<=reg_A[8:15]^reg_B[8:15];
								result[16:23]<=reg_A[16:23]^reg_B[16:23];
								result[24:31]<=reg_A[24:31]^reg_B[24:31];
								result[32:39]<=reg_A[32:39]^reg_B[32:39];
								result[40:47]<=reg_A[40:47]^reg_B[40:47];
								result[48:55]<=reg_A[48:55]^reg_B[48:55];
								result[56:63]<=reg_A[56:63]^reg_B[56:63];
								result[64:71]<=reg_A[64:71]^reg_B[64:71];
								result[72:79]<=reg_A[72:79]^reg_B[72:79];
								result[80:87]<=reg_A[80:87]^reg_B[80:87];
								result[88:95]<=reg_A[88:95]^reg_B[88:95];
								result[96:103]<=reg_A[96:103]^reg_B[96:103];
								result[104:111]<=reg_A[104:111]^reg_B[104:111];
								result[112:119]<=reg_A[112:119]^reg_B[112:119];
								result[120:127]<=reg_A[120:127]^reg_B[120:127];
							end
							`w16:	// aluwxor AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]^reg_B[0:15];
								result[16:31]<=reg_A[16:31]^reg_B[16:31];
								result[32:47]<=reg_A[32:47]^reg_B[32:47];
								result[48:63]<=reg_A[48:63]^reg_B[48:63];
								result[64:79]<=reg_A[64:79]^reg_B[64:79];
								result[80:95]<=reg_A[80:95]^reg_B[80:95];
								result[96:111]<=reg_A[96:111]^reg_B[96:111];
								result[112:127]<=reg_A[112:127]^reg_B[112:127];
							end
							`w32:	// aluwxor AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]^reg_B[0:31];
								result[32:63]<=reg_A[32:63]^reg_B[32:63];
								result[64:95]<=reg_A[64:95]^reg_B[64:95];
								result[96:127]<=reg_A[96:127]^reg_B[96:127];
							end
							
							default:	// aluwxor AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwxor AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwxor AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]^reg_B[0:7];
								result[8:15]<=reg_A[8:15]^reg_B[8:15];
								result[16:23]<=reg_A[16:23]^reg_B[16:23];
								result[24:31]<=reg_A[24:31]^reg_B[24:31];
								result[32:39]<=reg_A[32:39]^reg_B[32:39];
								result[40:47]<=reg_A[40:47]^reg_B[40:47];
								result[48:55]<=reg_A[48:55]^reg_B[48:55];
								result[56:63]<=reg_A[56:63]^reg_B[56:63];
							end
							`w16:	// aluwxor AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]^reg_B[0:15];
								result[16:31]<=reg_A[16:31]^reg_B[16:31];
								result[32:47]<=reg_A[32:47]^reg_B[32:47];
								result[48:63]<=reg_A[48:63]^reg_B[48:63];
							end
							`w32:	// aluwxor AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]^reg_B[0:31];
								result[32:63]<=reg_A[32:63]^reg_B[32:63];
							end
							
							default:
							begin
								// aluwxor AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwxor AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwxor AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]^reg_B[64:71];
								result[72:79]<=reg_A[72:79]^reg_B[72:79];
								result[80:87]<=reg_A[80:87]^reg_B[80:87];
								result[88:95]<=reg_A[88:95]^reg_B[88:95];
								result[96:103]<=reg_A[96:103]^reg_B[96:103];
								result[104:111]<=reg_A[104:111]^reg_B[104:111];
								result[112:119]<=reg_A[112:119]^reg_B[112:119];
								result[120:127]<=reg_A[120:127]^reg_B[120:127];
							end
							`w16:	// aluwxor AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]^reg_B[64:79];
								result[80:95]<=reg_A[80:95]^reg_B[80:95];
								result[96:111]<=reg_A[96:111]^reg_B[96:111];
								result[112:127]<=reg_A[112:127]^reg_B[112:127];
							end
							`w32:	// aluwxor AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]^reg_B[64:95];
								result[96:127]<=reg_A[96:127]^reg_B[96:127];
							end
							
							default:
							begin
									// aluwxor AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwxor AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwxor AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]^reg_B[0:7];
								result[16:23]<=reg_A[16:23]^reg_B[16:23];
								result[32:39]<=reg_A[32:39]^reg_B[32:39];
								result[48:55]<=reg_A[48:55]^reg_B[48:55];
								result[64:71]<=reg_A[64:71]^reg_B[64:71];
								result[80:87]<=reg_A[80:87]^reg_B[80:87];
								result[96:103]<=reg_A[96:103]^reg_B[96:103];
								result[112:119]<=reg_A[112:119]^reg_B[112:119];
							end
							`w16:	// aluwxor AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]^reg_B[0:15];
								result[32:47]<=reg_A[32:47]^reg_B[32:47];
								result[64:79]<=reg_A[64:79]^reg_B[64:79];
								result[96:111]<=reg_A[96:111]^reg_B[96:111];
							end
							`w32:	// aluwxor AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]^reg_B[0:31];
								result[64:95]<=reg_A[64:95]^reg_B[64:95];
							end
							
							default:
							begin
								// aluwxor AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwxor AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwxor AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]^reg_B[8:15];
								result[24:31]<=reg_A[24:31]^reg_B[24:31];
								result[40:47]<=reg_A[40:47]^reg_B[40:47];
								result[56:63]<=reg_A[56:63]^reg_B[56:63];
								result[72:79]<=reg_A[72:79]^reg_B[72:79];
								result[88:95]<=reg_A[88:95]^reg_B[88:95];
								result[104:111]<=reg_A[104:111]^reg_B[104:111];
								result[120:127]<=reg_A[120:127]^reg_B[120:127];
							end
							`w16:	// aluwxor AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]^reg_B[16:31];
								result[48:63]<=reg_A[48:63]^reg_B[48:63];
								result[80:95]<=reg_A[80:95]^reg_B[80:95];
								result[112:127]<=reg_A[112:127]^reg_B[112:127];
							end
							`w32:	// aluwxor AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]^reg_B[32:63];
								result[96:127]<=reg_A[96:127]^reg_B[96:127];
							end
							
							default:
							begin
								// aluwxor AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwxor AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwxor AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]^reg_B[0:7];
							end
							`w16:	// aluwxor AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]^reg_B[0:15];
							end
							`w32:	// aluwxor AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]^reg_B[0:31];
							end
							
							default:
							begin
								// aluwxor AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwxor AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwxor AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]^reg_B[120:127];
							end
							`w16:	// aluwxor AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]^reg_B[112:127];
							end
							`w32:	// aluwxor AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]^reg_B[96:127];
							end
							
							default:
							begin
								// aluwxor AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwxor AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end

			
			// ======================================================
			
			// SUB instruction
			`aluwsub:
			begin
				case(ctrl_ppp)
					`aa:	// aluwsub AND `aa
					begin
						case(ctrl_ww)
							`w8:	// aluwsub AND `aa AND `w8
							begin
								result[0:7]<=reg_A[0:7]-reg_B[0:7];
								result[8:15]<=reg_A[8:15]-reg_B[8:15];
								result[16:23]<=reg_A[16:23]-reg_B[16:23];
								result[24:31]<=reg_A[24:31]-reg_B[24:31];
								result[32:39]<=reg_A[32:39]-reg_B[32:39];
								result[40:47]<=reg_A[40:47]-reg_B[40:47];
								result[48:55]<=reg_A[48:55]-reg_B[48:55];
								result[56:63]<=reg_A[56:63]-reg_B[56:63];
								result[64:71]<=reg_A[64:71]-reg_B[64:71];
								result[72:79]<=reg_A[72:79]-reg_B[72:79];
								result[80:87]<=reg_A[80:87]-reg_B[80:87];
								result[88:95]<=reg_A[88:95]-reg_B[88:95];
								result[96:103]<=reg_A[96:103]-reg_B[96:103];
								result[104:111]<=reg_A[104:111]-reg_B[104:111];
								result[112:119]<=reg_A[112:119]-reg_B[112:119];
								result[120:127]<=reg_A[120:127]-reg_B[120:127];
							end
							`w16:	// aluwsub AND `aa AND `w16
							begin
								result[0:15]<=reg_A[0:15]-reg_B[0:15];
								result[16:31]<=reg_A[16:31]-reg_B[16:31];
								result[32:47]<=reg_A[32:47]-reg_B[32:47];
								result[48:63]<=reg_A[48:63]-reg_B[48:63];
								result[64:79]<=reg_A[64:79]-reg_B[64:79];
								result[80:95]<=reg_A[80:95]-reg_B[80:95];
								result[96:111]<=reg_A[96:111]-reg_B[96:111];
								result[112:127]<=reg_A[112:127]-reg_B[112:127];
							end
							`w32:	// aluwsub AND `aa AND `w32
							begin
								result[0:31]<=reg_A[0:31]-reg_B[0:31];
								result[32:63]<=reg_A[32:63]-reg_B[32:63];
								result[64:95]<=reg_A[64:95]-reg_B[64:95];
								result[96:127]<=reg_A[96:127]-reg_B[96:127];
							end
							
							default:	// aluwsub AND `aa AND Default
							begin
								result<=128'd0;
							end
						endcase
					
					end
					`uu:	// aluwsub AND `uu
					begin
						case(ctrl_ww)
							`w8:	// aluwsub AND `uu AND `w8
							begin
								result[0:7]<=reg_A[0:7]-reg_B[0:7];
								result[8:15]<=reg_A[8:15]-reg_B[8:15];
								result[16:23]<=reg_A[16:23]-reg_B[16:23];
								result[24:31]<=reg_A[24:31]-reg_B[24:31];
								result[32:39]<=reg_A[32:39]-reg_B[32:39];
								result[40:47]<=reg_A[40:47]-reg_B[40:47];
								result[48:55]<=reg_A[48:55]-reg_B[48:55];
								result[56:63]<=reg_A[56:63]-reg_B[56:63];
							end
							`w16:	// aluwsub AND `uu AND `w16
							begin
								result[0:15]<=reg_A[0:15]-reg_B[0:15];
								result[16:31]<=reg_A[16:31]-reg_B[16:31];
								result[32:47]<=reg_A[32:47]-reg_B[32:47];
								result[48:63]<=reg_A[48:63]-reg_B[48:63];
							end
							`w32:	// aluwsub AND `uu AND `w32
							begin
								result[0:31]<=reg_A[0:31]-reg_B[0:31];
								result[32:63]<=reg_A[32:63]-reg_B[32:63];
							end
							
							default:
							begin
								// aluwsub AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`dd:	// aluwsub AND `dd
					begin
						case(ctrl_ww)
							`w8:	// aluwsub AND `dd AND `w8
							begin
								result[64:71]<=reg_A[64:71]-reg_B[64:71];
								result[72:79]<=reg_A[72:79]-reg_B[72:79];
								result[80:87]<=reg_A[80:87]-reg_B[80:87];
								result[88:95]<=reg_A[88:95]-reg_B[88:95];
								result[96:103]<=reg_A[96:103]-reg_B[96:103];
								result[104:111]<=reg_A[104:111]-reg_B[104:111];
								result[112:119]<=reg_A[112:119]-reg_B[112:119];
								result[120:127]<=reg_A[120:127]-reg_B[120:127];
							end
							`w16:	// aluwsub AND `dd AND `w16
							begin
								result[64:79]<=reg_A[64:79]-reg_B[64:79];
								result[80:95]<=reg_A[80:95]-reg_B[80:95];
								result[96:111]<=reg_A[96:111]-reg_B[96:111];
								result[112:127]<=reg_A[112:127]-reg_B[112:127];
							end
							`w32:	// aluwsub AND `dd AND `w32
							begin
								result[64:95]<=reg_A[64:95]-reg_B[64:95];
								result[96:127]<=reg_A[96:127]-reg_B[96:127];
							end
							
							default:
							begin
									// aluwsub AND `dd AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`ee:	// aluwsub AND `ee
					begin
						case(ctrl_ww)
							`w8:	// aluwsub AND `ee AND `w8
							begin
								result[0:7]<=reg_A[0:7]-reg_B[0:7];
								result[16:23]<=reg_A[16:23]-reg_B[16:23];
								result[32:39]<=reg_A[32:39]-reg_B[32:39];
								result[48:55]<=reg_A[48:55]-reg_B[48:55];
								result[64:71]<=reg_A[64:71]-reg_B[64:71];
								result[80:87]<=reg_A[80:87]-reg_B[80:87];
								result[96:103]<=reg_A[96:103]-reg_B[96:103];
								result[112:119]<=reg_A[112:119]-reg_B[112:119];
							end
							`w16:	// aluwsub AND `ee AND `w16
							begin
								result[0:15]<=reg_A[0:15]-reg_B[0:15];
								result[32:47]<=reg_A[32:47]-reg_B[32:47];
								result[64:79]<=reg_A[64:79]-reg_B[64:79];
								result[96:111]<=reg_A[96:111]-reg_B[96:111];
							end
							`w32:	// aluwsub AND `ee AND `w32
							begin
								result[0:31]<=reg_A[0:31]-reg_B[0:31];
								result[64:95]<=reg_A[64:95]-reg_B[64:95];
							end
							
							default:
							begin
								// aluwsub AND `ee AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`oo:	// aluwsub AND `oo
					begin
						case(ctrl_ww)
							`w8:	// aluwsub AND `oo AND `w8
							begin
								result[8:15]<=reg_A[8:15]-reg_B[8:15];
								result[24:31]<=reg_A[24:31]-reg_B[24:31];
								result[40:47]<=reg_A[40:47]-reg_B[40:47];
								result[56:63]<=reg_A[56:63]-reg_B[56:63];
								result[72:79]<=reg_A[72:79]-reg_B[72:79];
								result[88:95]<=reg_A[88:95]-reg_B[88:95];
								result[104:111]<=reg_A[104:111]-reg_B[104:111];
								result[120:127]<=reg_A[120:127]-reg_B[120:127];
							end
							`w16:	// aluwsub AND `oo AND `w16
							begin
								result[16:31]<=reg_A[16:31]-reg_B[16:31];
								result[48:63]<=reg_A[48:63]-reg_B[48:63];
								result[80:95]<=reg_A[80:95]-reg_B[80:95];
								result[112:127]<=reg_A[112:127]-reg_B[112:127];
							end
							`w32:	// aluwsub AND `oo AND `w32
							begin
								result[32:63]<=reg_A[32:63]-reg_B[32:63];
								result[96:127]<=reg_A[96:127]-reg_B[96:127];
							end
							
							default:
							begin
								// aluwsub AND `oo AND Default
								result<=128'd0;
							end
						endcase
					
					end
					`mm:	// aluwsub AND `mm
					begin
						case(ctrl_ww)
							`w8:	// aluwsub AND `mm AND `w8
							begin
								result[0:7]<=reg_A[0:7]-reg_B[0:7];
							end
							`w16:	// aluwsub AND `mm AND `w16
							begin
								result[0:15]<=reg_A[0:15]-reg_B[0:15];
							end
							`w32:	// aluwsub AND `mm AND `w32
							begin
								result[0:31]<=reg_A[0:31]-reg_B[0:31];
							end
							
							default:
							begin
								// aluwsub AND `mm AND `w8
								result<=128'd0;
							end
						endcase
					
					end
					`ll:	// aluwsub AND `ll
					begin
						case(ctrl_ww)
							`w8:	// aluwsub AND `ll AND `w8
							begin
								result[120:127]<=reg_A[120:127]-reg_B[120:127];
							end
							`w16:	// aluwsub AND `ll AND `w16
							begin
								result[112:127]<=reg_A[112:127]-reg_B[112:127];
							end
							`w32:	// aluwsub AND `ll AND `w32
							begin
								result[96:127]<=reg_A[96:127]-reg_B[96:127];
							end
							
							default:
							begin
								// aluwsub AND `ll AND Default
								result<=128'd0;
							end
						endcase
					
					end
					default:	// aluwsub AND Default
					begin
						result<=128'd0;
					end
				endcase
				
			end

			

//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================
//================================================================================




			// ================================================
			
			// PRM instruction
			
			`aluwprm:
			begin
				case(ctrl_ppp)
					`aa:	// aluwprm PRM `aa
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase

						case(reg_B[12:15]) //byte1
						4'd0:
							result[8:15]<=reg_A[0:7];
						4'd1:
							result[8:15]<=reg_A[8:15];
						4'd2:
							result[8:15]<=reg_A[16:23];
						4'd3:
							result[8:15]<=reg_A[24:31];
						4'd4:
							result[8:15]<=reg_A[32:39];
						4'd5:
							result[8:15]<=reg_A[40:47];
						4'd6:
							result[8:15]<=reg_A[48:55];
						4'd7:
							result[8:15]<=reg_A[56:63];
						4'd8:
							result[8:15]<=reg_A[64:71];
						4'd9:
							result[8:15]<=reg_A[72:79];
						4'd10:
							result[8:15]<=reg_A[80:87];
						4'd11:
							result[8:15]<=reg_A[88:95];
						4'd12:
							result[8:15]<=reg_A[96:103];
						4'd13:
							result[8:15]<=reg_A[104:111];
						4'd14:
							result[8:15]<=reg_A[112:119];
						4'd15:
							result[8:15]<=reg_A[120:127];
						endcase

						case(reg_B[20:23]) //byte2
						4'd0:
							result[16:23]<=reg_A[0:7];
						4'd1:
							result[16:23]<=reg_A[8:15];
						4'd2:
							result[16:23]<=reg_A[16:23];
						4'd3:
							result[16:23]<=reg_A[24:31];
						4'd4:
							result[16:23]<=reg_A[32:39];
						4'd5:
							result[16:23]<=reg_A[40:47];
						4'd6:
							result[16:23]<=reg_A[48:55];
						4'd7:
							result[16:23]<=reg_A[56:63];
						4'd8:
							result[16:23]<=reg_A[64:71];
						4'd9:
							result[16:23]<=reg_A[72:79];
						4'd10:
							result[16:23]<=reg_A[80:87];
						4'd11:
							result[16:23]<=reg_A[88:95];
						4'd12:
							result[16:23]<=reg_A[96:103];
						4'd13:
							result[16:23]<=reg_A[104:111];
						4'd14:
							result[16:23]<=reg_A[112:119];
						4'd15:
							result[16:23]<=reg_A[120:127];
						endcase

						case(reg_B[28:31]) //byte3
						4'd0:
							result[24:31]<=reg_A[0:7];
						4'd1:
							result[24:31]<=reg_A[8:15];
						4'd2:
							result[24:31]<=reg_A[16:23];
						4'd3:
							result[24:31]<=reg_A[24:31];
						4'd4:
							result[24:31]<=reg_A[32:39];
						4'd5:
							result[24:31]<=reg_A[40:47];
						4'd6:
							result[24:31]<=reg_A[48:55];
						4'd7:
							result[24:31]<=reg_A[56:63];
						4'd8:
							result[24:31]<=reg_A[64:71];
						4'd9:
							result[24:31]<=reg_A[72:79];
						4'd10:
							result[24:31]<=reg_A[80:87];
						4'd11:
							result[24:31]<=reg_A[88:95];
						4'd12:
							result[24:31]<=reg_A[96:103];
						4'd13:
							result[24:31]<=reg_A[104:111];
						4'd14:
							result[24:31]<=reg_A[112:119];
						4'd15:
							result[24:31]<=reg_A[120:127];
						endcase

						case(reg_B[36:39]) //byte4
						4'd0:
							result[32:39]<=reg_A[0:7];
						4'd1:
							result[32:39]<=reg_A[8:15];
						4'd2:
							result[32:39]<=reg_A[16:23];
						4'd3:
							result[32:39]<=reg_A[24:31];
						4'd4:
							result[32:39]<=reg_A[32:39];
						4'd5:
							result[32:39]<=reg_A[40:47];
						4'd6:
							result[32:39]<=reg_A[48:55];
						4'd7:
							result[32:39]<=reg_A[56:63];
						4'd8:
							result[32:39]<=reg_A[64:71];
						4'd9:
							result[32:39]<=reg_A[72:79];
						4'd10:
							result[32:39]<=reg_A[80:87];
						4'd11:
							result[32:39]<=reg_A[88:95];
						4'd12:
							result[32:39]<=reg_A[96:103];
						4'd13:
							result[32:39]<=reg_A[104:111];
						4'd14:
							result[32:39]<=reg_A[112:119];
						4'd15:
							result[32:39]<=reg_A[120:127];
						endcase

						case(reg_B[44:47]) //byte5
						4'd0:
							result[40:47]<=reg_A[0:7];
						4'd1:
							result[40:47]<=reg_A[8:15];
						4'd2:
							result[40:47]<=reg_A[16:23];
						4'd3:
							result[40:47]<=reg_A[24:31];
						4'd4:
							result[40:47]<=reg_A[32:39];
						4'd5:
							result[40:47]<=reg_A[40:47];
						4'd6:
							result[40:47]<=reg_A[48:55];
						4'd7:
							result[40:47]<=reg_A[56:63];
						4'd8:
							result[40:47]<=reg_A[64:71];
						4'd9:
							result[40:47]<=reg_A[72:79];
						4'd10:
							result[40:47]<=reg_A[80:87];
						4'd11:
							result[40:47]<=reg_A[88:95];
						4'd12:
							result[40:47]<=reg_A[96:103];
						4'd13:
							result[40:47]<=reg_A[104:111];
						4'd14:
							result[40:47]<=reg_A[112:119];
						4'd15:
							result[40:47]<=reg_A[120:127];
						endcase

						case(reg_B[52:55]) //byte6
						4'd0:
							result[48:55]<=reg_A[0:7];
						4'd1:
							result[48:55]<=reg_A[8:15];
						4'd2:
							result[48:55]<=reg_A[16:23];
						4'd3:
							result[48:55]<=reg_A[24:31];
						4'd4:
							result[48:55]<=reg_A[32:39];
						4'd5:
							result[48:55]<=reg_A[40:47];
						4'd6:
							result[48:55]<=reg_A[48:55];
						4'd7:
							result[48:55]<=reg_A[56:63];
						4'd8:
							result[48:55]<=reg_A[64:71];
						4'd9:
							result[48:55]<=reg_A[72:79];
						4'd10:
							result[48:55]<=reg_A[80:87];
						4'd11:
							result[48:55]<=reg_A[88:95];
						4'd12:
							result[48:55]<=reg_A[96:103];
						4'd13:
							result[48:55]<=reg_A[104:111];
						4'd14:
							result[48:55]<=reg_A[112:119];
						4'd15:
							result[48:55]<=reg_A[120:127];
						endcase

						case(reg_B[60:63]) //byte7
						4'd0:
							result[56:63]<=reg_A[0:7];
						4'd1:
							result[56:63]<=reg_A[8:15];
						4'd2:
							result[56:63]<=reg_A[16:23];
						4'd3:
							result[56:63]<=reg_A[24:31];
						4'd4:
							result[56:63]<=reg_A[32:39];
						4'd5:
							result[56:63]<=reg_A[40:47];
						4'd6:
							result[56:63]<=reg_A[48:55];
						4'd7:
							result[56:63]<=reg_A[56:63];
						4'd8:
							result[56:63]<=reg_A[64:71];
						4'd9:
							result[56:63]<=reg_A[72:79];
						4'd10:
							result[56:63]<=reg_A[80:87];
						4'd11:
							result[56:63]<=reg_A[88:95];
						4'd12:
							result[56:63]<=reg_A[96:103];
						4'd13:
							result[56:63]<=reg_A[104:111];
						4'd14:
							result[56:63]<=reg_A[112:119];
						4'd15:
							result[56:63]<=reg_A[120:127];
						endcase

						case(reg_B[68:71]) //byte8
						4'd0:
							result[64:71]<=reg_A[0:7];
						4'd1:
							result[64:71]<=reg_A[8:15];
						4'd2:
							result[64:71]<=reg_A[16:23];
						4'd3:
							result[64:71]<=reg_A[24:31];
						4'd4:
							result[64:71]<=reg_A[32:39];
						4'd5:
							result[64:71]<=reg_A[40:47];
						4'd6:
							result[64:71]<=reg_A[48:55];
						4'd7:
							result[64:71]<=reg_A[56:63];
						4'd8:
							result[64:71]<=reg_A[64:71];
						4'd9:
							result[64:71]<=reg_A[72:79];
						4'd10:
							result[64:71]<=reg_A[80:87];
						4'd11:
							result[64:71]<=reg_A[88:95];
						4'd12:
							result[64:71]<=reg_A[96:103];
						4'd13:
							result[64:71]<=reg_A[104:111];
						4'd14:
							result[64:71]<=reg_A[112:119];
						4'd15:
							result[64:71]<=reg_A[120:127];
						endcase

						case(reg_B[76:79]) //byte9
						4'd0:
							result[72:79]<=reg_A[0:7];
						4'd1:
							result[72:79]<=reg_A[8:15];
						4'd2:
							result[72:79]<=reg_A[16:23];
						4'd3:
							result[72:79]<=reg_A[24:31];
						4'd4:
							result[72:79]<=reg_A[32:39];
						4'd5:
							result[72:79]<=reg_A[40:47];
						4'd6:
							result[72:79]<=reg_A[48:55];
						4'd7:
							result[72:79]<=reg_A[56:63];
						4'd8:
							result[72:79]<=reg_A[64:71];
						4'd9:
							result[72:79]<=reg_A[72:79];
						4'd10:
							result[72:79]<=reg_A[80:87];
						4'd11:
							result[72:79]<=reg_A[88:95];
						4'd12:
							result[72:79]<=reg_A[96:103];
						4'd13:
							result[72:79]<=reg_A[104:111];
						4'd14:
							result[72:79]<=reg_A[112:119];
						4'd15:
							result[72:79]<=reg_A[120:127];
						endcase

						case(reg_B[84:87]) //byte10
						4'd0:
							result[80:87]<=reg_A[0:7];
						4'd1:
							result[80:87]<=reg_A[8:15];
						4'd2:
							result[80:87]<=reg_A[16:23];
						4'd3:
							result[80:87]<=reg_A[24:31];
						4'd4:
							result[80:87]<=reg_A[32:39];
						4'd5:
							result[80:87]<=reg_A[40:47];
						4'd6:
							result[80:87]<=reg_A[48:55];
						4'd7:
							result[80:87]<=reg_A[56:63];
						4'd8:
							result[80:87]<=reg_A[64:71];
						4'd9:
							result[80:87]<=reg_A[72:79];
						4'd10:
							result[80:87]<=reg_A[80:87];
						4'd11:
							result[80:87]<=reg_A[88:95];
						4'd12:
							result[80:87]<=reg_A[96:103];
						4'd13:
							result[80:87]<=reg_A[104:111];
						4'd14:
							result[80:87]<=reg_A[112:119];
						4'd15:
							result[80:87]<=reg_A[120:127];
						endcase

						case(reg_B[92:95]) //byte11
						4'd0:
							result[88:95]<=reg_A[0:7];
						4'd1:
							result[88:95]<=reg_A[8:15];
						4'd2:
							result[88:95]<=reg_A[16:23];
						4'd3:
							result[88:95]<=reg_A[24:31];
						4'd4:
							result[88:95]<=reg_A[32:39];
						4'd5:
							result[88:95]<=reg_A[40:47];
						4'd6:
							result[88:95]<=reg_A[48:55];
						4'd7:
							result[88:95]<=reg_A[56:63];
						4'd8:
							result[88:95]<=reg_A[64:71];
						4'd9:
							result[88:95]<=reg_A[72:79];
						4'd10:
							result[88:95]<=reg_A[80:87];
						4'd11:
							result[88:95]<=reg_A[88:95];
						4'd12:
							result[88:95]<=reg_A[96:103];
						4'd13:
							result[88:95]<=reg_A[104:111];
						4'd14:
							result[88:95]<=reg_A[112:119];
						4'd15:
							result[88:95]<=reg_A[120:127];
						endcase

						case(reg_B[100:103]) //byte12
						4'd0:
							result[96:103]<=reg_A[0:7];
						4'd1:
							result[96:103]<=reg_A[8:15];
						4'd2:
							result[96:103]<=reg_A[16:23];
						4'd3:
							result[96:103]<=reg_A[24:31];
						4'd4:
							result[96:103]<=reg_A[32:39];
						4'd5:
							result[96:103]<=reg_A[40:47];
						4'd6:
							result[96:103]<=reg_A[48:55];
						4'd7:
							result[96:103]<=reg_A[56:63];
						4'd8:
							result[96:103]<=reg_A[64:71];
						4'd9:
							result[96:103]<=reg_A[72:79];
						4'd10:
							result[96:103]<=reg_A[80:87];
						4'd11:
							result[96:103]<=reg_A[88:95];
						4'd12:
							result[96:103]<=reg_A[96:103];
						4'd13:
							result[96:103]<=reg_A[104:111];
						4'd14:
							result[96:103]<=reg_A[112:119];
						4'd15:
							result[96:103]<=reg_A[120:127];
						endcase

						case(reg_B[108:111]) //byte13
						4'd0:
							result[104:111]<=reg_A[0:7];
						4'd1:
							result[104:111]<=reg_A[8:15];
						4'd2:
							result[104:111]<=reg_A[16:23];
						4'd3:
							result[104:111]<=reg_A[24:31];
						4'd4:
							result[104:111]<=reg_A[32:39];
						4'd5:
							result[104:111]<=reg_A[40:47];
						4'd6:
							result[104:111]<=reg_A[48:55];
						4'd7:
							result[104:111]<=reg_A[56:63];
						4'd8:
							result[104:111]<=reg_A[64:71];
						4'd9:
							result[104:111]<=reg_A[72:79];
						4'd10:
							result[104:111]<=reg_A[80:87];
						4'd11:
							result[104:111]<=reg_A[88:95];
						4'd12:
							result[104:111]<=reg_A[96:103];
						4'd13:
							result[104:111]<=reg_A[104:111];
						4'd14:
							result[104:111]<=reg_A[112:119];
						4'd15:
							result[104:111]<=reg_A[120:127];
						endcase

						case(reg_B[116:119]) //byte14
						4'd0:
							result[112:119]<=reg_A[112:119];
						4'd1:
							result[112:119]<=reg_A[8:15];
						4'd2:
							result[112:119]<=reg_A[16:23];
						4'd3:
							result[112:119]<=reg_A[24:31];
						4'd4:
							result[112:119]<=reg_A[32:39];
						4'd5:
							result[112:119]<=reg_A[40:47];
						4'd6:
							result[112:119]<=reg_A[48:55];
						4'd7:
							result[112:119]<=reg_A[56:63];
						4'd8:
							result[112:119]<=reg_A[64:71];
						4'd9:
							result[112:119]<=reg_A[72:79];
						4'd10:
							result[112:119]<=reg_A[80:87];
						4'd11:
							result[112:119]<=reg_A[88:95];
						4'd12:
							result[112:119]<=reg_A[96:103];
						4'd13:
							result[112:119]<=reg_A[104:111];
						4'd14:
							result[112:119]<=reg_A[112:119];
						4'd15:
							result[112:119]<=reg_A[120:127];
						endcase

						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					`uu:	// aluwprm PRM `uu
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase

						case(reg_B[12:15]) //byte1
						4'd0:
							result[8:15]<=reg_A[0:7];
						4'd1:
							result[8:15]<=reg_A[8:15];
						4'd2:
							result[8:15]<=reg_A[16:23];
						4'd3:
							result[8:15]<=reg_A[24:31];
						4'd4:
							result[8:15]<=reg_A[32:39];
						4'd5:
							result[8:15]<=reg_A[40:47];
						4'd6:
							result[8:15]<=reg_A[48:55];
						4'd7:
							result[8:15]<=reg_A[56:63];
						4'd8:
							result[8:15]<=reg_A[64:71];
						4'd9:
							result[8:15]<=reg_A[72:79];
						4'd10:
							result[8:15]<=reg_A[80:87];
						4'd11:
							result[8:15]<=reg_A[88:95];
						4'd12:
							result[8:15]<=reg_A[96:103];
						4'd13:
							result[8:15]<=reg_A[104:111];
						4'd14:
							result[8:15]<=reg_A[112:119];
						4'd15:
							result[8:15]<=reg_A[120:127];
						endcase

						case(reg_B[20:23]) //byte2
						4'd0:
							result[16:23]<=reg_A[0:7];
						4'd1:
							result[16:23]<=reg_A[8:15];
						4'd2:
							result[16:23]<=reg_A[16:23];
						4'd3:
							result[16:23]<=reg_A[24:31];
						4'd4:
							result[16:23]<=reg_A[32:39];
						4'd5:
							result[16:23]<=reg_A[40:47];
						4'd6:
							result[16:23]<=reg_A[48:55];
						4'd7:
							result[16:23]<=reg_A[56:63];
						4'd8:
							result[16:23]<=reg_A[64:71];
						4'd9:
							result[16:23]<=reg_A[72:79];
						4'd10:
							result[16:23]<=reg_A[80:87];
						4'd11:
							result[16:23]<=reg_A[88:95];
						4'd12:
							result[16:23]<=reg_A[96:103];
						4'd13:
							result[16:23]<=reg_A[104:111];
						4'd14:
							result[16:23]<=reg_A[112:119];
						4'd15:
							result[16:23]<=reg_A[120:127];
						endcase

						case(reg_B[28:31]) //byte3
						4'd0:
							result[24:31]<=reg_A[0:7];
						4'd1:
							result[24:31]<=reg_A[8:15];
						4'd2:
							result[24:31]<=reg_A[16:23];
						4'd3:
							result[24:31]<=reg_A[24:31];
						4'd4:
							result[24:31]<=reg_A[32:39];
						4'd5:
							result[24:31]<=reg_A[40:47];
						4'd6:
							result[24:31]<=reg_A[48:55];
						4'd7:
							result[24:31]<=reg_A[56:63];
						4'd8:
							result[24:31]<=reg_A[64:71];
						4'd9:
							result[24:31]<=reg_A[72:79];
						4'd10:
							result[24:31]<=reg_A[80:87];
						4'd11:
							result[24:31]<=reg_A[88:95];
						4'd12:
							result[24:31]<=reg_A[96:103];
						4'd13:
							result[24:31]<=reg_A[104:111];
						4'd14:
							result[24:31]<=reg_A[112:119];
						4'd15:
							result[24:31]<=reg_A[120:127];
						endcase

						case(reg_B[36:39]) //byte4
						4'd0:
							result[32:39]<=reg_A[0:7];
						4'd1:
							result[32:39]<=reg_A[8:15];
						4'd2:
							result[32:39]<=reg_A[16:23];
						4'd3:
							result[32:39]<=reg_A[24:31];
						4'd4:
							result[32:39]<=reg_A[32:39];
						4'd5:
							result[32:39]<=reg_A[40:47];
						4'd6:
							result[32:39]<=reg_A[48:55];
						4'd7:
							result[32:39]<=reg_A[56:63];
						4'd8:
							result[32:39]<=reg_A[64:71];
						4'd9:
							result[32:39]<=reg_A[72:79];
						4'd10:
							result[32:39]<=reg_A[80:87];
						4'd11:
							result[32:39]<=reg_A[88:95];
						4'd12:
							result[32:39]<=reg_A[96:103];
						4'd13:
							result[32:39]<=reg_A[104:111];
						4'd14:
							result[32:39]<=reg_A[112:119];
						4'd15:
							result[32:39]<=reg_A[120:127];
						endcase

						case(reg_B[44:47]) //byte5
						4'd0:
							result[40:47]<=reg_A[0:7];
						4'd1:
							result[40:47]<=reg_A[8:15];
						4'd2:
							result[40:47]<=reg_A[16:23];
						4'd3:
							result[40:47]<=reg_A[24:31];
						4'd4:
							result[40:47]<=reg_A[32:39];
						4'd5:
							result[40:47]<=reg_A[40:47];
						4'd6:
							result[40:47]<=reg_A[48:55];
						4'd7:
							result[40:47]<=reg_A[56:63];
						4'd8:
							result[40:47]<=reg_A[64:71];
						4'd9:
							result[40:47]<=reg_A[72:79];
						4'd10:
							result[40:47]<=reg_A[80:87];
						4'd11:
							result[40:47]<=reg_A[88:95];
						4'd12:
							result[40:47]<=reg_A[96:103];
						4'd13:
							result[40:47]<=reg_A[104:111];
						4'd14:
							result[40:47]<=reg_A[112:119];
						4'd15:
							result[40:47]<=reg_A[120:127];
						endcase

						case(reg_B[52:55]) //byte6
						4'd0:
							result[48:55]<=reg_A[0:7];
						4'd1:
							result[48:55]<=reg_A[8:15];
						4'd2:
							result[48:55]<=reg_A[16:23];
						4'd3:
							result[48:55]<=reg_A[24:31];
						4'd4:
							result[48:55]<=reg_A[32:39];
						4'd5:
							result[48:55]<=reg_A[40:47];
						4'd6:
							result[48:55]<=reg_A[48:55];
						4'd7:
							result[48:55]<=reg_A[56:63];
						4'd8:
							result[48:55]<=reg_A[64:71];
						4'd9:
							result[48:55]<=reg_A[72:79];
						4'd10:
							result[48:55]<=reg_A[80:87];
						4'd11:
							result[48:55]<=reg_A[88:95];
						4'd12:
							result[48:55]<=reg_A[96:103];
						4'd13:
							result[48:55]<=reg_A[104:111];
						4'd14:
							result[48:55]<=reg_A[112:119];
						4'd15:
							result[48:55]<=reg_A[120:127];
						endcase

						case(reg_B[60:63]) //byte7
						4'd0:
							result[56:63]<=reg_A[0:7];
						4'd1:
							result[56:63]<=reg_A[8:15];
						4'd2:
							result[56:63]<=reg_A[16:23];
						4'd3:
							result[56:63]<=reg_A[24:31];
						4'd4:
							result[56:63]<=reg_A[32:39];
						4'd5:
							result[56:63]<=reg_A[40:47];
						4'd6:
							result[56:63]<=reg_A[48:55];
						4'd7:
							result[56:63]<=reg_A[56:63];
						4'd8:
							result[56:63]<=reg_A[64:71];
						4'd9:
							result[56:63]<=reg_A[72:79];
						4'd10:
							result[56:63]<=reg_A[80:87];
						4'd11:
							result[56:63]<=reg_A[88:95];
						4'd12:
							result[56:63]<=reg_A[96:103];
						4'd13:
							result[56:63]<=reg_A[104:111];
						4'd14:
							result[56:63]<=reg_A[112:119];
						4'd15:
							result[56:63]<=reg_A[120:127];
						endcase

						//bytes8-15
						result[64:127]<=64'd0;
					end
					`dd:	// aluwprm PRM `dd
					begin
						//bytes0-7
						result[0:63]<=64'd0;

						case(reg_B[68:71]) //byte8
						4'd0:
							result[64:71]<=reg_A[0:7];
						4'd1:
							result[64:71]<=reg_A[8:15];
						4'd2:
							result[64:71]<=reg_A[16:23];
						4'd3:
							result[64:71]<=reg_A[24:31];
						4'd4:
							result[64:71]<=reg_A[32:39];
						4'd5:
							result[64:71]<=reg_A[40:47];
						4'd6:
							result[64:71]<=reg_A[48:55];
						4'd7:
							result[64:71]<=reg_A[56:63];
						4'd8:
							result[64:71]<=reg_A[64:71];
						4'd9:
							result[64:71]<=reg_A[72:79];
						4'd10:
							result[64:71]<=reg_A[80:87];
						4'd11:
							result[64:71]<=reg_A[88:95];
						4'd12:
							result[64:71]<=reg_A[96:103];
						4'd13:
							result[64:71]<=reg_A[104:111];
						4'd14:
							result[64:71]<=reg_A[112:119];
						4'd15:
							result[64:71]<=reg_A[120:127];
						endcase

						case(reg_B[76:79]) //byte9
						4'd0:
							result[72:79]<=reg_A[0:7];
						4'd1:
							result[72:79]<=reg_A[8:15];
						4'd2:
							result[72:79]<=reg_A[16:23];
						4'd3:
							result[72:79]<=reg_A[24:31];
						4'd4:
							result[72:79]<=reg_A[32:39];
						4'd5:
							result[72:79]<=reg_A[40:47];
						4'd6:
							result[72:79]<=reg_A[48:55];
						4'd7:
							result[72:79]<=reg_A[56:63];
						4'd8:
							result[72:79]<=reg_A[64:71];
						4'd9:
							result[72:79]<=reg_A[72:79];
						4'd10:
							result[72:79]<=reg_A[80:87];
						4'd11:
							result[72:79]<=reg_A[88:95];
						4'd12:
							result[72:79]<=reg_A[96:103];
						4'd13:
							result[72:79]<=reg_A[104:111];
						4'd14:
							result[72:79]<=reg_A[112:119];
						4'd15:
							result[72:79]<=reg_A[120:127];
						endcase

						case(reg_B[84:87]) //byte10
						4'd0:
							result[80:87]<=reg_A[0:7];
						4'd1:
							result[80:87]<=reg_A[8:15];
						4'd2:
							result[80:87]<=reg_A[16:23];
						4'd3:
							result[80:87]<=reg_A[24:31];
						4'd4:
							result[80:87]<=reg_A[32:39];
						4'd5:
							result[80:87]<=reg_A[40:47];
						4'd6:
							result[80:87]<=reg_A[48:55];
						4'd7:
							result[80:87]<=reg_A[56:63];
						4'd8:
							result[80:87]<=reg_A[64:71];
						4'd9:
							result[80:87]<=reg_A[72:79];
						4'd10:
							result[80:87]<=reg_A[80:87];
						4'd11:
							result[80:87]<=reg_A[88:95];
						4'd12:
							result[80:87]<=reg_A[96:103];
						4'd13:
							result[80:87]<=reg_A[104:111];
						4'd14:
							result[80:87]<=reg_A[112:119];
						4'd15:
							result[80:87]<=reg_A[120:127];
						endcase

						case(reg_B[92:95]) //byte11
						4'd0:
							result[88:95]<=reg_A[0:7];
						4'd1:
							result[88:95]<=reg_A[8:15];
						4'd2:
							result[88:95]<=reg_A[16:23];
						4'd3:
							result[88:95]<=reg_A[24:31];
						4'd4:
							result[88:95]<=reg_A[32:39];
						4'd5:
							result[88:95]<=reg_A[40:47];
						4'd6:
							result[88:95]<=reg_A[48:55];
						4'd7:
							result[88:95]<=reg_A[56:63];
						4'd8:
							result[88:95]<=reg_A[64:71];
						4'd9:
							result[88:95]<=reg_A[72:79];
						4'd10:
							result[88:95]<=reg_A[80:87];
						4'd11:
							result[88:95]<=reg_A[88:95];
						4'd12:
							result[88:95]<=reg_A[96:103];
						4'd13:
							result[88:95]<=reg_A[104:111];
						4'd14:
							result[88:95]<=reg_A[112:119];
						4'd15:
							result[88:95]<=reg_A[120:127];
						endcase

						case(reg_B[100:103]) //byte12
						4'd0:
							result[96:103]<=reg_A[0:7];
						4'd1:
							result[96:103]<=reg_A[8:15];
						4'd2:
							result[96:103]<=reg_A[16:23];
						4'd3:
							result[96:103]<=reg_A[24:31];
						4'd4:
							result[96:103]<=reg_A[32:39];
						4'd5:
							result[96:103]<=reg_A[40:47];
						4'd6:
							result[96:103]<=reg_A[48:55];
						4'd7:
							result[96:103]<=reg_A[56:63];
						4'd8:
							result[96:103]<=reg_A[64:71];
						4'd9:
							result[96:103]<=reg_A[72:79];
						4'd10:
							result[96:103]<=reg_A[80:87];
						4'd11:
							result[96:103]<=reg_A[88:95];
						4'd12:
							result[96:103]<=reg_A[96:103];
						4'd13:
							result[96:103]<=reg_A[104:111];
						4'd14:
							result[96:103]<=reg_A[112:119];
						4'd15:
							result[96:103]<=reg_A[120:127];
						endcase

						case(reg_B[108:111]) //byte13
						4'd0:
							result[104:111]<=reg_A[0:7];
						4'd1:
							result[104:111]<=reg_A[8:15];
						4'd2:
							result[104:111]<=reg_A[16:23];
						4'd3:
							result[104:111]<=reg_A[24:31];
						4'd4:
							result[104:111]<=reg_A[32:39];
						4'd5:
							result[104:111]<=reg_A[40:47];
						4'd6:
							result[104:111]<=reg_A[48:55];
						4'd7:
							result[104:111]<=reg_A[56:63];
						4'd8:
							result[104:111]<=reg_A[64:71];
						4'd9:
							result[104:111]<=reg_A[72:79];
						4'd10:
							result[104:111]<=reg_A[80:87];
						4'd11:
							result[104:111]<=reg_A[88:95];
						4'd12:
							result[104:111]<=reg_A[96:103];
						4'd13:
							result[104:111]<=reg_A[104:111];
						4'd14:
							result[104:111]<=reg_A[112:119];
						4'd15:
							result[104:111]<=reg_A[120:127];
						endcase

						case(reg_B[116:119]) //byte14
						4'd0:
							result[112:119]<=reg_A[0:7];
						4'd1:
							result[112:119]<=reg_A[8:15];
						4'd2:
							result[112:119]<=reg_A[16:23];
						4'd3:
							result[112:119]<=reg_A[24:31];
						4'd4:
							result[112:119]<=reg_A[32:39];
						4'd5:
							result[112:119]<=reg_A[40:47];
						4'd6:
							result[112:119]<=reg_A[48:55];
						4'd7:
							result[112:119]<=reg_A[56:63];
						4'd8:
							result[112:119]<=reg_A[64:71];
						4'd9:
							result[112:119]<=reg_A[72:79];
						4'd10:
							result[112:119]<=reg_A[80:87];
						4'd11:
							result[112:119]<=reg_A[88:95];
						4'd12:
							result[112:119]<=reg_A[96:103];
						4'd13:
							result[112:119]<=reg_A[104:111];
						4'd14:
							result[112:119]<=reg_A[112:119];
						4'd15:
							result[112:119]<=reg_A[120:127];
						endcase

						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					`ee:	// aluwprm PRM `ee
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase

						//byte1
						result[8:15]<=8'd0;

						case(reg_B[20:23]) //byte2
						4'd0:
							result[16:23]<=reg_A[0:7];
						4'd1:
							result[16:23]<=reg_A[8:15];
						4'd2:
							result[16:23]<=reg_A[16:23];
						4'd3:
							result[16:23]<=reg_A[24:31];
						4'd4:
							result[16:23]<=reg_A[32:39];
						4'd5:
							result[16:23]<=reg_A[40:47];
						4'd6:
							result[16:23]<=reg_A[48:55];
						4'd7:
							result[16:23]<=reg_A[56:63];
						4'd8:
							result[16:23]<=reg_A[64:71];
						4'd9:
							result[16:23]<=reg_A[72:79];
						4'd10:
							result[16:23]<=reg_A[80:87];
						4'd11:
							result[16:23]<=reg_A[88:95];
						4'd12:
							result[16:23]<=reg_A[96:103];
						4'd13:
							result[16:23]<=reg_A[104:111];
						4'd14:
							result[16:23]<=reg_A[112:119];
						4'd15:
							result[16:23]<=reg_A[120:127];
						endcase

						//byte3
						result[24:31]<=8'd0;

						case(reg_B[36:39]) //byte4
						4'd0:
							result[32:39]<=reg_A[0:7];
						4'd1:
							result[32:39]<=reg_A[8:15];
						4'd2:
							result[32:39]<=reg_A[16:23];
						4'd3:
							result[32:39]<=reg_A[24:31];
						4'd4:
							result[32:39]<=reg_A[32:39];
						4'd5:
							result[32:39]<=reg_A[40:47];
						4'd6:
							result[32:39]<=reg_A[48:55];
						4'd7:
							result[32:39]<=reg_A[56:63];
						4'd8:
							result[32:39]<=reg_A[64:71];
						4'd9:
							result[32:39]<=reg_A[72:79];
						4'd10:
							result[32:39]<=reg_A[80:87];
						4'd11:
							result[32:39]<=reg_A[88:95];
						4'd12:
							result[32:39]<=reg_A[96:103];
						4'd13:
							result[32:39]<=reg_A[104:111];
						4'd14:
							result[32:39]<=reg_A[112:119];
						4'd15:
							result[32:39]<=reg_A[120:127];
						endcase

						//byte5
						result[40:47]<=8'd0;

						case(reg_B[52:55]) //byte6
						4'd0:
							result[48:55]<=reg_A[0:7];
						4'd1:
							result[48:55]<=reg_A[8:15];
						4'd2:
							result[48:55]<=reg_A[16:23];
						4'd3:
							result[48:55]<=reg_A[24:31];
						4'd4:
							result[48:55]<=reg_A[32:39];
						4'd5:
							result[48:55]<=reg_A[40:47];
						4'd6:
							result[48:55]<=reg_A[48:55];
						4'd7:
							result[48:55]<=reg_A[56:63];
						4'd8:
							result[48:55]<=reg_A[64:71];
						4'd9:
							result[48:55]<=reg_A[72:79];
						4'd10:
							result[48:55]<=reg_A[80:87];
						4'd11:
							result[48:55]<=reg_A[88:95];
						4'd12:
							result[48:55]<=reg_A[96:103];
						4'd13:
							result[48:55]<=reg_A[104:111];
						4'd14:
							result[48:55]<=reg_A[112:119];
						4'd15:
							result[48:55]<=reg_A[120:127];
						endcase

						//byte7
						result[56:63]<=8'd0;

						case(reg_B[68:71]) //byte8
						4'd0:
							result[64:71]<=reg_A[0:7];
						4'd1:
							result[64:71]<=reg_A[8:15];
						4'd2:
							result[64:71]<=reg_A[16:23];
						4'd3:
							result[64:71]<=reg_A[24:31];
						4'd4:
							result[64:71]<=reg_A[32:39];
						4'd5:
							result[64:71]<=reg_A[40:47];
						4'd6:
							result[64:71]<=reg_A[48:55];
						4'd7:
							result[64:71]<=reg_A[56:63];
						4'd8:
							result[64:71]<=reg_A[64:71];
						4'd9:
							result[64:71]<=reg_A[72:79];
						4'd10:
							result[64:71]<=reg_A[80:87];
						4'd11:
							result[64:71]<=reg_A[88:95];
						4'd12:
							result[64:71]<=reg_A[96:103];
						4'd13:
							result[64:71]<=reg_A[104:111];
						4'd14:
							result[64:71]<=reg_A[112:119];
						4'd15:
							result[64:71]<=reg_A[120:127];
						endcase

						//byte9
						result[72:79]<=8'd0;

						case(reg_B[84:87]) //byte10
						4'd0:
							result[80:87]<=reg_A[0:7];
						4'd1:
							result[80:87]<=reg_A[8:15];
						4'd2:
							result[80:87]<=reg_A[16:23];
						4'd3:
							result[80:87]<=reg_A[24:31];
						4'd4:
							result[80:87]<=reg_A[32:39];
						4'd5:
							result[80:87]<=reg_A[40:47];
						4'd6:
							result[80:87]<=reg_A[48:55];
						4'd7:
							result[80:87]<=reg_A[56:63];
						4'd8:
							result[80:87]<=reg_A[64:71];
						4'd9:
							result[80:87]<=reg_A[72:79];
						4'd10:
							result[80:87]<=reg_A[80:87];
						4'd11:
							result[80:87]<=reg_A[88:95];
						4'd12:
							result[80:87]<=reg_A[96:103];
						4'd13:
							result[80:87]<=reg_A[104:111];
						4'd14:
							result[80:87]<=reg_A[112:119];
						4'd15:
							result[80:87]<=reg_A[120:127];
						endcase

						//byte11
						result[88:95]<=8'd0;

						case(reg_B[100:103]) //byte12
						4'd0:
							result[96:103]<=reg_A[0:7];
						4'd1:
							result[96:103]<=reg_A[8:15];
						4'd2:
							result[96:103]<=reg_A[16:23];
						4'd3:
							result[96:103]<=reg_A[24:31];
						4'd4:
							result[96:103]<=reg_A[32:39];
						4'd5:
							result[96:103]<=reg_A[40:47];
						4'd6:
							result[96:103]<=reg_A[48:55];
						4'd7:
							result[96:103]<=reg_A[56:63];
						4'd8:
							result[96:103]<=reg_A[64:71];
						4'd9:
							result[96:103]<=reg_A[72:79];
						4'd10:
							result[96:103]<=reg_A[80:87];
						4'd11:
							result[96:103]<=reg_A[88:95];
						4'd12:
							result[96:103]<=reg_A[96:103];
						4'd13:
							result[96:103]<=reg_A[104:111];
						4'd14:
							result[96:103]<=reg_A[112:119];
						4'd15:
							result[96:103]<=reg_A[120:127];
						endcase

						//byte13
						result[104:111]<=8'd0;

						case(reg_B[116:119]) //byte14
						4'd0:
							result[112:119]<=reg_A[112:119];
						4'd1:
							result[112:119]<=reg_A[8:15];
						4'd2:
							result[112:119]<=reg_A[16:23];
						4'd3:
							result[112:119]<=reg_A[24:31];
						4'd4:
							result[112:119]<=reg_A[32:39];
						4'd5:
							result[112:119]<=reg_A[40:47];
						4'd6:
							result[112:119]<=reg_A[48:55];
						4'd7:
							result[112:119]<=reg_A[56:63];
						4'd8:
							result[112:119]<=reg_A[64:71];
						4'd9:
							result[112:119]<=reg_A[72:79];
						4'd10:
							result[112:119]<=reg_A[80:87];
						4'd11:
							result[112:119]<=reg_A[88:95];
						4'd12:
							result[112:119]<=reg_A[96:103];
						4'd13:
							result[112:119]<=reg_A[104:111];
						4'd14:
							result[112:119]<=reg_A[112:119];
						4'd15:
							result[112:119]<=reg_A[120:127];
						endcase

						//byte15
						result[120:127]<=8'd0;

					end
					`oo:	// aluwprm PRM `oo
					begin
						//byte0
						result[0:7]<=8'd0;

						case(reg_B[12:15]) //byte1
						4'd0:
							result[8:15]<=reg_A[0:7];
						4'd1:
							result[8:15]<=reg_A[8:15];
						4'd2:
							result[8:15]<=reg_A[16:23];
						4'd3:
							result[8:15]<=reg_A[24:31];
						4'd4:
							result[8:15]<=reg_A[32:39];
						4'd5:
							result[8:15]<=reg_A[40:47];
						4'd6:
							result[8:15]<=reg_A[48:55];
						4'd7:
							result[8:15]<=reg_A[56:63];
						4'd8:
							result[8:15]<=reg_A[64:71];
						4'd9:
							result[8:15]<=reg_A[72:79];
						4'd10:
							result[8:15]<=reg_A[80:87];
						4'd11:
							result[8:15]<=reg_A[88:95];
						4'd12:
							result[8:15]<=reg_A[96:103];
						4'd13:
							result[8:15]<=reg_A[104:111];
						4'd14:
							result[8:15]<=reg_A[112:119];
						4'd15:
							result[8:15]<=reg_A[120:127];
						endcase

						//byte2
						result[16:23]<=8'd0;

						case(reg_B[28:31]) //byte3
						4'd0:
							result[24:31]<=reg_A[0:7];
						4'd1:
							result[24:31]<=reg_A[8:15];
						4'd2:
							result[24:31]<=reg_A[16:23];
						4'd3:
							result[24:31]<=reg_A[24:31];
						4'd4:
							result[24:31]<=reg_A[32:39];
						4'd5:
							result[24:31]<=reg_A[40:47];
						4'd6:
							result[24:31]<=reg_A[48:55];
						4'd7:
							result[24:31]<=reg_A[56:63];
						4'd8:
							result[24:31]<=reg_A[64:71];
						4'd9:
							result[24:31]<=reg_A[72:79];
						4'd10:
							result[24:31]<=reg_A[80:87];
						4'd11:
							result[24:31]<=reg_A[88:95];
						4'd12:
							result[24:31]<=reg_A[96:103];
						4'd13:
							result[24:31]<=reg_A[104:111];
						4'd14:
							result[24:31]<=reg_A[112:119];
						4'd15:
							result[24:31]<=reg_A[120:127];
						endcase

						//byte4
						result[32:39]<=8'd0;

						case(reg_B[44:47]) //byte5
						4'd0:
							result[40:47]<=reg_A[0:7];
						4'd1:
							result[40:47]<=reg_A[8:15];
						4'd2:
							result[40:47]<=reg_A[16:23];
						4'd3:
							result[40:47]<=reg_A[24:31];
						4'd4:
							result[40:47]<=reg_A[32:39];
						4'd5:
							result[40:47]<=reg_A[40:47];
						4'd6:
							result[40:47]<=reg_A[48:55];
						4'd7:
							result[40:47]<=reg_A[56:63];
						4'd8:
							result[40:47]<=reg_A[64:71];
						4'd9:
							result[40:47]<=reg_A[72:79];
						4'd10:
							result[40:47]<=reg_A[80:87];
						4'd11:
							result[40:47]<=reg_A[88:95];
						4'd12:
							result[40:47]<=reg_A[96:103];
						4'd13:
							result[40:47]<=reg_A[104:111];
						4'd14:
							result[40:47]<=reg_A[112:119];
						4'd15:
							result[40:47]<=reg_A[120:127];
						endcase

						//byte6
						result[48:55]<=8'd0;

						case(reg_B[60:63]) //byte7
						4'd0:
							result[56:63]<=reg_A[0:7];
						4'd1:
							result[56:63]<=reg_A[8:15];
						4'd2:
							result[56:63]<=reg_A[16:23];
						4'd3:
							result[56:63]<=reg_A[24:31];
						4'd4:
							result[56:63]<=reg_A[32:39];
						4'd5:
							result[56:63]<=reg_A[40:47];
						4'd6:
							result[56:63]<=reg_A[48:55];
						4'd7:
							result[56:63]<=reg_A[56:63];
						4'd8:
							result[56:63]<=reg_A[64:71];
						4'd9:
							result[56:63]<=reg_A[72:79];
						4'd10:
							result[56:63]<=reg_A[80:87];
						4'd11:
							result[56:63]<=reg_A[88:95];
						4'd12:
							result[56:63]<=reg_A[96:103];
						4'd13:
							result[56:63]<=reg_A[104:111];
						4'd14:
							result[56:63]<=reg_A[112:119];
						4'd15:
							result[56:63]<=reg_A[120:127];
						endcase

						//byte8
						result[64:71]<=8'd0;

						case(reg_B[76:79]) //byte9
						4'd0:
							result[72:79]<=reg_A[0:7];
						4'd1:
							result[72:79]<=reg_A[8:15];
						4'd2:
							result[72:79]<=reg_A[16:23];
						4'd3:
							result[72:79]<=reg_A[24:31];
						4'd4:
							result[72:79]<=reg_A[32:39];
						4'd5:
							result[72:79]<=reg_A[40:47];
						4'd6:
							result[72:79]<=reg_A[48:55];
						4'd7:
							result[72:79]<=reg_A[56:63];
						4'd8:
							result[72:79]<=reg_A[64:71];
						4'd9:
							result[72:79]<=reg_A[72:79];
						4'd10:
							result[72:79]<=reg_A[80:87];
						4'd11:
							result[72:79]<=reg_A[88:95];
						4'd12:
							result[72:79]<=reg_A[96:103];
						4'd13:
							result[72:79]<=reg_A[104:111];
						4'd14:
							result[72:79]<=reg_A[112:119];
						4'd15:
							result[72:79]<=reg_A[120:127];
						endcase

						//byte10
						result[80:87]<=8'd0;
						
						case(reg_B[92:95]) //byte11
						4'd0:
							result[88:95]<=reg_A[0:7];
						4'd1:
							result[88:95]<=reg_A[8:15];
						4'd2:
							result[88:95]<=reg_A[16:23];
						4'd3:
							result[88:95]<=reg_A[24:31];
						4'd4:
							result[88:95]<=reg_A[32:39];
						4'd5:
							result[88:95]<=reg_A[40:47];
						4'd6:
							result[88:95]<=reg_A[48:55];
						4'd7:
							result[88:95]<=reg_A[56:63];
						4'd8:
							result[88:95]<=reg_A[64:71];
						4'd9:
							result[88:95]<=reg_A[72:79];
						4'd10:
							result[88:95]<=reg_A[80:87];
						4'd11:
							result[88:95]<=reg_A[88:95];
						4'd12:
							result[88:95]<=reg_A[96:103];
						4'd13:
							result[88:95]<=reg_A[104:111];
						4'd14:
							result[88:95]<=reg_A[112:119];
						4'd15:
							result[88:95]<=reg_A[120:127];
						endcase

						//byte12
						result[96:103]<=8'd0;
						
						case(reg_B[108:111]) //byte13
						4'd0:
							result[104:111]<=reg_A[0:7];
						4'd1:
							result[104:111]<=reg_A[8:15];
						4'd2:
							result[104:111]<=reg_A[16:23];
						4'd3:
							result[104:111]<=reg_A[24:31];
						4'd4:
							result[104:111]<=reg_A[32:39];
						4'd5:
							result[104:111]<=reg_A[40:47];
						4'd6:
							result[104:111]<=reg_A[48:55];
						4'd7:
							result[104:111]<=reg_A[56:63];
						4'd8:
							result[104:111]<=reg_A[64:71];
						4'd9:
							result[104:111]<=reg_A[72:79];
						4'd10:
							result[104:111]<=reg_A[80:87];
						4'd11:
							result[104:111]<=reg_A[88:95];
						4'd12:
							result[104:111]<=reg_A[96:103];
						4'd13:
							result[104:111]<=reg_A[104:111];
						4'd14:
							result[104:111]<=reg_A[112:119];
						4'd15:
							result[104:111]<=reg_A[120:127];
						endcase
						
						//byte14
						result[112:119]<=8'd0;
						
						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					`mm:	// aluwprm PRM `mm
					begin
						case(reg_B[4:7]) //byte0
						4'd0:
							result[0:7]<=reg_A[0:7];
						4'd1:
							result[0:7]<=reg_A[8:15];
						4'd2:
							result[0:7]<=reg_A[16:23];
						4'd3:
							result[0:7]<=reg_A[24:31];
						4'd4:
							result[0:7]<=reg_A[32:39];
						4'd5:
							result[0:7]<=reg_A[40:47];
						4'd6:
							result[0:7]<=reg_A[48:55];
						4'd7:
							result[0:7]<=reg_A[56:63];
						4'd8:
							result[0:7]<=reg_A[64:71];
						4'd9:
							result[0:7]<=reg_A[72:79];
						4'd10:
							result[0:7]<=reg_A[80:87];
						4'd11:
							result[0:7]<=reg_A[88:95];
						4'd12:
							result[0:7]<=reg_A[96:103];
						4'd13:
							result[0:7]<=reg_A[104:111];
						4'd14:
							result[0:7]<=reg_A[112:119];
						4'd15:
							result[0:7]<=reg_A[120:127];
						endcase
						
						//bytes1-14
						result[8:127]<=120'd0;
						
					end
					`ll:	// aluwprm PRM `ll
					begin
						//bytes0-14
						result[0:119]<=120'd0;
						
						case(reg_B[124:127]) //byte15
						4'd0:
							result[120:127]<=reg_A[0:7];
						4'd1:
							result[120:127]<=reg_A[8:15];
						4'd2:
							result[120:127]<=reg_A[16:23];
						4'd3:
							result[120:127]<=reg_A[24:31];
						4'd4:
							result[120:127]<=reg_A[32:39];
						4'd5:
							result[120:127]<=reg_A[40:47];
						4'd6:
							result[120:127]<=reg_A[48:55];
						4'd7:
							result[120:127]<=reg_A[56:63];
						4'd8:
							result[120:127]<=reg_A[64:71];
						4'd9:
							result[120:127]<=reg_A[72:79];
						4'd10:
							result[120:127]<=reg_A[80:87];
						4'd11:
							result[120:127]<=reg_A[88:95];
						4'd12:
							result[120:127]<=reg_A[96:103];
						4'd13:
							result[120:127]<=reg_A[104:111];
						4'd14:
							result[120:127]<=reg_A[112:119];
						4'd15:
							result[120:127]<=reg_A[120:127];
						endcase
					end
					default:	// aluwprm PRM Default
					begin
						result<=128'd0;
					end
				endcase
			end
			
			
			
			
			
/*
 * ========================================================
 *=========================================================
 *========================================================
 *=========================================================
 *========================================================
 *========================================================
 *=======================================================
 *========================================================
 *=======================================================
 *=======================================================
  *=========================================================
 *========================================================
 *=========================================================
 *========================================================
 *========================================================
 *=======================================================
 *========================================================
 *=======================================================
 *=======================================================
  *=========================================================
 *========================================================
 *=========================================================
 *========================================================
 *========================================================
 *=======================================================
 *========================================================
 *=======================================================
 *=======================================================
  *=========================================================
 *========================================================
 *=========================================================
 *========================================================
 *========================================================
 *=======================================================
 *========================================================
 *=======================================================
 *=======================================================
  *=========================================================
 *========================================================
 *=========================================================
 *========================================================
 *========================================================
 *=======================================================
 *========================================================
 *=======================================================
 *=======================================================
 */
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			
			// ================================================
			
			// SLLI instruction
			
			`aluwslli:
			begin
				case(ctrl_ppp)
					`aa:	// aluwslli SLLI `aa
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:15]<={reg_A[9:15],{1'b0}};
								result[16:23]<={reg_A[17:23],{1'b0}};
								result[24:31]<={reg_A[25:31],{1'b0}};
								result[32:39]<={reg_A[33:39],{1'b0}};
								result[40:47]<={reg_A[41:47],{1'b0}};
								result[48:55]<={reg_A[49:55],{1'b0}};
								result[56:63]<={reg_A[57:63],{1'b0}};
								result[64:71]<={reg_A[65:71],{1'b0}};
								result[72:79]<={reg_A[73:79],{1'b0}};
								result[80:87]<={reg_A[81:87],{1'b0}};
								result[88:95]<={reg_A[89:95],{1'b0}};
								result[96:103]<={reg_A[97:103],{1'b0}};
								result[104:111]<={reg_A[105:111],{1'b0}};
								result[112:119]<={reg_A[113:119],{1'b0}};
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:15]<={reg_A[10:15],{2{1'b0}}};
								result[16:23]<={reg_A[18:23],{2{1'b0}}};
								result[24:31]<={reg_A[26:31],{2{1'b0}}};
								result[32:39]<={reg_A[34:39],{2{1'b0}}};
								result[40:47]<={reg_A[42:47],{2{1'b0}}};
								result[48:55]<={reg_A[50:55],{2{1'b0}}};
								result[56:63]<={reg_A[58:63],{2{1'b0}}};
								result[64:71]<={reg_A[66:71],{2{1'b0}}};
								result[72:79]<={reg_A[74:79],{2{1'b0}}};
								result[80:87]<={reg_A[82:87],{2{1'b0}}};
								result[88:95]<={reg_A[90:95],{2{1'b0}}};
								result[96:103]<={reg_A[98:103],{2{1'b0}}};
								result[104:111]<={reg_A[106:111],{2{1'b0}}};
								result[112:119]<={reg_A[114:119],{2{1'b0}}};
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:15]<={reg_A[11:15],{3{1'b0}}};
								result[16:23]<={reg_A[19:23],{3{1'b0}}};
								result[24:31]<={reg_A[27:31],{3{1'b0}}};
								result[32:39]<={reg_A[35:39],{3{1'b0}}};
								result[40:47]<={reg_A[43:47],{3{1'b0}}};
								result[48:55]<={reg_A[51:55],{3{1'b0}}};
								result[56:63]<={reg_A[59:63],{3{1'b0}}};
								result[64:71]<={reg_A[67:71],{3{1'b0}}};
								result[72:79]<={reg_A[75:79],{3{1'b0}}};
								result[80:87]<={reg_A[83:87],{3{1'b0}}};
								result[88:95]<={reg_A[91:95],{3{1'b0}}};
								result[96:103]<={reg_A[99:103],{3{1'b0}}};
								result[104:111]<={reg_A[107:111],{3{1'b0}}};
								result[112:119]<={reg_A[115:119],{3{1'b0}}};
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:15]<={reg_A[12:15],{4{1'b0}}};
								result[16:23]<={reg_A[20:23],{4{1'b0}}};
								result[24:31]<={reg_A[28:31],{4{1'b0}}};
								result[32:39]<={reg_A[36:39],{4{1'b0}}};
								result[40:47]<={reg_A[44:47],{4{1'b0}}};
								result[48:55]<={reg_A[52:55],{4{1'b0}}};
								result[56:63]<={reg_A[60:63],{4{1'b0}}};
								result[64:71]<={reg_A[68:71],{4{1'b0}}};
								result[72:79]<={reg_A[76:79],{4{1'b0}}};
								result[80:87]<={reg_A[84:87],{4{1'b0}}};
								result[88:95]<={reg_A[92:95],{4{1'b0}}};
								result[96:103]<={reg_A[100:103],{4{1'b0}}};
								result[104:111]<={reg_A[108:111],{4{1'b0}}};
								result[112:119]<={reg_A[116:119],{4{1'b0}}};
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:15]<={reg_A[13:15],{5{1'b0}}};
								result[16:23]<={reg_A[21:23],{5{1'b0}}};
								result[24:31]<={reg_A[29:31],{5{1'b0}}};
								result[32:39]<={reg_A[37:39],{5{1'b0}}};
								result[40:47]<={reg_A[45:47],{5{1'b0}}};
								result[48:55]<={reg_A[53:55],{5{1'b0}}};
								result[56:63]<={reg_A[61:63],{5{1'b0}}};
								result[64:71]<={reg_A[69:71],{5{1'b0}}};
								result[72:79]<={reg_A[77:79],{5{1'b0}}};
								result[80:87]<={reg_A[85:87],{5{1'b0}}};
								result[88:95]<={reg_A[93:95],{5{1'b0}}};
								result[96:103]<={reg_A[101:103],{5{1'b0}}};
								result[104:111]<={reg_A[109:111],{5{1'b0}}};
								result[112:119]<={reg_A[117:119],{5{1'b0}}};
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:15]<={reg_A[14:15],{6{1'b0}}};
								result[16:23]<={reg_A[22:23],{6{1'b0}}};
								result[24:31]<={reg_A[30:31],{6{1'b0}}};
								result[32:39]<={reg_A[38:39],{6{1'b0}}};
								result[40:47]<={reg_A[46:47],{6{1'b0}}};
								result[48:55]<={reg_A[54:55],{6{1'b0}}};
								result[56:63]<={reg_A[62:63],{6{1'b0}}};
								result[64:71]<={reg_A[70:71],{6{1'b0}}};
								result[72:79]<={reg_A[78:79],{6{1'b0}}};
								result[80:87]<={reg_A[86:87],{6{1'b0}}};
								result[88:95]<={reg_A[94:95],{6{1'b0}}};
								result[96:103]<={reg_A[102:103],{6{1'b0}}};
								result[104:111]<={reg_A[110:111],{6{1'b0}}};
								result[112:119]<={reg_A[118:119],{6{1'b0}}};
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:15]<={reg_A[15],{7{1'b0}}};
								result[16:23]<={reg_A[23],{7{1'b0}}};
								result[24:31]<={reg_A[31],{7{1'b0}}};
								result[32:39]<={reg_A[39],{7{1'b0}}};
								result[40:47]<={reg_A[47],{7{1'b0}}};
								result[48:55]<={reg_A[55],{7{1'b0}}};
								result[56:63]<={reg_A[63],{7{1'b0}}};
								result[64:71]<={reg_A[71],{7{1'b0}}};
								result[72:79]<={reg_A[79],{7{1'b0}}};
								result[80:87]<={reg_A[87],{7{1'b0}}};
								result[88:95]<={reg_A[95],{7{1'b0}}};
								result[96:103]<={reg_A[103],{7{1'b0}}};
								result[104:111]<={reg_A[111],{7{1'b0}}};
								result[112:119]<={reg_A[119],{7{1'b0}}};
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:31]<={reg_A[17:31],{1'b0}};
								result[32:47]<={reg_A[33:47],{1'b0}};
								result[48:63]<={reg_A[49:63],{1'b0}};
								result[64:79]<={reg_A[65:79],{1'b0}};
								result[80:95]<={reg_A[81:95],{1'b0}};
								result[96:111]<={reg_A[97:111],{1'b0}};
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:31]<={reg_A[18:31],{2{1'b0}}};
								result[32:47]<={reg_A[34:47],{2{1'b0}}};
								result[48:63]<={reg_A[50:63],{2{1'b0}}};
								result[64:79]<={reg_A[66:79],{2{1'b0}}};
								result[80:95]<={reg_A[82:95],{2{1'b0}}};
								result[96:111]<={reg_A[98:111],{2{1'b0}}};
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:31]<={reg_A[19:31],{3{1'b0}}};
								result[32:47]<={reg_A[35:47],{3{1'b0}}};
								result[48:63]<={reg_A[51:63],{3{1'b0}}};
								result[64:79]<={reg_A[67:79],{3{1'b0}}};
								result[80:95]<={reg_A[83:95],{3{1'b0}}};
								result[96:111]<={reg_A[99:111],{3{1'b0}}};
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:31]<={reg_A[20:31],{4{1'b0}}};
								result[32:47]<={reg_A[36:47],{4{1'b0}}};
								result[48:63]<={reg_A[52:63],{4{1'b0}}};
								result[64:79]<={reg_A[68:79],{4{1'b0}}};
								result[80:95]<={reg_A[84:95],{4{1'b0}}};
								result[96:111]<={reg_A[100:111],{4{1'b0}}};
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:31]<={reg_A[21:31],{5{1'b0}}};
								result[32:47]<={reg_A[37:47],{5{1'b0}}};
								result[48:63]<={reg_A[52:63],{5{1'b0}}};
								result[64:79]<={reg_A[69:79],{5{1'b0}}};
								result[80:95]<={reg_A[85:95],{5{1'b0}}};
								result[96:111]<={reg_A[101:111],{5{1'b0}}};
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:31]<={reg_A[22:31],{6{1'b0}}};
								result[32:47]<={reg_A[38:47],{6{1'b0}}};
								result[48:63]<={reg_A[53:63],{6{1'b0}}};
								result[64:79]<={reg_A[70:79],{6{1'b0}}};
								result[80:95]<={reg_A[86:95],{6{1'b0}}};
								result[96:111]<={reg_A[102:111],{6{1'b0}}};
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:31]<={reg_A[23:31],{7{1'b0}}};
								result[32:47]<={reg_A[39:47],{7{1'b0}}};
								result[48:63]<={reg_A[54:63],{7{1'b0}}};
								result[64:79]<={reg_A[71:79],{7{1'b0}}};
								result[80:95]<={reg_A[87:95],{7{1'b0}}};
								result[96:111]<={reg_A[103:111],{7{1'b0}}};
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:31]<={reg_A[24:31],{8{1'b0}}};
								result[32:47]<={reg_A[40:47],{8{1'b0}}};
								result[48:63]<={reg_A[55:63],{8{1'b0}}};
								result[64:79]<={reg_A[72:79],{8{1'b0}}};
								result[80:95]<={reg_A[88:95],{8{1'b0}}};
								result[96:111]<={reg_A[104:111],{8{1'b0}}};
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:31]<={reg_A[25:31],{9{1'b0}}};
								result[32:47]<={reg_A[41:47],{9{1'b0}}};
								result[48:63]<={reg_A[56:63],{9{1'b0}}};
								result[64:79]<={reg_A[73:79],{9{1'b0}}};
								result[80:95]<={reg_A[89:95],{9{1'b0}}};
								result[96:111]<={reg_A[105:111],{9{1'b0}}};
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:31]<={reg_A[26:31],{10{1'b0}}};
								result[32:47]<={reg_A[42:47],{10{1'b0}}};
								result[48:63]<={reg_A[58:63],{10{1'b0}}};
								result[64:79]<={reg_A[74:79],{10{1'b0}}};
								result[80:95]<={reg_A[90:95],{10{1'b0}}};
								result[96:111]<={reg_A[106:111],{10{1'b0}}};
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:31]<={reg_A[27:31],{11{1'b0}}};
								result[32:47]<={reg_A[43:47],{11{1'b0}}};
								result[48:63]<={reg_A[59:63],{11{1'b0}}};
								result[64:79]<={reg_A[75:79],{11{1'b0}}};
								result[80:95]<={reg_A[91:95],{11{1'b0}}};
								result[96:111]<={reg_A[107:111],{11{1'b0}}};
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:31]<={reg_A[28:31],{12{1'b0}}};
								result[32:47]<={reg_A[44:47],{12{1'b0}}};
								result[48:63]<={reg_A[60:63],{12{1'b0}}};
								result[64:79]<={reg_A[76:79],{12{1'b0}}};
								result[80:95]<={reg_A[92:95],{12{1'b0}}};
								result[96:111]<={reg_A[108:111],{12{1'b0}}};
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:31]<={reg_A[29:31],{13{1'b0}}};
								result[32:47]<={reg_A[45:47],{13{1'b0}}};
								result[48:63]<={reg_A[61:63],{13{1'b0}}};
								result[64:79]<={reg_A[77:79],{13{1'b0}}};
								result[80:95]<={reg_A[93:95],{13{1'b0}}};
								result[96:111]<={reg_A[109:111],{13{1'b0}}};
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:31]<={reg_A[30:31],{14{1'b0}}};
								result[32:47]<={reg_A[46:47],{14{1'b0}}};
								result[48:63]<={reg_A[62:63],{14{1'b0}}};
								result[64:79]<={reg_A[78:79],{14{1'b0}}};
								result[80:95]<={reg_A[94:95],{14{1'b0}}};
								result[96:111]<={reg_A[110:111],{14{1'b0}}};
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:31]<={reg_A[31],{15{1'b0}}};
								result[32:47]<={reg_A[47],{15{1'b0}}};
								result[48:63]<={reg_A[63],{15{1'b0}}};
								result[64:79]<={reg_A[79],{15{1'b0}}};
								result[80:95]<={reg_A[95],{15{1'b0}}};
								result[96:111]<={reg_A[111],{15{1'b0}}};
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:63]<={reg_A[33:63],{1'b0}};
								result[64:95]<={reg_A[65:95],{1'b0}};
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:63]<={reg_A[34:63],{2{1'b0}}};
								result[64:95]<={reg_A[66:95],{2{1'b0}}};
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:63]<={reg_A[35:63],{3{1'b0}}};
								result[64:95]<={reg_A[67:95],{3{1'b0}}};
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:63]<={reg_A[36:63],{4{1'b0}}};
								result[64:95]<={reg_A[68:95],{4{1'b0}}};
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:63]<={reg_A[37:63],{5{1'b0}}};
								result[64:95]<={reg_A[69:95],{5{1'b0}}};
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:63]<={reg_A[38:63],{6{1'b0}}};
								result[64:95]<={reg_A[70:95],{6{1'b0}}};
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:63]<={reg_A[39:63],{7{1'b0}}};
								result[64:95]<={reg_A[71:95],{7{1'b0}}};
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:63]<={reg_A[40:63],{8{1'b0}}};
								result[64:95]<={reg_A[72:95],{8{1'b0}}};
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:63]<={reg_A[41:63],{9{1'b0}}};
								result[64:95]<={reg_A[73:95],{9{1'b0}}};
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:63]<={reg_A[42:63],{10{1'b0}}};
								result[64:95]<={reg_A[74:95],{10{1'b0}}};
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:63]<={reg_A[43:63],{11{1'b0}}};
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:63]<={reg_A[44:63],{12{1'b0}}};
								result[64:95]<={reg_A[76:95],{12{1'b0}}};
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:63]<={reg_A[45:63],{13{1'b0}}};
								result[64:95]<={reg_A[77:95],{13{1'b0}}};
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:63]<={reg_A[46:63],{14{1'b0}}};
								result[64:95]<={reg_A[78:95],{14{1'b0}}};
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:63]<={reg_A[47:63],{15{1'b0}}};
								result[64:95]<={reg_A[79:95],{15{1'b0}}};
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:63]<={reg_A[48:63],{16{1'b0}}};
								result[64:95]<={reg_A[80:95],{16{1'b0}}};
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:63]<={reg_A[49:63],{17{1'b0}}};
								result[64:95]<={reg_A[81:95],{17{1'b0}}};
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:63]<={reg_A[50:63],{18{1'b0}}};
								result[64:95]<={reg_A[82:95],{18{1'b0}}};
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:63]<={reg_A[51:63],{19{1'b0}}};
								result[64:95]<={reg_A[83:95],{19{1'b0}}};
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:63]<={reg_A[52:63],{20{1'b0}}};
								result[64:95]<={reg_A[84:95],{20{1'b0}}};
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:63]<={reg_A[53:63],{21{1'b0}}};
								result[64:95]<={reg_A[85:95],{21{1'b0}}};
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:63]<={reg_A[54:63],{22{1'b0}}};
								result[64:95]<={reg_A[86:95],{22{1'b0}}};
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:63]<={reg_A[55:63],{23{1'b0}}};
								result[64:95]<={reg_A[87:95],{23{1'b0}}};
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:63]<={reg_A[56:63],{24{1'b0}}};
								result[64:95]<={reg_A[88:95],{24{1'b0}}};
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:63]<={reg_A[57:63],{25{1'b0}}};
								result[64:95]<={reg_A[89:95],{25{1'b0}}};
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:63]<={reg_A[58:63],{26{1'b0}}};
								result[64:95]<={reg_A[90:95],{26{1'b0}}};
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:63]<={reg_A[59:63],{27{1'b0}}};
								result[64:95]<={reg_A[91:95],{27{1'b0}}};
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:63]<={reg_A[60:63],{28{1'b0}}};
								result[64:95]<={reg_A[92:95],{28{1'b0}}};
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:63]<={reg_A[61:63],{29{1'b0}}};
								result[64:95]<={reg_A[93:95],{29{1'b0}}};
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:63]<={reg_A[62:63],{30{1'b0}}};
								result[64:95]<={reg_A[94:95],{30{1'b0}}};
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:63]<={reg_A[63],{31{1'b0}}};
								result[64:95]<={reg_A[95],{31{1'b0}}};
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end
					

					`uu:	// aluwslli SLLI `uu
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:63]<=reg_A[0:63];
								result[64:127]<=64'd0;
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:15]<={reg_A[9:15],{1'b0}};
								result[16:23]<={reg_A[17:23],{1'b0}};
								result[24:31]<={reg_A[25:31],{1'b0}};
								result[32:39]<={reg_A[33:39],{1'b0}};
								result[40:47]<={reg_A[41:47],{1'b0}};
								result[48:55]<={reg_A[49:55],{1'b0}};
								result[56:63]<={reg_A[57:63],{1'b0}};
								result[64:127]<=64'd0;
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:15]<={reg_A[10:15],{2{1'b0}}};
								result[16:23]<={reg_A[18:23],{2{1'b0}}};
								result[24:31]<={reg_A[26:31],{2{1'b0}}};
								result[32:39]<={reg_A[34:39],{2{1'b0}}};
								result[40:47]<={reg_A[42:47],{2{1'b0}}};
								result[48:55]<={reg_A[50:55],{2{1'b0}}};
								result[56:63]<={reg_A[58:63],{2{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:15]<={reg_A[11:15],{3{1'b0}}};
								result[16:23]<={reg_A[19:23],{3{1'b0}}};
								result[24:31]<={reg_A[27:31],{3{1'b0}}};
								result[32:39]<={reg_A[35:39],{3{1'b0}}};
								result[40:47]<={reg_A[43:47],{3{1'b0}}};
								result[48:55]<={reg_A[51:55],{3{1'b0}}};
								result[56:63]<={reg_A[59:63],{3{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:15]<={reg_A[12:15],{4{1'b0}}};
								result[16:23]<={reg_A[20:23],{4{1'b0}}};
								result[24:31]<={reg_A[28:31],{4{1'b0}}};
								result[32:39]<={reg_A[36:39],{4{1'b0}}};
								result[40:47]<={reg_A[44:47],{4{1'b0}}};
								result[48:55]<={reg_A[52:55],{4{1'b0}}};
								result[56:63]<={reg_A[60:63],{4{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:15]<={reg_A[13:15],{5{1'b0}}};
								result[16:23]<={reg_A[21:23],{5{1'b0}}};
								result[24:31]<={reg_A[29:31],{5{1'b0}}};
								result[32:39]<={reg_A[37:39],{5{1'b0}}};
								result[40:47]<={reg_A[45:47],{5{1'b0}}};
								result[48:55]<={reg_A[53:55],{5{1'b0}}};
								result[56:63]<={reg_A[61:63],{5{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:15]<={reg_A[14:15],{6{1'b0}}};
								result[16:23]<={reg_A[22:23],{6{1'b0}}};
								result[24:31]<={reg_A[30:31],{6{1'b0}}};
								result[32:39]<={reg_A[38:39],{6{1'b0}}};
								result[40:47]<={reg_A[46:47],{6{1'b0}}};
								result[48:55]<={reg_A[54:55],{6{1'b0}}};
								result[56:63]<={reg_A[62:63],{6{1'b0}}};
								result[64:127]<=64'd0;
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:15]<={reg_A[15],{7{1'b0}}};
								result[16:23]<={reg_A[23],{7{1'b0}}};
								result[24:31]<={reg_A[31],{7{1'b0}}};
								result[32:39]<={reg_A[39],{7{1'b0}}};
								result[40:47]<={reg_A[47],{7{1'b0}}};
								result[48:55]<={reg_A[55],{7{1'b0}}};
								result[56:63]<={reg_A[63],{7{1'b0}}};
								result[64:127]<=64'd0;
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:63]<=reg_A[0:63];
								result[64:127]<=64'd0;
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:31]<={reg_A[17:31],{1'b0}};
								result[32:47]<={reg_A[33:47],{1'b0}};
								result[48:63]<={reg_A[49:63],{1'b0}};
								result[64:127]<=64'd0;
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:31]<={reg_A[18:31],{2{1'b0}}};
								result[32:47]<={reg_A[34:47],{2{1'b0}}};
								result[48:63]<={reg_A[50:63],{2{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:31]<={reg_A[19:31],{3{1'b0}}};
								result[32:47]<={reg_A[35:47],{3{1'b0}}};
								result[48:63]<={reg_A[51:63],{3{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:31]<={reg_A[20:31],{4{1'b0}}};
								result[32:47]<={reg_A[36:47],{4{1'b0}}};
								result[48:63]<={reg_A[52:63],{4{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:31]<={reg_A[21:31],{5{1'b0}}};
								result[32:47]<={reg_A[37:47],{5{1'b0}}};
								result[48:63]<={reg_A[52:63],{5{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:31]<={reg_A[22:31],{6{1'b0}}};
								result[32:47]<={reg_A[38:47],{6{1'b0}}};
								result[48:63]<={reg_A[53:63],{6{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:31]<={reg_A[23:31],{7{1'b0}}};
								result[32:47]<={reg_A[39:47],{7{1'b0}}};
								result[48:63]<={reg_A[54:63],{7{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:31]<={reg_A[24:31],{8{1'b0}}};
								result[32:47]<={reg_A[40:47],{8{1'b0}}};
								result[48:63]<={reg_A[55:63],{8{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:31]<={reg_A[25:31],{9{1'b0}}};
								result[32:47]<={reg_A[41:47],{9{1'b0}}};
								result[48:63]<={reg_A[56:63],{9{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:31]<={reg_A[26:31],{10{1'b0}}};
								result[32:47]<={reg_A[42:47],{10{1'b0}}};
								result[48:63]<={reg_A[58:63],{10{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:31]<={reg_A[27:31],{11{1'b0}}};
								result[32:47]<={reg_A[43:47],{11{1'b0}}};
								result[48:63]<={reg_A[59:63],{11{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:31]<={reg_A[28:31],{12{1'b0}}};
								result[32:47]<={reg_A[44:47],{12{1'b0}}};
								result[48:63]<={reg_A[60:63],{12{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:31]<={reg_A[29:31],{13{1'b0}}};
								result[32:47]<={reg_A[45:47],{13{1'b0}}};
								result[48:63]<={reg_A[61:63],{13{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:31]<={reg_A[30:31],{14{1'b0}}};
								result[32:47]<={reg_A[46:47],{14{1'b0}}};
								result[48:63]<={reg_A[62:63],{14{1'b0}}};
								result[64:127]<=64'd0;
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:31]<={reg_A[31],{15{1'b0}}};
								result[32:47]<={reg_A[47],{15{1'b0}}};
								result[48:63]<={reg_A[63],{15{1'b0}}};
								result[64:127]<=64'd0;
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:63]<=reg_A[0:63];
								result[64:127]<=64'd0;
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:63]<={reg_A[33:63],{1'b0}};
								result[64:127]<=64'd0;
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:63]<={reg_A[34:63],{2{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:63]<={reg_A[35:63],{3{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:63]<={reg_A[36:63],{4{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:63]<={reg_A[37:63],{5{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:63]<={reg_A[38:63],{6{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:63]<={reg_A[39:63],{7{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:63]<={reg_A[40:63],{8{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:63]<={reg_A[41:63],{9{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:63]<={reg_A[42:63],{10{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:63]<={reg_A[43:63],{11{1'b0}}};
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:63]<={reg_A[44:63],{12{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:63]<={reg_A[45:63],{13{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:63]<={reg_A[46:63],{14{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:63]<={reg_A[47:63],{15{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:63]<={reg_A[48:63],{16{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:63]<={reg_A[49:63],{17{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:63]<={reg_A[50:63],{18{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:63]<={reg_A[51:63],{19{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:63]<={reg_A[52:63],{20{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:63]<={reg_A[53:63],{21{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:63]<={reg_A[54:63],{22{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:63]<={reg_A[55:63],{23{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:63]<={reg_A[56:63],{24{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:63]<={reg_A[57:63],{25{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:63]<={reg_A[58:63],{26{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:63]<={reg_A[59:63],{27{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:63]<={reg_A[60:63],{28{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:63]<={reg_A[61:63],{29{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:63]<={reg_A[62:63],{30{1'b0}}};
								result[64:127]<=64'd0;
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:63]<={reg_A[63],{31{1'b0}}};
								result[64:127]<=64'd0;
								end
						endcase
						end
					endcase
					end

					`dd:	// aluwslli SLLI `dd
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:63]<=64'd0;
								result[64:127]<=reg_A[64:127];
								end
							3'd1:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[65:71],{1'b0}};
								result[72:79]<={reg_A[73:79],{1'b0}};
								result[80:87]<={reg_A[81:87],{1'b0}};
								result[88:95]<={reg_A[89:95],{1'b0}};
								result[96:103]<={reg_A[97:103],{1'b0}};
								result[104:111]<={reg_A[105:111],{1'b0}};
								result[112:119]<={reg_A[113:119],{1'b0}};
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[66:71],{2{1'b0}}};
								result[72:79]<={reg_A[74:79],{2{1'b0}}};
								result[80:87]<={reg_A[82:87],{2{1'b0}}};
								result[88:95]<={reg_A[90:95],{2{1'b0}}};
								result[96:103]<={reg_A[98:103],{2{1'b0}}};
								result[104:111]<={reg_A[106:111],{2{1'b0}}};
								result[112:119]<={reg_A[114:119],{2{1'b0}}};
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[67:71],{3{1'b0}}};
								result[72:79]<={reg_A[75:79],{3{1'b0}}};
								result[80:87]<={reg_A[83:87],{3{1'b0}}};
								result[88:95]<={reg_A[91:95],{3{1'b0}}};
								result[96:103]<={reg_A[99:103],{3{1'b0}}};
								result[104:111]<={reg_A[107:111],{3{1'b0}}};
								result[112:119]<={reg_A[115:119],{3{1'b0}}};
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[68:71],{4{1'b0}}};
								result[72:79]<={reg_A[76:79],{4{1'b0}}};
								result[80:87]<={reg_A[84:87],{4{1'b0}}};
								result[88:95]<={reg_A[92:95],{4{1'b0}}};
								result[96:103]<={reg_A[100:103],{4{1'b0}}};
								result[104:111]<={reg_A[108:111],{4{1'b0}}};
								result[112:119]<={reg_A[116:119],{4{1'b0}}};
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[69:71],{5{1'b0}}};
								result[72:79]<={reg_A[77:79],{5{1'b0}}};
								result[80:87]<={reg_A[85:87],{5{1'b0}}};
								result[88:95]<={reg_A[93:95],{5{1'b0}}};
								result[96:103]<={reg_A[101:103],{5{1'b0}}};
								result[104:111]<={reg_A[109:111],{5{1'b0}}};
								result[112:119]<={reg_A[117:119],{5{1'b0}}};
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[70:71],{6{1'b0}}};
								result[72:79]<={reg_A[78:79],{6{1'b0}}};
								result[80:87]<={reg_A[86:87],{6{1'b0}}};
								result[88:95]<={reg_A[94:95],{6{1'b0}}};
								result[96:103]<={reg_A[102:103],{6{1'b0}}};
								result[104:111]<={reg_A[110:111],{6{1'b0}}};
								result[112:119]<={reg_A[118:119],{6{1'b0}}};
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:63]<=64'd0;
								result[64:71]<={reg_A[71],{7{1'b0}}};
								result[72:79]<={reg_A[79],{7{1'b0}}};
								result[80:87]<={reg_A[87],{7{1'b0}}};
								result[88:95]<={reg_A[95],{7{1'b0}}};
								result[96:103]<={reg_A[103],{7{1'b0}}};
								result[104:111]<={reg_A[111],{7{1'b0}}};
								result[112:119]<={reg_A[119],{7{1'b0}}};
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:63]<=64'd0;
								result[64:127]<=reg_A[64:127];
								end
							4'd1:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[65:79],{1'b0}};
								result[80:95]<={reg_A[81:95],{1'b0}};
								result[96:111]<={reg_A[97:111],{1'b0}};
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[66:79],{2{1'b0}}};
								result[80:95]<={reg_A[82:95],{2{1'b0}}};
								result[96:111]<={reg_A[98:111],{2{1'b0}}};
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[67:79],{3{1'b0}}};
								result[80:95]<={reg_A[83:95],{3{1'b0}}};
								result[96:111]<={reg_A[99:111],{3{1'b0}}};
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[68:79],{4{1'b0}}};
								result[80:95]<={reg_A[84:95],{4{1'b0}}};
								result[96:111]<={reg_A[100:111],{4{1'b0}}};
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[69:79],{5{1'b0}}};
								result[80:95]<={reg_A[85:95],{5{1'b0}}};
								result[96:111]<={reg_A[101:111],{5{1'b0}}};
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[70:79],{6{1'b0}}};
								result[80:95]<={reg_A[86:95],{6{1'b0}}};
								result[96:111]<={reg_A[102:111],{6{1'b0}}};
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[71:79],{7{1'b0}}};
								result[80:95]<={reg_A[87:95],{7{1'b0}}};
								result[96:111]<={reg_A[103:111],{7{1'b0}}};
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[72:79],{8{1'b0}}};
								result[80:95]<={reg_A[88:95],{8{1'b0}}};
								result[96:111]<={reg_A[104:111],{8{1'b0}}};
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[73:79],{9{1'b0}}};
								result[80:95]<={reg_A[89:95],{9{1'b0}}};
								result[96:111]<={reg_A[105:111],{9{1'b0}}};
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[74:79],{10{1'b0}}};
								result[80:95]<={reg_A[90:95],{10{1'b0}}};
								result[96:111]<={reg_A[106:111],{10{1'b0}}};
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[75:79],{11{1'b0}}};
								result[80:95]<={reg_A[91:95],{11{1'b0}}};
								result[96:111]<={reg_A[107:111],{11{1'b0}}};
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[76:79],{12{1'b0}}};
								result[80:95]<={reg_A[92:95],{12{1'b0}}};
								result[96:111]<={reg_A[108:111],{12{1'b0}}};
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[77:79],{13{1'b0}}};
								result[80:95]<={reg_A[93:95],{13{1'b0}}};
								result[96:111]<={reg_A[109:111],{13{1'b0}}};
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[78:79],{14{1'b0}}};
								result[80:95]<={reg_A[94:95],{14{1'b0}}};
								result[96:111]<={reg_A[110:111],{14{1'b0}}};
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:63]<=64'd0;
								result[64:79]<={reg_A[79],{15{1'b0}}};
								result[80:95]<={reg_A[95],{15{1'b0}}};
								result[96:111]<={reg_A[111],{15{1'b0}}};
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:63]<=64'd0;
								result[64:127]<=reg_A[64:127];
								end
							5'd1:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[65:95],{1'b0}};
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[66:95],{2{1'b0}}};
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[67:95],{3{1'b0}}};
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[68:95],{4{1'b0}}};
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[69:95],{5{1'b0}}};
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[70:95],{6{1'b0}}};
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[71:95],{7{1'b0}}};
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[72:95],{8{1'b0}}};
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[73:95],{9{1'b0}}};
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[74:95],{10{1'b0}}};
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[76:95],{12{1'b0}}};
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[77:95],{13{1'b0}}};
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[78:95],{14{1'b0}}};
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[79:95],{15{1'b0}}};
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[80:95],{16{1'b0}}};
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[81:95],{17{1'b0}}};
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[82:95],{18{1'b0}}};
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[83:95],{19{1'b0}}};
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[84:95],{20{1'b0}}};
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[85:95],{21{1'b0}}};
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[86:95],{22{1'b0}}};
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[87:95],{23{1'b0}}};
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[88:95],{24{1'b0}}};
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[89:95],{25{1'b0}}};
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[90:95],{26{1'b0}}};
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[91:95],{27{1'b0}}};
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[92:95],{28{1'b0}}};
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[93:95],{29{1'b0}}};
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[94:95],{30{1'b0}}};
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:63]<=64'd0;
								result[64:95]<={reg_A[95],{31{1'b0}}};
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end

					`ee:	// aluwslli SLLI `ee
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:7]<=reg_A[0:7];
								result[8:15]<=8'b0;
								result[16:23]<=reg_A[16:23];
								result[24:31]<=8'b0;
								result[32:39]<=reg_A[33:39];
								result[40:47]<=8'b0;
								result[48:55]<=reg_A[48:55];
								result[56:63]<=8'b0;
								result[64:71]<=reg_A[64:71];
								result[72:79]<=8'b0;
								result[80:87]<=reg_A[80:87];
								result[88:95]<=8'b0;
								result[96:103]<=reg_A[96:103];
								result[104:111]<=8'b0;
								result[112:119]<=reg_A[112:119];
								result[120:127]<=8'b0;
								
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[17:23],{1'b0}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[33:39],{1'b0}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[49:55],{1'b0}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[65:71],{1'b0}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[81:87],{1'b0}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[97:103],{1'b0}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[113:119],{1'b0}};
								result[120:127]<=8'b0;
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[18:23],{2{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[34:39],{2{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[50:55],{2{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[66:71],{2{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[82:87],{2{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[98:103],{2{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[114:119],{2{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[19:23],{3{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[35:39],{3{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[51:55],{3{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[67:71],{3{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[83:87],{3{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[99:103],{3{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[115:119],{3{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[20:23],{4{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[36:39],{4{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[52:55],{4{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[68:71],{4{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[84:87],{4{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[100:103],{4{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[116:119],{4{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[21:23],{5{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[37:39],{5{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[53:55],{5{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[69:71],{5{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[85:87],{5{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[101:103],{5{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[117:119],{5{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[22:23],{6{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[38:39],{6{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[54:55],{6{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[70:71],{6{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[86:87],{6{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[102:103],{6{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[118:119],{6{1'b0}}};
								result[120:127]<=8'b0;
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:15]<=8'b0;
								result[16:23]<={reg_A[23],{7{1'b0}}};
								result[24:31]<=8'b0;
								result[32:39]<={reg_A[39],{7{1'b0}}};
								result[40:47]<=8'b0;
								result[48:55]<={reg_A[55],{7{1'b0}}};
								result[56:63]<=8'b0;
								result[64:71]<={reg_A[71],{7{1'b0}}};
								result[72:79]<=8'b0;
								result[80:87]<={reg_A[87],{7{1'b0}}};
								result[88:95]<=8'b0;
								result[96:103]<={reg_A[103],{7{1'b0}}};
								result[104:111]<=8'b0;
								result[112:119]<={reg_A[119],{7{1'b0}}};
								result[120:127]<=8'b0;
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[33:47],{1'b0}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[65:79],{1'b0}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[97:111],{1'b0}};
								result[112:127]<=16'b0;
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[34:47],{2{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[66:79],{2{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[98:111],{2{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[35:47],{3{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[67:79],{3{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[99:111],{3{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[36:47],{4{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[68:79],{4{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[100:111],{4{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[37:47],{5{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[69:79],{5{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[101:111],{5{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[38:47],{6{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[70:79],{6{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[102:111],{6{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[39:47],{7{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[71:79],{7{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[103:111],{7{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[40:47],{8{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[72:79],{8{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[104:111],{8{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[41:47],{9{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[73:79],{9{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[105:111],{9{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[42:47],{10{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[74:79],{10{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[106:111],{10{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[43:47],{11{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[75:79],{11{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[107:111],{11{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[44:47],{12{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[76:79],{12{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[108:111],{12{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[45:47],{13{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[77:79],{13{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[109:111],{13{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[46:47],{14{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[78:79],{14{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[110:111],{14{1'b0}}};
								result[112:127]<=16'b0;
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:31]<=16'b0;
								result[32:47]<={reg_A[47],{15{1'b0}}};
								result[48:63]<=16'b0;
								result[64:79]<={reg_A[79],{15{1'b0}}};
								result[80:95]<=16'b0;
								result[96:111]<={reg_A[111],{15{1'b0}}};
								result[112:127]<=16'b0;
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[65:95],{1'b0}};
								result[96:127]<=32'b0;
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[66:95],{2{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[67:95],{3{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[68:95],{4{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[69:95],{5{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[70:95],{6{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[71:95],{7{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[72:95],{8{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[73:95],{9{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[74:95],{10{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[75:95],{11{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[76:95],{12{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[77:95],{13{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[78:95],{14{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[79:95],{15{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[80:95],{16{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[81:95],{17{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[82:95],{18{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[83:95],{19{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[84:95],{20{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[85:95],{21{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[86:95],{22{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[87:95],{23{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[88:95],{24{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[89:95],{25{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[90:95],{26{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[91:95],{27{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[92:95],{28{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[93:95],{29{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[94:95],{30{1'b0}}};
								result[96:127]<=32'b0;
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:63]<=32'b0;
								result[64:95]<={reg_A[95],{31{1'b0}}};
								result[96:127]<=32'b0;
								end
						endcase
						end
					endcase
					end

					`oo:	// aluwslli SLLI `oo
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							3'd1:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[9:15],{1'b0}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[25:31],{1'b0}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[41:47],{1'b0}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[57:63],{1'b0}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[73:79],{1'b0}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[89:95],{1'b0}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[105:111],{1'b0}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[10:15],{2{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[26:31],{2{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[42:47],{2{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[58:63],{2{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[74:79],{2{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[90:95],{2{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[106:111],{2{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[11:15],{3{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[27:31],{3{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[43:47],{3{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[59:63],{3{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[75:79],{3{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[91:95],{3{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[107:111],{3{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[12:15],{4{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[28:31],{4{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[44:47],{4{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[60:63],{4{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[76:79],{4{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[92:95],{4{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[108:111],{4{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[13:15],{5{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[29:31],{5{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[45:47],{5{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[61:63],{5{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[77:79],{5{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[93:95],{5{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[109:111],{5{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[14:15],{6{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[30:31],{6{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[46:47],{6{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[62:63],{6{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[78:79],{6{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[94:95],{6{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[110:111],{6{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:7]<=8'b0;
								result[8:15]<={reg_A[15],{7{1'b0}}};
								result[16:23]<=8'b0;
								result[24:31]<={reg_A[31],{7{1'b0}}};
								result[32:39]<=8'b0;
								result[40:47]<={reg_A[47],{7{1'b0}}};
								result[48:55]<=8'b0;
								result[56:63]<={reg_A[63],{7{1'b0}}};
								result[64:71]<=8'b0;
								result[72:79]<={reg_A[79],{7{1'b0}}};
								result[80:87]<=8'b0;
								result[88:95]<={reg_A[95],{7{1'b0}}};
								result[96:103]<=8'b0;
								result[104:111]<={reg_A[111],{7{1'b0}}};
								result[112:119]<=8'b0;
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							4'd1:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[17:31],{1'b0}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[49:63],{1'b0}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[81:95],{1'b0}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[18:31],{2{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[50:63],{2{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[82:95],{2{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[19:31],{3{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[51:63],{3{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[83:95],{3{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[20:31],{4{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[52:63],{4{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[84:95],{4{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[21:31],{5{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[52:63],{5{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[85:95],{5{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[22:31],{6{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[53:63],{6{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[86:95],{6{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[23:31],{7{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[54:63],{7{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[87:95],{7{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[24:31],{8{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[55:63],{8{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[88:95],{8{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[25:31],{9{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[56:63],{9{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[89:95],{9{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[26:31],{10{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[58:63],{10{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[90:95],{10{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[27:31],{11{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[59:63],{11{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[91:95],{11{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[28:31],{12{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[60:63],{12{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[92:95],{12{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[29:31],{13{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[61:63],{13{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[93:95],{13{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[30:31],{14{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[62:63],{14{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[94:95],{14{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:15]<=16'b0;
								result[16:31]<={reg_A[31],{15{1'b0}}};
								result[32:47]<=16'b0;
								result[48:63]<={reg_A[63],{15{1'b0}}};
								result[64:79]<=16'b0;
								result[80:95]<={reg_A[95],{15{1'b0}}};
								result[96:111]<=16'b0;
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:127]<=reg_A[0:127];
								end
							5'd1:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[33:63],{1'b0}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[34:63],{2{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[35:63],{3{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[36:63],{4{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[37:63],{5{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[38:63],{6{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[39:63],{7{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[40:63],{8{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[41:63],{9{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[42:63],{10{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[43:63],{11{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[44:63],{12{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[45:63],{13{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[46:63],{14{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[47:63],{15{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[48:63],{16{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[49:63],{17{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[50:63],{18{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[51:63],{19{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[52:63],{20{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[53:63],{21{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[54:63],{22{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[55:63],{23{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[56:63],{24{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[57:63],{25{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[58:63],{26{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[59:63],{27{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[60:63],{28{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[61:63],{29{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[62:63],{30{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:31]<=32'b0;
								result[32:63]<={reg_A[63],{31{1'b0}}};
								result[64:95]<=32'b0;
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end

					`mm:	// aluwslli SLLI `mm
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:7]<=reg_A[0:7];
								result[8:127]<=119'b0;
								end
							3'd1:
								begin
								result[0:7]<={reg_A[1:7],{1'b0}};
								result[8:127]<=119'b0;
								end
							3'd2:
								begin
								result[0:7]<={reg_A[2:7],{2{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd3:
								begin
								result[0:7]<={reg_A[3:7],{3{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd4:
								begin
								result[0:7]<={reg_A[4:7],{4{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd5:
								begin
								result[0:7]<={reg_A[5:7],{5{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd6:
								begin
								result[0:7]<={reg_A[6:7],{6{1'b0}}};
								result[8:127]<=119'b0;
								end
							3'd7:
								begin
								result[0:7]<={reg_A[7],{7{1'b0}}};
								result[8:127]<=119'b0;
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:15]<=reg_A[0:15];
								result[16:127]<=112'b0;
								end
							4'd1:
								begin
								result[0:15]<={reg_A[1:15],{1'b0}};
								result[16:127]<=112'b0;
								end
							4'd2:
								begin
								result[0:15]<={reg_A[2:15],{2{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd3:
								begin
								result[0:15]<={reg_A[3:15],{3{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd4:
								begin
								result[0:15]<={reg_A[4:15],{4{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd5:
								begin
								result[0:15]<={reg_A[5:15],{5{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd6:
								begin
								result[0:15]<={reg_A[6:15],{6{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd7:
								begin
								result[0:15]<={reg_A[7:15],{7{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd8:
								begin
								result[0:15]<={reg_A[8:15],{8{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd9:
								begin
								result[0:15]<={reg_A[9:15],{9{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd10:
								begin
								result[0:15]<={reg_A[10:15],{10{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd11:
								begin
								result[0:15]<={reg_A[11:15],{11{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd12:
								begin
								result[0:15]<={reg_A[12:15],{12{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd13:
								begin
								result[0:15]<={reg_A[13:15],{13{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd14:
								begin
								result[0:15]<={reg_A[14:15],{14{1'b0}}};
								result[16:127]<=112'b0;
								end
							4'd15:
								begin
								result[0:15]<={reg_A[15],{15{1'b0}}};
								result[16:127]<=112'b0;
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:31]<=reg_A[0:31];
								result[32:127]<=96'b0;
								end
							5'd1:
								begin
								result[0:31]<={reg_A[1:31],{1'b0}};
								result[32:127]<=96'b0;
								end
							5'd2:
								begin
								result[0:31]<={reg_A[2:31],{2{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd3:
								begin
								result[0:31]<={reg_A[3:31],{3{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd4:
								begin
								result[0:31]<={reg_A[4:31],{4{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd5:
								begin
								result[0:31]<={reg_A[5:31],{5{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd6:
								begin
								result[0:31]<={reg_A[6:31],{6{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd7:
								begin
								result[0:31]<={reg_A[7:31],{7{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd8:
								begin
								result[0:31]<={reg_A[8:31],{8{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd9:
								begin
								result[0:31]<={reg_A[9:31],{9{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd10:
								begin
								result[0:31]<={reg_A[10:31],{10{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd11:
								begin
								result[0:31]<={reg_A[11:31],{11{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd12:
								begin
								result[0:31]<={reg_A[12:31],{12{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd13:
								begin
								result[0:31]<={reg_A[13:31],{13{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd14:
								begin
								result[0:31]<={reg_A[14:31],{14{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd15:
								begin
								result[0:31]<={reg_A[15:31],{15{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd16:
								begin
								result[0:31]<={reg_A[16:31],{16{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd17:
								begin
								result[0:31]<={reg_A[17:31],{17{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd18:
								begin
								result[0:31]<={reg_A[18:31],{18{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd19:
								begin
								result[0:31]<={reg_A[19:31],{19{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd20:
								begin
								result[0:31]<={reg_A[20:31],{20{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd21:
								begin
								result[0:31]<={reg_A[21:31],{21{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd22:
								begin
								result[0:31]<={reg_A[22:31],{22{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd23:
								begin
								result[0:31]<={reg_A[23:31],{23{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd24:
								begin
								result[0:31]<={reg_A[24:31],{24{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd25:
								begin
								result[0:31]<={reg_A[25:31],{25{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd26:
								begin
								result[0:31]<={reg_A[26:31],{26{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd27:
								begin
								result[0:31]<={reg_A[27:31],{27{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd28:
								begin
								result[0:31]<={reg_A[28:31],{28{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd29:
								begin
								result[0:31]<={reg_A[29:31],{29{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd30:
								begin
								result[0:31]<={reg_A[30:31],{30{1'b0}}};
								result[32:127]<=96'b0;
								end
							5'd31:
								begin
								result[0:31]<={reg_A[31],{31{1'b0}}};
								result[32:127]<=96'b0;
								end
						endcase
						end
					endcase
					end

					`ll:	// aluwslli SLLI `ll
					begin
					case(ctrl_ww)
						`w8:
						begin
						case(reg_B[2:4])
							3'd0:
								begin
								result[0:119]<=120'b0;
								result[120:127]<=reg_A[120:127];
								end
							3'd1:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[121:127],{1'b0}};
								end
							3'd2:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[122:127],{2{1'b0}}};
								end
							3'd3:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[123:127],{3{1'b0}}};
								end
							3'd4:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[124:127],{4{1'b0}}};
								end
							3'd5:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[125:127],{5{1'b0}}};
								end
							3'd6:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[126:127],{6{1'b0}}};
								end
							3'd7:
								begin
								result[0:119]<=120'b0;
								result[120:127]<={reg_A[127],{7{1'b0}}};
								end
						endcase
						end
						`w16:
						begin
						case(reg_B[1:4])
							4'd0:
								begin
								result[0:111]<=112'b0;
								result[112:127]<=reg_A[112:127];
								end
							4'd1:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[113:127],{1'b0}};
								end
							4'd2:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[114:127],{2{1'b0}}};
								end
							4'd3:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[115:127],{3{1'b0}}};
								end
							4'd4:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[116:127],{4{1'b0}}};
								end
							4'd5:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[117:127],{5{1'b0}}};
								end
							4'd6:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[118:127],{6{1'b0}}};
								end
							4'd7:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[119:127],{7{1'b0}}};
								end
							4'd8:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[120:127],{8{1'b0}}};
								end
							4'd9:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[121:127],{9{1'b0}}};
								end
							4'd10:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[122:127],{10{1'b0}}};
								end
							4'd11:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[123:127],{11{1'b0}}};
								end
							4'd12:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[124:127],{12{1'b0}}};
								end
							4'd13:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[125:127],{13{1'b0}}};
								end
							4'd14:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[126:127],{14{1'b0}}};
								end
							4'd15:
								begin
								result[0:111]<=112'b0;
								result[112:127]<={reg_A[127],{15{1'b0}}};
								end
						endcase
						end
						`w32:
						begin
						case(reg_B[0:4])
							5'd0:
								begin
								result[0:95]<=96'b0;
								result[96:127]<=reg_A[96:127];
								end
							5'd1:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[97:127],{1'b0}};
								end
							5'd2:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[98:127],{2{1'b0}}};
								end
							5'd3:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[99:127],{3{1'b0}}};
								end
							5'd4:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[100:127],{4{1'b0}}};
								end
							5'd5:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[101:127],{5{1'b0}}};
								end
							5'd6:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[102:127],{6{1'b0}}};
								end
							5'd7:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[103:127],{7{1'b0}}};
								end
							5'd8:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[104:127],{8{1'b0}}};
								end
							5'd9:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[105:127],{9{1'b0}}};
								end
							5'd10:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[106:127],{10{1'b0}}};
								end
							5'd11:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[107:127],{11{1'b0}}};
								end
							5'd12:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[108:127],{12{1'b0}}};
								end
							5'd13:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[109:127],{13{1'b0}}};
								end
							5'd14:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[110:127],{14{1'b0}}};
								end
							5'd15:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[111:127],{15{1'b0}}};
								end
							5'd16:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[112:127],{16{1'b0}}};
								end
							5'd17:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[113:127],{17{1'b0}}};
								end
							5'd18:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[114:127],{18{1'b0}}};
								end
							5'd19:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[115:127],{19{1'b0}}};
								end
							5'd20:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[116:127],{20{1'b0}}};
								end
							5'd21:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[117:127],{21{1'b0}}};
								end
							5'd22:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[118:127],{22{1'b0}}};
								end
							5'd23:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[119:127],{23{1'b0}}};
								end
							5'd24:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[120:127],{24{1'b0}}};
								end
							5'd25:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[121:127],{25{1'b0}}};
								end
							5'd26:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[122:127],{26{1'b0}}};
								end
							5'd27:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[123:127],{27{1'b0}}};
								end
							5'd28:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[124:127],{28{1'b0}}};
								end
							5'd29:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[125:127],{29{1'b0}}};
								end
							5'd30:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[126:127],{30{1'b0}}};
								end
							5'd31:
								begin
								result[0:95]<=96'b0;
								result[96:127]<={reg_A[127],{31{1'b0}}};
								end
						endcase
						end
					endcase
					end
				endcase
			end

			default:
			begin
				// Default arithmetic/logic operation
				result<=128'd0;
			end
		endcase
	end
	
	
	
	
endmodule
